-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 18 2019 12:11:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2drone
entity Pc2drone is
port (
    uart_input_pc : in std_logic;
    debug_CH5_31B : out std_logic;
    debug_CH3_20A : out std_logic;
    debug_CH0_16A : out std_logic;
    uart_input_drone : in std_logic;
    ppm_output : out std_logic;
    debug_CH6_5B : out std_logic;
    debug_CH2_18A : out std_logic;
    debug_CH4_2A : out std_logic;
    debug_CH1_0A : out std_logic;
    clk_system : in std_logic);
end Pc2drone;

-- Architecture of Pc2drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2drone is

signal \N__59697\ : std_logic;
signal \N__59683\ : std_logic;
signal \N__59682\ : std_logic;
signal \N__59681\ : std_logic;
signal \N__59674\ : std_logic;
signal \N__59673\ : std_logic;
signal \N__59672\ : std_logic;
signal \N__59665\ : std_logic;
signal \N__59664\ : std_logic;
signal \N__59663\ : std_logic;
signal \N__59656\ : std_logic;
signal \N__59655\ : std_logic;
signal \N__59654\ : std_logic;
signal \N__59647\ : std_logic;
signal \N__59646\ : std_logic;
signal \N__59645\ : std_logic;
signal \N__59638\ : std_logic;
signal \N__59637\ : std_logic;
signal \N__59636\ : std_logic;
signal \N__59629\ : std_logic;
signal \N__59628\ : std_logic;
signal \N__59627\ : std_logic;
signal \N__59620\ : std_logic;
signal \N__59619\ : std_logic;
signal \N__59618\ : std_logic;
signal \N__59611\ : std_logic;
signal \N__59610\ : std_logic;
signal \N__59609\ : std_logic;
signal \N__59602\ : std_logic;
signal \N__59601\ : std_logic;
signal \N__59600\ : std_logic;
signal \N__59583\ : std_logic;
signal \N__59580\ : std_logic;
signal \N__59577\ : std_logic;
signal \N__59574\ : std_logic;
signal \N__59573\ : std_logic;
signal \N__59572\ : std_logic;
signal \N__59569\ : std_logic;
signal \N__59566\ : std_logic;
signal \N__59563\ : std_logic;
signal \N__59560\ : std_logic;
signal \N__59557\ : std_logic;
signal \N__59554\ : std_logic;
signal \N__59551\ : std_logic;
signal \N__59546\ : std_logic;
signal \N__59543\ : std_logic;
signal \N__59538\ : std_logic;
signal \N__59535\ : std_logic;
signal \N__59532\ : std_logic;
signal \N__59529\ : std_logic;
signal \N__59528\ : std_logic;
signal \N__59527\ : std_logic;
signal \N__59520\ : std_logic;
signal \N__59517\ : std_logic;
signal \N__59514\ : std_logic;
signal \N__59511\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59505\ : std_logic;
signal \N__59502\ : std_logic;
signal \N__59501\ : std_logic;
signal \N__59500\ : std_logic;
signal \N__59497\ : std_logic;
signal \N__59492\ : std_logic;
signal \N__59487\ : std_logic;
signal \N__59484\ : std_logic;
signal \N__59481\ : std_logic;
signal \N__59478\ : std_logic;
signal \N__59475\ : std_logic;
signal \N__59472\ : std_logic;
signal \N__59469\ : std_logic;
signal \N__59466\ : std_logic;
signal \N__59463\ : std_logic;
signal \N__59460\ : std_logic;
signal \N__59459\ : std_logic;
signal \N__59458\ : std_logic;
signal \N__59455\ : std_logic;
signal \N__59452\ : std_logic;
signal \N__59449\ : std_logic;
signal \N__59446\ : std_logic;
signal \N__59443\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59433\ : std_logic;
signal \N__59430\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59426\ : std_logic;
signal \N__59425\ : std_logic;
signal \N__59418\ : std_logic;
signal \N__59415\ : std_logic;
signal \N__59412\ : std_logic;
signal \N__59409\ : std_logic;
signal \N__59406\ : std_logic;
signal \N__59403\ : std_logic;
signal \N__59400\ : std_logic;
signal \N__59397\ : std_logic;
signal \N__59396\ : std_logic;
signal \N__59395\ : std_logic;
signal \N__59392\ : std_logic;
signal \N__59387\ : std_logic;
signal \N__59382\ : std_logic;
signal \N__59379\ : std_logic;
signal \N__59376\ : std_logic;
signal \N__59373\ : std_logic;
signal \N__59370\ : std_logic;
signal \N__59367\ : std_logic;
signal \N__59364\ : std_logic;
signal \N__59361\ : std_logic;
signal \N__59360\ : std_logic;
signal \N__59359\ : std_logic;
signal \N__59352\ : std_logic;
signal \N__59349\ : std_logic;
signal \N__59346\ : std_logic;
signal \N__59343\ : std_logic;
signal \N__59340\ : std_logic;
signal \N__59337\ : std_logic;
signal \N__59336\ : std_logic;
signal \N__59335\ : std_logic;
signal \N__59334\ : std_logic;
signal \N__59333\ : std_logic;
signal \N__59332\ : std_logic;
signal \N__59331\ : std_logic;
signal \N__59330\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59328\ : std_logic;
signal \N__59327\ : std_logic;
signal \N__59326\ : std_logic;
signal \N__59325\ : std_logic;
signal \N__59324\ : std_logic;
signal \N__59323\ : std_logic;
signal \N__59322\ : std_logic;
signal \N__59321\ : std_logic;
signal \N__59320\ : std_logic;
signal \N__59319\ : std_logic;
signal \N__59318\ : std_logic;
signal \N__59317\ : std_logic;
signal \N__59316\ : std_logic;
signal \N__59315\ : std_logic;
signal \N__59314\ : std_logic;
signal \N__59313\ : std_logic;
signal \N__59312\ : std_logic;
signal \N__59311\ : std_logic;
signal \N__59310\ : std_logic;
signal \N__59309\ : std_logic;
signal \N__59308\ : std_logic;
signal \N__59307\ : std_logic;
signal \N__59306\ : std_logic;
signal \N__59305\ : std_logic;
signal \N__59304\ : std_logic;
signal \N__59303\ : std_logic;
signal \N__59302\ : std_logic;
signal \N__59301\ : std_logic;
signal \N__59300\ : std_logic;
signal \N__59299\ : std_logic;
signal \N__59298\ : std_logic;
signal \N__59297\ : std_logic;
signal \N__59296\ : std_logic;
signal \N__59295\ : std_logic;
signal \N__59294\ : std_logic;
signal \N__59293\ : std_logic;
signal \N__59292\ : std_logic;
signal \N__59291\ : std_logic;
signal \N__59290\ : std_logic;
signal \N__59289\ : std_logic;
signal \N__59288\ : std_logic;
signal \N__59287\ : std_logic;
signal \N__59286\ : std_logic;
signal \N__59285\ : std_logic;
signal \N__59284\ : std_logic;
signal \N__59283\ : std_logic;
signal \N__59282\ : std_logic;
signal \N__59281\ : std_logic;
signal \N__59280\ : std_logic;
signal \N__59279\ : std_logic;
signal \N__59278\ : std_logic;
signal \N__59277\ : std_logic;
signal \N__59276\ : std_logic;
signal \N__59275\ : std_logic;
signal \N__59274\ : std_logic;
signal \N__59273\ : std_logic;
signal \N__59272\ : std_logic;
signal \N__59271\ : std_logic;
signal \N__59270\ : std_logic;
signal \N__59269\ : std_logic;
signal \N__59268\ : std_logic;
signal \N__59267\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59265\ : std_logic;
signal \N__59264\ : std_logic;
signal \N__59263\ : std_logic;
signal \N__59262\ : std_logic;
signal \N__59261\ : std_logic;
signal \N__59260\ : std_logic;
signal \N__59259\ : std_logic;
signal \N__59258\ : std_logic;
signal \N__59257\ : std_logic;
signal \N__59256\ : std_logic;
signal \N__59255\ : std_logic;
signal \N__59254\ : std_logic;
signal \N__59253\ : std_logic;
signal \N__59252\ : std_logic;
signal \N__59251\ : std_logic;
signal \N__59250\ : std_logic;
signal \N__59249\ : std_logic;
signal \N__59248\ : std_logic;
signal \N__59247\ : std_logic;
signal \N__59246\ : std_logic;
signal \N__59245\ : std_logic;
signal \N__59244\ : std_logic;
signal \N__59243\ : std_logic;
signal \N__59242\ : std_logic;
signal \N__59241\ : std_logic;
signal \N__59240\ : std_logic;
signal \N__59239\ : std_logic;
signal \N__59238\ : std_logic;
signal \N__59237\ : std_logic;
signal \N__59236\ : std_logic;
signal \N__59235\ : std_logic;
signal \N__59234\ : std_logic;
signal \N__59233\ : std_logic;
signal \N__59232\ : std_logic;
signal \N__59231\ : std_logic;
signal \N__59230\ : std_logic;
signal \N__59229\ : std_logic;
signal \N__59228\ : std_logic;
signal \N__59227\ : std_logic;
signal \N__59226\ : std_logic;
signal \N__59225\ : std_logic;
signal \N__59224\ : std_logic;
signal \N__59223\ : std_logic;
signal \N__59222\ : std_logic;
signal \N__59221\ : std_logic;
signal \N__59220\ : std_logic;
signal \N__59219\ : std_logic;
signal \N__59218\ : std_logic;
signal \N__59217\ : std_logic;
signal \N__59216\ : std_logic;
signal \N__59215\ : std_logic;
signal \N__59214\ : std_logic;
signal \N__59213\ : std_logic;
signal \N__59212\ : std_logic;
signal \N__59211\ : std_logic;
signal \N__59210\ : std_logic;
signal \N__59209\ : std_logic;
signal \N__59208\ : std_logic;
signal \N__59207\ : std_logic;
signal \N__59206\ : std_logic;
signal \N__59205\ : std_logic;
signal \N__59204\ : std_logic;
signal \N__59203\ : std_logic;
signal \N__59202\ : std_logic;
signal \N__59201\ : std_logic;
signal \N__59200\ : std_logic;
signal \N__59199\ : std_logic;
signal \N__59198\ : std_logic;
signal \N__59197\ : std_logic;
signal \N__59196\ : std_logic;
signal \N__59195\ : std_logic;
signal \N__59194\ : std_logic;
signal \N__59193\ : std_logic;
signal \N__59192\ : std_logic;
signal \N__59191\ : std_logic;
signal \N__59190\ : std_logic;
signal \N__59189\ : std_logic;
signal \N__59188\ : std_logic;
signal \N__59187\ : std_logic;
signal \N__59186\ : std_logic;
signal \N__59185\ : std_logic;
signal \N__59184\ : std_logic;
signal \N__59183\ : std_logic;
signal \N__59182\ : std_logic;
signal \N__59181\ : std_logic;
signal \N__59180\ : std_logic;
signal \N__59179\ : std_logic;
signal \N__59178\ : std_logic;
signal \N__59177\ : std_logic;
signal \N__59176\ : std_logic;
signal \N__59175\ : std_logic;
signal \N__59174\ : std_logic;
signal \N__59173\ : std_logic;
signal \N__59172\ : std_logic;
signal \N__59171\ : std_logic;
signal \N__59170\ : std_logic;
signal \N__59169\ : std_logic;
signal \N__59168\ : std_logic;
signal \N__59167\ : std_logic;
signal \N__59166\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59164\ : std_logic;
signal \N__59163\ : std_logic;
signal \N__59162\ : std_logic;
signal \N__59161\ : std_logic;
signal \N__59160\ : std_logic;
signal \N__59159\ : std_logic;
signal \N__59158\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59156\ : std_logic;
signal \N__59155\ : std_logic;
signal \N__59154\ : std_logic;
signal \N__59153\ : std_logic;
signal \N__59152\ : std_logic;
signal \N__59151\ : std_logic;
signal \N__59150\ : std_logic;
signal \N__59149\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59147\ : std_logic;
signal \N__59146\ : std_logic;
signal \N__59145\ : std_logic;
signal \N__59144\ : std_logic;
signal \N__59143\ : std_logic;
signal \N__59142\ : std_logic;
signal \N__59141\ : std_logic;
signal \N__59140\ : std_logic;
signal \N__59139\ : std_logic;
signal \N__59138\ : std_logic;
signal \N__59137\ : std_logic;
signal \N__59136\ : std_logic;
signal \N__59135\ : std_logic;
signal \N__59134\ : std_logic;
signal \N__59133\ : std_logic;
signal \N__59132\ : std_logic;
signal \N__59131\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59129\ : std_logic;
signal \N__59128\ : std_logic;
signal \N__59127\ : std_logic;
signal \N__59126\ : std_logic;
signal \N__59125\ : std_logic;
signal \N__59124\ : std_logic;
signal \N__59123\ : std_logic;
signal \N__59122\ : std_logic;
signal \N__59121\ : std_logic;
signal \N__59120\ : std_logic;
signal \N__59119\ : std_logic;
signal \N__59118\ : std_logic;
signal \N__59117\ : std_logic;
signal \N__59116\ : std_logic;
signal \N__59115\ : std_logic;
signal \N__59114\ : std_logic;
signal \N__59113\ : std_logic;
signal \N__59112\ : std_logic;
signal \N__59111\ : std_logic;
signal \N__59110\ : std_logic;
signal \N__59109\ : std_logic;
signal \N__59108\ : std_logic;
signal \N__59107\ : std_logic;
signal \N__59106\ : std_logic;
signal \N__59105\ : std_logic;
signal \N__59104\ : std_logic;
signal \N__59103\ : std_logic;
signal \N__59102\ : std_logic;
signal \N__59101\ : std_logic;
signal \N__59100\ : std_logic;
signal \N__59099\ : std_logic;
signal \N__59098\ : std_logic;
signal \N__59097\ : std_logic;
signal \N__59096\ : std_logic;
signal \N__59095\ : std_logic;
signal \N__59094\ : std_logic;
signal \N__59093\ : std_logic;
signal \N__59092\ : std_logic;
signal \N__59091\ : std_logic;
signal \N__59090\ : std_logic;
signal \N__59089\ : std_logic;
signal \N__59088\ : std_logic;
signal \N__59087\ : std_logic;
signal \N__59086\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59084\ : std_logic;
signal \N__59083\ : std_logic;
signal \N__59082\ : std_logic;
signal \N__59081\ : std_logic;
signal \N__59080\ : std_logic;
signal \N__59079\ : std_logic;
signal \N__59078\ : std_logic;
signal \N__59077\ : std_logic;
signal \N__59076\ : std_logic;
signal \N__59075\ : std_logic;
signal \N__59074\ : std_logic;
signal \N__58545\ : std_logic;
signal \N__58542\ : std_logic;
signal \N__58539\ : std_logic;
signal \N__58538\ : std_logic;
signal \N__58537\ : std_logic;
signal \N__58536\ : std_logic;
signal \N__58535\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58531\ : std_logic;
signal \N__58528\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58524\ : std_logic;
signal \N__58523\ : std_logic;
signal \N__58520\ : std_logic;
signal \N__58517\ : std_logic;
signal \N__58514\ : std_logic;
signal \N__58511\ : std_logic;
signal \N__58508\ : std_logic;
signal \N__58507\ : std_logic;
signal \N__58504\ : std_logic;
signal \N__58503\ : std_logic;
signal \N__58502\ : std_logic;
signal \N__58499\ : std_logic;
signal \N__58496\ : std_logic;
signal \N__58495\ : std_logic;
signal \N__58494\ : std_logic;
signal \N__58491\ : std_logic;
signal \N__58486\ : std_logic;
signal \N__58483\ : std_logic;
signal \N__58480\ : std_logic;
signal \N__58477\ : std_logic;
signal \N__58474\ : std_logic;
signal \N__58471\ : std_logic;
signal \N__58468\ : std_logic;
signal \N__58465\ : std_logic;
signal \N__58462\ : std_logic;
signal \N__58459\ : std_logic;
signal \N__58456\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58450\ : std_logic;
signal \N__58449\ : std_logic;
signal \N__58446\ : std_logic;
signal \N__58443\ : std_logic;
signal \N__58440\ : std_logic;
signal \N__58435\ : std_logic;
signal \N__58432\ : std_logic;
signal \N__58423\ : std_logic;
signal \N__58420\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58414\ : std_logic;
signal \N__58411\ : std_logic;
signal \N__58408\ : std_logic;
signal \N__58405\ : std_logic;
signal \N__58402\ : std_logic;
signal \N__58395\ : std_logic;
signal \N__58392\ : std_logic;
signal \N__58389\ : std_logic;
signal \N__58386\ : std_logic;
signal \N__58383\ : std_logic;
signal \N__58378\ : std_logic;
signal \N__58375\ : std_logic;
signal \N__58370\ : std_logic;
signal \N__58359\ : std_logic;
signal \N__58358\ : std_logic;
signal \N__58357\ : std_logic;
signal \N__58356\ : std_logic;
signal \N__58355\ : std_logic;
signal \N__58354\ : std_logic;
signal \N__58353\ : std_logic;
signal \N__58352\ : std_logic;
signal \N__58351\ : std_logic;
signal \N__58350\ : std_logic;
signal \N__58349\ : std_logic;
signal \N__58348\ : std_logic;
signal \N__58347\ : std_logic;
signal \N__58346\ : std_logic;
signal \N__58345\ : std_logic;
signal \N__58344\ : std_logic;
signal \N__58343\ : std_logic;
signal \N__58342\ : std_logic;
signal \N__58341\ : std_logic;
signal \N__58340\ : std_logic;
signal \N__58339\ : std_logic;
signal \N__58338\ : std_logic;
signal \N__58337\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58335\ : std_logic;
signal \N__58334\ : std_logic;
signal \N__58333\ : std_logic;
signal \N__58332\ : std_logic;
signal \N__58331\ : std_logic;
signal \N__58330\ : std_logic;
signal \N__58329\ : std_logic;
signal \N__58328\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58326\ : std_logic;
signal \N__58325\ : std_logic;
signal \N__58324\ : std_logic;
signal \N__58323\ : std_logic;
signal \N__58322\ : std_logic;
signal \N__58321\ : std_logic;
signal \N__58320\ : std_logic;
signal \N__58319\ : std_logic;
signal \N__58314\ : std_logic;
signal \N__58305\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58295\ : std_logic;
signal \N__58286\ : std_logic;
signal \N__58281\ : std_logic;
signal \N__58276\ : std_logic;
signal \N__58265\ : std_logic;
signal \N__58262\ : std_logic;
signal \N__58257\ : std_logic;
signal \N__58252\ : std_logic;
signal \N__58247\ : std_logic;
signal \N__58232\ : std_logic;
signal \N__58229\ : std_logic;
signal \N__58226\ : std_logic;
signal \N__58223\ : std_logic;
signal \N__58220\ : std_logic;
signal \N__58219\ : std_logic;
signal \N__58218\ : std_logic;
signal \N__58217\ : std_logic;
signal \N__58216\ : std_logic;
signal \N__58215\ : std_logic;
signal \N__58214\ : std_logic;
signal \N__58213\ : std_logic;
signal \N__58212\ : std_logic;
signal \N__58211\ : std_logic;
signal \N__58210\ : std_logic;
signal \N__58209\ : std_logic;
signal \N__58208\ : std_logic;
signal \N__58207\ : std_logic;
signal \N__58206\ : std_logic;
signal \N__58205\ : std_logic;
signal \N__58204\ : std_logic;
signal \N__58203\ : std_logic;
signal \N__58202\ : std_logic;
signal \N__58201\ : std_logic;
signal \N__58200\ : std_logic;
signal \N__58199\ : std_logic;
signal \N__58198\ : std_logic;
signal \N__58197\ : std_logic;
signal \N__58196\ : std_logic;
signal \N__58195\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58193\ : std_logic;
signal \N__58192\ : std_logic;
signal \N__58191\ : std_logic;
signal \N__58190\ : std_logic;
signal \N__58189\ : std_logic;
signal \N__58188\ : std_logic;
signal \N__58187\ : std_logic;
signal \N__58186\ : std_logic;
signal \N__58185\ : std_logic;
signal \N__58184\ : std_logic;
signal \N__58183\ : std_logic;
signal \N__58182\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58180\ : std_logic;
signal \N__58179\ : std_logic;
signal \N__58176\ : std_logic;
signal \N__58173\ : std_logic;
signal \N__58170\ : std_logic;
signal \N__58167\ : std_logic;
signal \N__58164\ : std_logic;
signal \N__58161\ : std_logic;
signal \N__58158\ : std_logic;
signal \N__58155\ : std_logic;
signal \N__58152\ : std_logic;
signal \N__58149\ : std_logic;
signal \N__58146\ : std_logic;
signal \N__58143\ : std_logic;
signal \N__58140\ : std_logic;
signal \N__58137\ : std_logic;
signal \N__58134\ : std_logic;
signal \N__58131\ : std_logic;
signal \N__58128\ : std_logic;
signal \N__58011\ : std_logic;
signal \N__58008\ : std_logic;
signal \N__58005\ : std_logic;
signal \N__58004\ : std_logic;
signal \N__58001\ : std_logic;
signal \N__57998\ : std_logic;
signal \N__57997\ : std_logic;
signal \N__57994\ : std_logic;
signal \N__57991\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57981\ : std_logic;
signal \N__57980\ : std_logic;
signal \N__57977\ : std_logic;
signal \N__57974\ : std_logic;
signal \N__57969\ : std_logic;
signal \N__57966\ : std_logic;
signal \N__57965\ : std_logic;
signal \N__57964\ : std_logic;
signal \N__57963\ : std_logic;
signal \N__57962\ : std_logic;
signal \N__57961\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57959\ : std_logic;
signal \N__57958\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57956\ : std_logic;
signal \N__57955\ : std_logic;
signal \N__57954\ : std_logic;
signal \N__57953\ : std_logic;
signal \N__57952\ : std_logic;
signal \N__57951\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57949\ : std_logic;
signal \N__57948\ : std_logic;
signal \N__57909\ : std_logic;
signal \N__57906\ : std_logic;
signal \N__57903\ : std_logic;
signal \N__57902\ : std_logic;
signal \N__57901\ : std_logic;
signal \N__57900\ : std_logic;
signal \N__57897\ : std_logic;
signal \N__57896\ : std_logic;
signal \N__57895\ : std_logic;
signal \N__57894\ : std_logic;
signal \N__57891\ : std_logic;
signal \N__57890\ : std_logic;
signal \N__57889\ : std_logic;
signal \N__57888\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57886\ : std_logic;
signal \N__57885\ : std_logic;
signal \N__57884\ : std_logic;
signal \N__57883\ : std_logic;
signal \N__57882\ : std_logic;
signal \N__57881\ : std_logic;
signal \N__57880\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57878\ : std_logic;
signal \N__57877\ : std_logic;
signal \N__57876\ : std_logic;
signal \N__57875\ : std_logic;
signal \N__57872\ : std_logic;
signal \N__57871\ : std_logic;
signal \N__57870\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57868\ : std_logic;
signal \N__57867\ : std_logic;
signal \N__57866\ : std_logic;
signal \N__57865\ : std_logic;
signal \N__57864\ : std_logic;
signal \N__57863\ : std_logic;
signal \N__57862\ : std_logic;
signal \N__57861\ : std_logic;
signal \N__57860\ : std_logic;
signal \N__57859\ : std_logic;
signal \N__57858\ : std_logic;
signal \N__57857\ : std_logic;
signal \N__57856\ : std_logic;
signal \N__57855\ : std_logic;
signal \N__57854\ : std_logic;
signal \N__57853\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57851\ : std_logic;
signal \N__57850\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57848\ : std_logic;
signal \N__57847\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57845\ : std_logic;
signal \N__57844\ : std_logic;
signal \N__57843\ : std_logic;
signal \N__57842\ : std_logic;
signal \N__57841\ : std_logic;
signal \N__57838\ : std_logic;
signal \N__57837\ : std_logic;
signal \N__57836\ : std_logic;
signal \N__57835\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57833\ : std_logic;
signal \N__57832\ : std_logic;
signal \N__57831\ : std_logic;
signal \N__57830\ : std_logic;
signal \N__57829\ : std_logic;
signal \N__57828\ : std_logic;
signal \N__57827\ : std_logic;
signal \N__57824\ : std_logic;
signal \N__57821\ : std_logic;
signal \N__57818\ : std_logic;
signal \N__57811\ : std_logic;
signal \N__57808\ : std_logic;
signal \N__57799\ : std_logic;
signal \N__57794\ : std_logic;
signal \N__57787\ : std_logic;
signal \N__57782\ : std_logic;
signal \N__57775\ : std_logic;
signal \N__57770\ : std_logic;
signal \N__57767\ : std_logic;
signal \N__57760\ : std_logic;
signal \N__57757\ : std_logic;
signal \N__57754\ : std_logic;
signal \N__57751\ : std_logic;
signal \N__57746\ : std_logic;
signal \N__57743\ : std_logic;
signal \N__57740\ : std_logic;
signal \N__57737\ : std_logic;
signal \N__57734\ : std_logic;
signal \N__57727\ : std_logic;
signal \N__57724\ : std_logic;
signal \N__57719\ : std_logic;
signal \N__57716\ : std_logic;
signal \N__57713\ : std_logic;
signal \N__57710\ : std_logic;
signal \N__57707\ : std_logic;
signal \N__57704\ : std_logic;
signal \N__57701\ : std_logic;
signal \N__57698\ : std_logic;
signal \N__57695\ : std_logic;
signal \N__57690\ : std_logic;
signal \N__57687\ : std_logic;
signal \N__57684\ : std_logic;
signal \N__57681\ : std_logic;
signal \N__57678\ : std_logic;
signal \N__57675\ : std_logic;
signal \N__57672\ : std_logic;
signal \N__57669\ : std_logic;
signal \N__57666\ : std_logic;
signal \N__57663\ : std_logic;
signal \N__57660\ : std_logic;
signal \N__57657\ : std_logic;
signal \N__57654\ : std_logic;
signal \N__57651\ : std_logic;
signal \N__57650\ : std_logic;
signal \N__57649\ : std_logic;
signal \N__57648\ : std_logic;
signal \N__57647\ : std_logic;
signal \N__57646\ : std_logic;
signal \N__57645\ : std_logic;
signal \N__57644\ : std_logic;
signal \N__57643\ : std_logic;
signal \N__57642\ : std_logic;
signal \N__57641\ : std_logic;
signal \N__57640\ : std_logic;
signal \N__57639\ : std_logic;
signal \N__57638\ : std_logic;
signal \N__57637\ : std_logic;
signal \N__57636\ : std_logic;
signal \N__57635\ : std_logic;
signal \N__57634\ : std_logic;
signal \N__57633\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57631\ : std_logic;
signal \N__57630\ : std_logic;
signal \N__57629\ : std_logic;
signal \N__57628\ : std_logic;
signal \N__57627\ : std_logic;
signal \N__57626\ : std_logic;
signal \N__57625\ : std_logic;
signal \N__57624\ : std_logic;
signal \N__57623\ : std_logic;
signal \N__57622\ : std_logic;
signal \N__57621\ : std_logic;
signal \N__57620\ : std_logic;
signal \N__57619\ : std_logic;
signal \N__57618\ : std_logic;
signal \N__57617\ : std_logic;
signal \N__57616\ : std_logic;
signal \N__57615\ : std_logic;
signal \N__57614\ : std_logic;
signal \N__57613\ : std_logic;
signal \N__57612\ : std_logic;
signal \N__57611\ : std_logic;
signal \N__57610\ : std_logic;
signal \N__57609\ : std_logic;
signal \N__57608\ : std_logic;
signal \N__57607\ : std_logic;
signal \N__57606\ : std_logic;
signal \N__57605\ : std_logic;
signal \N__57604\ : std_logic;
signal \N__57603\ : std_logic;
signal \N__57602\ : std_logic;
signal \N__57601\ : std_logic;
signal \N__57600\ : std_logic;
signal \N__57599\ : std_logic;
signal \N__57598\ : std_logic;
signal \N__57597\ : std_logic;
signal \N__57596\ : std_logic;
signal \N__57595\ : std_logic;
signal \N__57594\ : std_logic;
signal \N__57593\ : std_logic;
signal \N__57592\ : std_logic;
signal \N__57591\ : std_logic;
signal \N__57590\ : std_logic;
signal \N__57589\ : std_logic;
signal \N__57588\ : std_logic;
signal \N__57587\ : std_logic;
signal \N__57586\ : std_logic;
signal \N__57585\ : std_logic;
signal \N__57584\ : std_logic;
signal \N__57583\ : std_logic;
signal \N__57582\ : std_logic;
signal \N__57581\ : std_logic;
signal \N__57580\ : std_logic;
signal \N__57579\ : std_logic;
signal \N__57578\ : std_logic;
signal \N__57577\ : std_logic;
signal \N__57576\ : std_logic;
signal \N__57575\ : std_logic;
signal \N__57574\ : std_logic;
signal \N__57573\ : std_logic;
signal \N__57572\ : std_logic;
signal \N__57571\ : std_logic;
signal \N__57570\ : std_logic;
signal \N__57569\ : std_logic;
signal \N__57568\ : std_logic;
signal \N__57567\ : std_logic;
signal \N__57566\ : std_logic;
signal \N__57565\ : std_logic;
signal \N__57564\ : std_logic;
signal \N__57563\ : std_logic;
signal \N__57562\ : std_logic;
signal \N__57561\ : std_logic;
signal \N__57560\ : std_logic;
signal \N__57559\ : std_logic;
signal \N__57558\ : std_logic;
signal \N__57557\ : std_logic;
signal \N__57556\ : std_logic;
signal \N__57555\ : std_logic;
signal \N__57554\ : std_logic;
signal \N__57553\ : std_logic;
signal \N__57552\ : std_logic;
signal \N__57551\ : std_logic;
signal \N__57550\ : std_logic;
signal \N__57549\ : std_logic;
signal \N__57548\ : std_logic;
signal \N__57547\ : std_logic;
signal \N__57546\ : std_logic;
signal \N__57545\ : std_logic;
signal \N__57544\ : std_logic;
signal \N__57543\ : std_logic;
signal \N__57542\ : std_logic;
signal \N__57541\ : std_logic;
signal \N__57540\ : std_logic;
signal \N__57539\ : std_logic;
signal \N__57538\ : std_logic;
signal \N__57537\ : std_logic;
signal \N__57536\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57534\ : std_logic;
signal \N__57533\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57531\ : std_logic;
signal \N__57530\ : std_logic;
signal \N__57529\ : std_logic;
signal \N__57528\ : std_logic;
signal \N__57527\ : std_logic;
signal \N__57526\ : std_logic;
signal \N__57525\ : std_logic;
signal \N__57524\ : std_logic;
signal \N__57523\ : std_logic;
signal \N__57522\ : std_logic;
signal \N__57521\ : std_logic;
signal \N__57520\ : std_logic;
signal \N__57519\ : std_logic;
signal \N__57518\ : std_logic;
signal \N__57517\ : std_logic;
signal \N__57516\ : std_logic;
signal \N__57515\ : std_logic;
signal \N__57514\ : std_logic;
signal \N__57513\ : std_logic;
signal \N__57512\ : std_logic;
signal \N__57511\ : std_logic;
signal \N__57510\ : std_logic;
signal \N__57509\ : std_logic;
signal \N__57508\ : std_logic;
signal \N__57507\ : std_logic;
signal \N__57506\ : std_logic;
signal \N__57505\ : std_logic;
signal \N__57504\ : std_logic;
signal \N__57503\ : std_logic;
signal \N__57502\ : std_logic;
signal \N__57501\ : std_logic;
signal \N__57500\ : std_logic;
signal \N__57499\ : std_logic;
signal \N__57498\ : std_logic;
signal \N__57497\ : std_logic;
signal \N__57496\ : std_logic;
signal \N__57493\ : std_logic;
signal \N__57490\ : std_logic;
signal \N__57487\ : std_logic;
signal \N__57484\ : std_logic;
signal \N__57481\ : std_logic;
signal \N__57478\ : std_logic;
signal \N__57475\ : std_logic;
signal \N__57472\ : std_logic;
signal \N__57469\ : std_logic;
signal \N__57466\ : std_logic;
signal \N__57463\ : std_logic;
signal \N__57460\ : std_logic;
signal \N__57457\ : std_logic;
signal \N__57454\ : std_logic;
signal \N__57451\ : std_logic;
signal \N__57448\ : std_logic;
signal \N__57445\ : std_logic;
signal \N__57442\ : std_logic;
signal \N__57439\ : std_logic;
signal \N__57436\ : std_logic;
signal \N__57433\ : std_logic;
signal \N__57430\ : std_logic;
signal \N__57427\ : std_logic;
signal \N__57424\ : std_logic;
signal \N__57421\ : std_logic;
signal \N__57418\ : std_logic;
signal \N__57415\ : std_logic;
signal \N__57412\ : std_logic;
signal \N__57409\ : std_logic;
signal \N__57406\ : std_logic;
signal \N__57403\ : std_logic;
signal \N__57400\ : std_logic;
signal \N__57397\ : std_logic;
signal \N__57394\ : std_logic;
signal \N__57391\ : std_logic;
signal \N__57388\ : std_logic;
signal \N__57385\ : std_logic;
signal \N__57382\ : std_logic;
signal \N__57379\ : std_logic;
signal \N__57376\ : std_logic;
signal \N__57373\ : std_logic;
signal \N__57370\ : std_logic;
signal \N__57367\ : std_logic;
signal \N__57364\ : std_logic;
signal \N__57361\ : std_logic;
signal \N__57358\ : std_logic;
signal \N__56955\ : std_logic;
signal \N__56952\ : std_logic;
signal \N__56949\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56943\ : std_logic;
signal \N__56940\ : std_logic;
signal \N__56939\ : std_logic;
signal \N__56936\ : std_logic;
signal \N__56935\ : std_logic;
signal \N__56932\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56926\ : std_logic;
signal \N__56923\ : std_logic;
signal \N__56920\ : std_logic;
signal \N__56915\ : std_logic;
signal \N__56912\ : std_logic;
signal \N__56909\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56901\ : std_logic;
signal \N__56898\ : std_logic;
signal \N__56895\ : std_logic;
signal \N__56894\ : std_logic;
signal \N__56893\ : std_logic;
signal \N__56890\ : std_logic;
signal \N__56887\ : std_logic;
signal \N__56884\ : std_logic;
signal \N__56881\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56868\ : std_logic;
signal \N__56865\ : std_logic;
signal \N__56862\ : std_logic;
signal \N__56859\ : std_logic;
signal \N__56856\ : std_logic;
signal \N__56853\ : std_logic;
signal \N__56850\ : std_logic;
signal \N__56849\ : std_logic;
signal \N__56848\ : std_logic;
signal \N__56841\ : std_logic;
signal \N__56838\ : std_logic;
signal \N__56835\ : std_logic;
signal \N__56832\ : std_logic;
signal \N__56829\ : std_logic;
signal \N__56826\ : std_logic;
signal \N__56823\ : std_logic;
signal \N__56822\ : std_logic;
signal \N__56819\ : std_logic;
signal \N__56816\ : std_logic;
signal \N__56815\ : std_logic;
signal \N__56812\ : std_logic;
signal \N__56809\ : std_logic;
signal \N__56806\ : std_logic;
signal \N__56803\ : std_logic;
signal \N__56800\ : std_logic;
signal \N__56797\ : std_logic;
signal \N__56794\ : std_logic;
signal \N__56787\ : std_logic;
signal \N__56784\ : std_logic;
signal \N__56781\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56775\ : std_logic;
signal \N__56774\ : std_logic;
signal \N__56773\ : std_logic;
signal \N__56770\ : std_logic;
signal \N__56765\ : std_logic;
signal \N__56762\ : std_logic;
signal \N__56759\ : std_logic;
signal \N__56756\ : std_logic;
signal \N__56753\ : std_logic;
signal \N__56750\ : std_logic;
signal \N__56747\ : std_logic;
signal \N__56744\ : std_logic;
signal \N__56741\ : std_logic;
signal \N__56736\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56730\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56724\ : std_logic;
signal \N__56723\ : std_logic;
signal \N__56720\ : std_logic;
signal \N__56717\ : std_logic;
signal \N__56714\ : std_logic;
signal \N__56711\ : std_logic;
signal \N__56710\ : std_logic;
signal \N__56705\ : std_logic;
signal \N__56702\ : std_logic;
signal \N__56699\ : std_logic;
signal \N__56696\ : std_logic;
signal \N__56693\ : std_logic;
signal \N__56690\ : std_logic;
signal \N__56687\ : std_logic;
signal \N__56682\ : std_logic;
signal \N__56679\ : std_logic;
signal \N__56676\ : std_logic;
signal \N__56673\ : std_logic;
signal \N__56672\ : std_logic;
signal \N__56671\ : std_logic;
signal \N__56664\ : std_logic;
signal \N__56661\ : std_logic;
signal \N__56658\ : std_logic;
signal \N__56655\ : std_logic;
signal \N__56652\ : std_logic;
signal \N__56649\ : std_logic;
signal \N__56648\ : std_logic;
signal \N__56647\ : std_logic;
signal \N__56640\ : std_logic;
signal \N__56637\ : std_logic;
signal \N__56634\ : std_logic;
signal \N__56631\ : std_logic;
signal \N__56628\ : std_logic;
signal \N__56627\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56619\ : std_logic;
signal \N__56616\ : std_logic;
signal \N__56613\ : std_logic;
signal \N__56610\ : std_logic;
signal \N__56609\ : std_logic;
signal \N__56608\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56604\ : std_logic;
signal \N__56603\ : std_logic;
signal \N__56600\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56597\ : std_logic;
signal \N__56594\ : std_logic;
signal \N__56593\ : std_logic;
signal \N__56592\ : std_logic;
signal \N__56589\ : std_logic;
signal \N__56586\ : std_logic;
signal \N__56583\ : std_logic;
signal \N__56580\ : std_logic;
signal \N__56577\ : std_logic;
signal \N__56574\ : std_logic;
signal \N__56571\ : std_logic;
signal \N__56568\ : std_logic;
signal \N__56565\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56561\ : std_logic;
signal \N__56558\ : std_logic;
signal \N__56553\ : std_logic;
signal \N__56544\ : std_logic;
signal \N__56541\ : std_logic;
signal \N__56538\ : std_logic;
signal \N__56535\ : std_logic;
signal \N__56532\ : std_logic;
signal \N__56529\ : std_logic;
signal \N__56522\ : std_logic;
signal \N__56515\ : std_logic;
signal \N__56508\ : std_logic;
signal \N__56507\ : std_logic;
signal \N__56506\ : std_logic;
signal \N__56503\ : std_logic;
signal \N__56500\ : std_logic;
signal \N__56497\ : std_logic;
signal \N__56494\ : std_logic;
signal \N__56491\ : std_logic;
signal \N__56488\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56486\ : std_logic;
signal \N__56483\ : std_logic;
signal \N__56480\ : std_logic;
signal \N__56479\ : std_logic;
signal \N__56476\ : std_logic;
signal \N__56473\ : std_logic;
signal \N__56470\ : std_logic;
signal \N__56467\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56465\ : std_logic;
signal \N__56464\ : std_logic;
signal \N__56461\ : std_logic;
signal \N__56458\ : std_logic;
signal \N__56455\ : std_logic;
signal \N__56454\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56448\ : std_logic;
signal \N__56445\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56437\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56433\ : std_logic;
signal \N__56428\ : std_logic;
signal \N__56425\ : std_logic;
signal \N__56422\ : std_logic;
signal \N__56417\ : std_logic;
signal \N__56412\ : std_logic;
signal \N__56409\ : std_logic;
signal \N__56406\ : std_logic;
signal \N__56403\ : std_logic;
signal \N__56400\ : std_logic;
signal \N__56397\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56389\ : std_logic;
signal \N__56388\ : std_logic;
signal \N__56385\ : std_logic;
signal \N__56384\ : std_logic;
signal \N__56381\ : std_logic;
signal \N__56378\ : std_logic;
signal \N__56375\ : std_logic;
signal \N__56368\ : std_logic;
signal \N__56363\ : std_logic;
signal \N__56360\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56334\ : std_logic;
signal \N__56331\ : std_logic;
signal \N__56328\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56324\ : std_logic;
signal \N__56321\ : std_logic;
signal \N__56318\ : std_logic;
signal \N__56313\ : std_logic;
signal \N__56312\ : std_logic;
signal \N__56311\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56305\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56295\ : std_logic;
signal \N__56292\ : std_logic;
signal \N__56289\ : std_logic;
signal \N__56286\ : std_logic;
signal \N__56285\ : std_logic;
signal \N__56284\ : std_logic;
signal \N__56279\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56275\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56270\ : std_logic;
signal \N__56267\ : std_logic;
signal \N__56266\ : std_logic;
signal \N__56263\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56257\ : std_logic;
signal \N__56252\ : std_logic;
signal \N__56249\ : std_logic;
signal \N__56246\ : std_logic;
signal \N__56243\ : std_logic;
signal \N__56242\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56221\ : std_logic;
signal \N__56220\ : std_logic;
signal \N__56217\ : std_logic;
signal \N__56214\ : std_logic;
signal \N__56211\ : std_logic;
signal \N__56208\ : std_logic;
signal \N__56203\ : std_logic;
signal \N__56200\ : std_logic;
signal \N__56197\ : std_logic;
signal \N__56194\ : std_logic;
signal \N__56191\ : std_logic;
signal \N__56186\ : std_logic;
signal \N__56183\ : std_logic;
signal \N__56174\ : std_logic;
signal \N__56163\ : std_logic;
signal \N__56160\ : std_logic;
signal \N__56157\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56153\ : std_logic;
signal \N__56150\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56142\ : std_logic;
signal \N__56141\ : std_logic;
signal \N__56140\ : std_logic;
signal \N__56139\ : std_logic;
signal \N__56136\ : std_logic;
signal \N__56133\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56129\ : std_logic;
signal \N__56126\ : std_logic;
signal \N__56125\ : std_logic;
signal \N__56124\ : std_logic;
signal \N__56121\ : std_logic;
signal \N__56118\ : std_logic;
signal \N__56115\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56111\ : std_logic;
signal \N__56110\ : std_logic;
signal \N__56107\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56105\ : std_logic;
signal \N__56102\ : std_logic;
signal \N__56099\ : std_logic;
signal \N__56096\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56090\ : std_logic;
signal \N__56087\ : std_logic;
signal \N__56084\ : std_logic;
signal \N__56081\ : std_logic;
signal \N__56078\ : std_logic;
signal \N__56075\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56073\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56067\ : std_logic;
signal \N__56064\ : std_logic;
signal \N__56061\ : std_logic;
signal \N__56058\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56046\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56034\ : std_logic;
signal \N__56031\ : std_logic;
signal \N__56028\ : std_logic;
signal \N__56025\ : std_logic;
signal \N__56020\ : std_logic;
signal \N__56017\ : std_logic;
signal \N__56016\ : std_logic;
signal \N__56013\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56002\ : std_logic;
signal \N__56001\ : std_logic;
signal \N__55998\ : std_logic;
signal \N__55995\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55983\ : std_logic;
signal \N__55980\ : std_logic;
signal \N__55971\ : std_logic;
signal \N__55968\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55947\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55943\ : std_logic;
signal \N__55940\ : std_logic;
signal \N__55937\ : std_logic;
signal \N__55932\ : std_logic;
signal \N__55931\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55927\ : std_logic;
signal \N__55926\ : std_logic;
signal \N__55923\ : std_logic;
signal \N__55922\ : std_logic;
signal \N__55919\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55913\ : std_logic;
signal \N__55910\ : std_logic;
signal \N__55907\ : std_logic;
signal \N__55904\ : std_logic;
signal \N__55903\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55899\ : std_logic;
signal \N__55898\ : std_logic;
signal \N__55895\ : std_logic;
signal \N__55892\ : std_logic;
signal \N__55889\ : std_logic;
signal \N__55886\ : std_logic;
signal \N__55883\ : std_logic;
signal \N__55880\ : std_logic;
signal \N__55877\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55867\ : std_logic;
signal \N__55864\ : std_logic;
signal \N__55859\ : std_logic;
signal \N__55856\ : std_logic;
signal \N__55853\ : std_logic;
signal \N__55850\ : std_logic;
signal \N__55847\ : std_logic;
signal \N__55846\ : std_logic;
signal \N__55845\ : std_logic;
signal \N__55842\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55836\ : std_logic;
signal \N__55835\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55825\ : std_logic;
signal \N__55822\ : std_logic;
signal \N__55819\ : std_logic;
signal \N__55818\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55814\ : std_logic;
signal \N__55811\ : std_logic;
signal \N__55806\ : std_logic;
signal \N__55803\ : std_logic;
signal \N__55794\ : std_logic;
signal \N__55789\ : std_logic;
signal \N__55786\ : std_logic;
signal \N__55773\ : std_logic;
signal \N__55770\ : std_logic;
signal \N__55767\ : std_logic;
signal \N__55766\ : std_logic;
signal \N__55763\ : std_logic;
signal \N__55760\ : std_logic;
signal \N__55755\ : std_logic;
signal \N__55754\ : std_logic;
signal \N__55751\ : std_logic;
signal \N__55750\ : std_logic;
signal \N__55749\ : std_logic;
signal \N__55746\ : std_logic;
signal \N__55743\ : std_logic;
signal \N__55740\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55734\ : std_logic;
signal \N__55733\ : std_logic;
signal \N__55732\ : std_logic;
signal \N__55731\ : std_logic;
signal \N__55730\ : std_logic;
signal \N__55727\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55723\ : std_logic;
signal \N__55720\ : std_logic;
signal \N__55717\ : std_logic;
signal \N__55716\ : std_logic;
signal \N__55713\ : std_logic;
signal \N__55710\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55705\ : std_logic;
signal \N__55702\ : std_logic;
signal \N__55699\ : std_logic;
signal \N__55696\ : std_logic;
signal \N__55693\ : std_logic;
signal \N__55688\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55682\ : std_logic;
signal \N__55679\ : std_logic;
signal \N__55676\ : std_logic;
signal \N__55673\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55667\ : std_logic;
signal \N__55666\ : std_logic;
signal \N__55659\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55644\ : std_logic;
signal \N__55639\ : std_logic;
signal \N__55636\ : std_logic;
signal \N__55633\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55625\ : std_logic;
signal \N__55616\ : std_logic;
signal \N__55605\ : std_logic;
signal \N__55602\ : std_logic;
signal \N__55599\ : std_logic;
signal \N__55596\ : std_logic;
signal \N__55595\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55589\ : std_logic;
signal \N__55584\ : std_logic;
signal \N__55583\ : std_logic;
signal \N__55582\ : std_logic;
signal \N__55581\ : std_logic;
signal \N__55578\ : std_logic;
signal \N__55575\ : std_logic;
signal \N__55574\ : std_logic;
signal \N__55571\ : std_logic;
signal \N__55568\ : std_logic;
signal \N__55567\ : std_logic;
signal \N__55566\ : std_logic;
signal \N__55565\ : std_logic;
signal \N__55562\ : std_logic;
signal \N__55559\ : std_logic;
signal \N__55556\ : std_logic;
signal \N__55553\ : std_logic;
signal \N__55550\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55545\ : std_logic;
signal \N__55542\ : std_logic;
signal \N__55541\ : std_logic;
signal \N__55538\ : std_logic;
signal \N__55535\ : std_logic;
signal \N__55534\ : std_logic;
signal \N__55531\ : std_logic;
signal \N__55528\ : std_logic;
signal \N__55525\ : std_logic;
signal \N__55522\ : std_logic;
signal \N__55521\ : std_logic;
signal \N__55518\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55503\ : std_logic;
signal \N__55500\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55494\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55486\ : std_logic;
signal \N__55483\ : std_logic;
signal \N__55480\ : std_logic;
signal \N__55477\ : std_logic;
signal \N__55474\ : std_logic;
signal \N__55471\ : std_logic;
signal \N__55468\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55462\ : std_logic;
signal \N__55459\ : std_logic;
signal \N__55456\ : std_logic;
signal \N__55453\ : std_logic;
signal \N__55450\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55446\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55436\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55428\ : std_logic;
signal \N__55421\ : std_logic;
signal \N__55416\ : std_logic;
signal \N__55413\ : std_logic;
signal \N__55410\ : std_logic;
signal \N__55395\ : std_logic;
signal \N__55392\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55388\ : std_logic;
signal \N__55385\ : std_logic;
signal \N__55382\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55374\ : std_logic;
signal \N__55373\ : std_logic;
signal \N__55372\ : std_logic;
signal \N__55369\ : std_logic;
signal \N__55366\ : std_logic;
signal \N__55363\ : std_logic;
signal \N__55362\ : std_logic;
signal \N__55357\ : std_logic;
signal \N__55356\ : std_logic;
signal \N__55355\ : std_logic;
signal \N__55354\ : std_logic;
signal \N__55353\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55347\ : std_logic;
signal \N__55344\ : std_logic;
signal \N__55343\ : std_logic;
signal \N__55342\ : std_logic;
signal \N__55339\ : std_logic;
signal \N__55336\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55332\ : std_logic;
signal \N__55329\ : std_logic;
signal \N__55326\ : std_logic;
signal \N__55323\ : std_logic;
signal \N__55320\ : std_logic;
signal \N__55317\ : std_logic;
signal \N__55314\ : std_logic;
signal \N__55311\ : std_logic;
signal \N__55308\ : std_logic;
signal \N__55305\ : std_logic;
signal \N__55302\ : std_logic;
signal \N__55299\ : std_logic;
signal \N__55296\ : std_logic;
signal \N__55293\ : std_logic;
signal \N__55290\ : std_logic;
signal \N__55285\ : std_logic;
signal \N__55284\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55270\ : std_logic;
signal \N__55265\ : std_logic;
signal \N__55260\ : std_logic;
signal \N__55257\ : std_logic;
signal \N__55254\ : std_logic;
signal \N__55251\ : std_logic;
signal \N__55248\ : std_logic;
signal \N__55239\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55227\ : std_logic;
signal \N__55224\ : std_logic;
signal \N__55223\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55206\ : std_logic;
signal \N__55205\ : std_logic;
signal \N__55202\ : std_logic;
signal \N__55199\ : std_logic;
signal \N__55194\ : std_logic;
signal \N__55191\ : std_logic;
signal \N__55188\ : std_logic;
signal \N__55185\ : std_logic;
signal \N__55182\ : std_logic;
signal \N__55179\ : std_logic;
signal \N__55176\ : std_logic;
signal \N__55173\ : std_logic;
signal \N__55170\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55168\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55159\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55148\ : std_logic;
signal \N__55145\ : std_logic;
signal \N__55140\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55134\ : std_logic;
signal \N__55133\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55122\ : std_logic;
signal \N__55119\ : std_logic;
signal \N__55116\ : std_logic;
signal \N__55113\ : std_logic;
signal \N__55110\ : std_logic;
signal \N__55107\ : std_logic;
signal \N__55104\ : std_logic;
signal \N__55103\ : std_logic;
signal \N__55102\ : std_logic;
signal \N__55095\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55089\ : std_logic;
signal \N__55086\ : std_logic;
signal \N__55083\ : std_logic;
signal \N__55080\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55078\ : std_logic;
signal \N__55075\ : std_logic;
signal \N__55070\ : std_logic;
signal \N__55067\ : std_logic;
signal \N__55064\ : std_logic;
signal \N__55061\ : std_logic;
signal \N__55058\ : std_logic;
signal \N__55053\ : std_logic;
signal \N__55050\ : std_logic;
signal \N__55047\ : std_logic;
signal \N__55044\ : std_logic;
signal \N__55043\ : std_logic;
signal \N__55042\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55032\ : std_logic;
signal \N__55029\ : std_logic;
signal \N__55026\ : std_logic;
signal \N__55023\ : std_logic;
signal \N__55020\ : std_logic;
signal \N__55017\ : std_logic;
signal \N__55014\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55010\ : std_logic;
signal \N__55009\ : std_logic;
signal \N__55006\ : std_logic;
signal \N__55001\ : std_logic;
signal \N__54996\ : std_logic;
signal \N__54993\ : std_logic;
signal \N__54990\ : std_logic;
signal \N__54987\ : std_logic;
signal \N__54984\ : std_logic;
signal \N__54983\ : std_logic;
signal \N__54982\ : std_logic;
signal \N__54975\ : std_logic;
signal \N__54972\ : std_logic;
signal \N__54969\ : std_logic;
signal \N__54966\ : std_logic;
signal \N__54963\ : std_logic;
signal \N__54960\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54958\ : std_logic;
signal \N__54957\ : std_logic;
signal \N__54954\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54942\ : std_logic;
signal \N__54939\ : std_logic;
signal \N__54936\ : std_logic;
signal \N__54933\ : std_logic;
signal \N__54930\ : std_logic;
signal \N__54929\ : std_logic;
signal \N__54928\ : std_logic;
signal \N__54927\ : std_logic;
signal \N__54924\ : std_logic;
signal \N__54917\ : std_logic;
signal \N__54912\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54910\ : std_logic;
signal \N__54909\ : std_logic;
signal \N__54906\ : std_logic;
signal \N__54899\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54891\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54882\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54876\ : std_logic;
signal \N__54873\ : std_logic;
signal \N__54870\ : std_logic;
signal \N__54869\ : std_logic;
signal \N__54868\ : std_logic;
signal \N__54865\ : std_logic;
signal \N__54860\ : std_logic;
signal \N__54857\ : std_logic;
signal \N__54854\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54846\ : std_logic;
signal \N__54843\ : std_logic;
signal \N__54840\ : std_logic;
signal \N__54837\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54832\ : std_logic;
signal \N__54827\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54819\ : std_logic;
signal \N__54816\ : std_logic;
signal \N__54813\ : std_logic;
signal \N__54812\ : std_logic;
signal \N__54809\ : std_logic;
signal \N__54808\ : std_logic;
signal \N__54805\ : std_logic;
signal \N__54802\ : std_logic;
signal \N__54799\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54786\ : std_logic;
signal \N__54783\ : std_logic;
signal \N__54780\ : std_logic;
signal \N__54777\ : std_logic;
signal \N__54776\ : std_logic;
signal \N__54775\ : std_logic;
signal \N__54768\ : std_logic;
signal \N__54765\ : std_logic;
signal \N__54762\ : std_logic;
signal \N__54759\ : std_logic;
signal \N__54756\ : std_logic;
signal \N__54753\ : std_logic;
signal \N__54752\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54748\ : std_logic;
signal \N__54743\ : std_logic;
signal \N__54740\ : std_logic;
signal \N__54737\ : std_logic;
signal \N__54734\ : std_logic;
signal \N__54731\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54725\ : std_logic;
signal \N__54720\ : std_logic;
signal \N__54717\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54710\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54699\ : std_logic;
signal \N__54696\ : std_logic;
signal \N__54693\ : std_logic;
signal \N__54690\ : std_logic;
signal \N__54687\ : std_logic;
signal \N__54684\ : std_logic;
signal \N__54681\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54675\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54669\ : std_logic;
signal \N__54666\ : std_logic;
signal \N__54663\ : std_logic;
signal \N__54660\ : std_logic;
signal \N__54657\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54650\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54642\ : std_logic;
signal \N__54639\ : std_logic;
signal \N__54636\ : std_logic;
signal \N__54633\ : std_logic;
signal \N__54630\ : std_logic;
signal \N__54629\ : std_logic;
signal \N__54626\ : std_logic;
signal \N__54623\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54615\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54606\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54597\ : std_logic;
signal \N__54594\ : std_logic;
signal \N__54591\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54579\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54570\ : std_logic;
signal \N__54569\ : std_logic;
signal \N__54568\ : std_logic;
signal \N__54567\ : std_logic;
signal \N__54564\ : std_logic;
signal \N__54557\ : std_logic;
signal \N__54552\ : std_logic;
signal \N__54549\ : std_logic;
signal \N__54546\ : std_logic;
signal \N__54543\ : std_logic;
signal \N__54540\ : std_logic;
signal \N__54537\ : std_logic;
signal \N__54536\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54532\ : std_logic;
signal \N__54527\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54516\ : std_logic;
signal \N__54513\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54498\ : std_logic;
signal \N__54495\ : std_logic;
signal \N__54494\ : std_logic;
signal \N__54493\ : std_logic;
signal \N__54490\ : std_logic;
signal \N__54489\ : std_logic;
signal \N__54482\ : std_logic;
signal \N__54479\ : std_logic;
signal \N__54476\ : std_logic;
signal \N__54471\ : std_logic;
signal \N__54468\ : std_logic;
signal \N__54465\ : std_logic;
signal \N__54462\ : std_logic;
signal \N__54459\ : std_logic;
signal \N__54458\ : std_logic;
signal \N__54455\ : std_logic;
signal \N__54452\ : std_logic;
signal \N__54447\ : std_logic;
signal \N__54444\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54438\ : std_logic;
signal \N__54435\ : std_logic;
signal \N__54432\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54428\ : std_logic;
signal \N__54425\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54411\ : std_logic;
signal \N__54408\ : std_logic;
signal \N__54405\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54398\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54392\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54384\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54378\ : std_logic;
signal \N__54377\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54371\ : std_logic;
signal \N__54366\ : std_logic;
signal \N__54363\ : std_logic;
signal \N__54360\ : std_logic;
signal \N__54357\ : std_logic;
signal \N__54354\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54348\ : std_logic;
signal \N__54347\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54340\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54334\ : std_logic;
signal \N__54327\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54321\ : std_logic;
signal \N__54318\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54314\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54305\ : std_logic;
signal \N__54302\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54294\ : std_logic;
signal \N__54291\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54282\ : std_logic;
signal \N__54279\ : std_logic;
signal \N__54278\ : std_logic;
signal \N__54273\ : std_logic;
signal \N__54270\ : std_logic;
signal \N__54267\ : std_logic;
signal \N__54264\ : std_logic;
signal \N__54261\ : std_logic;
signal \N__54258\ : std_logic;
signal \N__54257\ : std_logic;
signal \N__54252\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54243\ : std_logic;
signal \N__54240\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54234\ : std_logic;
signal \N__54231\ : std_logic;
signal \N__54228\ : std_logic;
signal \N__54225\ : std_logic;
signal \N__54222\ : std_logic;
signal \N__54219\ : std_logic;
signal \N__54218\ : std_logic;
signal \N__54213\ : std_logic;
signal \N__54210\ : std_logic;
signal \N__54207\ : std_logic;
signal \N__54204\ : std_logic;
signal \N__54201\ : std_logic;
signal \N__54198\ : std_logic;
signal \N__54197\ : std_logic;
signal \N__54192\ : std_logic;
signal \N__54189\ : std_logic;
signal \N__54186\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54180\ : std_logic;
signal \N__54179\ : std_logic;
signal \N__54174\ : std_logic;
signal \N__54171\ : std_logic;
signal \N__54168\ : std_logic;
signal \N__54165\ : std_logic;
signal \N__54162\ : std_logic;
signal \N__54159\ : std_logic;
signal \N__54156\ : std_logic;
signal \N__54153\ : std_logic;
signal \N__54152\ : std_logic;
signal \N__54147\ : std_logic;
signal \N__54144\ : std_logic;
signal \N__54141\ : std_logic;
signal \N__54140\ : std_logic;
signal \N__54139\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54133\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54123\ : std_logic;
signal \N__54122\ : std_logic;
signal \N__54121\ : std_logic;
signal \N__54118\ : std_logic;
signal \N__54113\ : std_logic;
signal \N__54110\ : std_logic;
signal \N__54107\ : std_logic;
signal \N__54102\ : std_logic;
signal \N__54099\ : std_logic;
signal \N__54096\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54094\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54078\ : std_logic;
signal \N__54077\ : std_logic;
signal \N__54072\ : std_logic;
signal \N__54069\ : std_logic;
signal \N__54066\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54057\ : std_logic;
signal \N__54054\ : std_logic;
signal \N__54053\ : std_logic;
signal \N__54052\ : std_logic;
signal \N__54049\ : std_logic;
signal \N__54044\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54035\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54030\ : std_logic;
signal \N__54029\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54010\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__53999\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53991\ : std_logic;
signal \N__53990\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53984\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53982\ : std_logic;
signal \N__53981\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53978\ : std_logic;
signal \N__53975\ : std_logic;
signal \N__53974\ : std_logic;
signal \N__53971\ : std_logic;
signal \N__53962\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53954\ : std_logic;
signal \N__53951\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53936\ : std_logic;
signal \N__53933\ : std_logic;
signal \N__53928\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53919\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53915\ : std_logic;
signal \N__53912\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53891\ : std_logic;
signal \N__53888\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53882\ : std_logic;
signal \N__53879\ : std_logic;
signal \N__53876\ : std_logic;
signal \N__53873\ : std_logic;
signal \N__53870\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53850\ : std_logic;
signal \N__53849\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53840\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53826\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53820\ : std_logic;
signal \N__53819\ : std_logic;
signal \N__53816\ : std_logic;
signal \N__53815\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53803\ : std_logic;
signal \N__53796\ : std_logic;
signal \N__53795\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53784\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53776\ : std_logic;
signal \N__53773\ : std_logic;
signal \N__53770\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53760\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53747\ : std_logic;
signal \N__53744\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53738\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53730\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53724\ : std_logic;
signal \N__53721\ : std_logic;
signal \N__53718\ : std_logic;
signal \N__53715\ : std_logic;
signal \N__53712\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53706\ : std_logic;
signal \N__53703\ : std_logic;
signal \N__53700\ : std_logic;
signal \N__53697\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53688\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53678\ : std_logic;
signal \N__53673\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53663\ : std_logic;
signal \N__53658\ : std_logic;
signal \N__53655\ : std_logic;
signal \N__53652\ : std_logic;
signal \N__53649\ : std_logic;
signal \N__53646\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53644\ : std_logic;
signal \N__53639\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53628\ : std_logic;
signal \N__53625\ : std_logic;
signal \N__53624\ : std_logic;
signal \N__53623\ : std_logic;
signal \N__53620\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53610\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53604\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53600\ : std_logic;
signal \N__53599\ : std_logic;
signal \N__53596\ : std_logic;
signal \N__53591\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53582\ : std_logic;
signal \N__53577\ : std_logic;
signal \N__53574\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53567\ : std_logic;
signal \N__53564\ : std_logic;
signal \N__53561\ : std_logic;
signal \N__53556\ : std_logic;
signal \N__53553\ : std_logic;
signal \N__53550\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53544\ : std_logic;
signal \N__53541\ : std_logic;
signal \N__53538\ : std_logic;
signal \N__53537\ : std_logic;
signal \N__53534\ : std_logic;
signal \N__53531\ : std_logic;
signal \N__53528\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53514\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53509\ : std_logic;
signal \N__53506\ : std_logic;
signal \N__53503\ : std_logic;
signal \N__53500\ : std_logic;
signal \N__53497\ : std_logic;
signal \N__53494\ : std_logic;
signal \N__53491\ : std_logic;
signal \N__53486\ : std_logic;
signal \N__53483\ : std_logic;
signal \N__53480\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53472\ : std_logic;
signal \N__53469\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53463\ : std_logic;
signal \N__53460\ : std_logic;
signal \N__53459\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53451\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53432\ : std_logic;
signal \N__53431\ : std_logic;
signal \N__53428\ : std_logic;
signal \N__53425\ : std_logic;
signal \N__53420\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53412\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53402\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53398\ : std_logic;
signal \N__53397\ : std_logic;
signal \N__53396\ : std_logic;
signal \N__53393\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53386\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53380\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53376\ : std_logic;
signal \N__53371\ : std_logic;
signal \N__53370\ : std_logic;
signal \N__53367\ : std_logic;
signal \N__53364\ : std_logic;
signal \N__53361\ : std_logic;
signal \N__53360\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53354\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53337\ : std_logic;
signal \N__53334\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53324\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53315\ : std_logic;
signal \N__53312\ : std_logic;
signal \N__53309\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53297\ : std_logic;
signal \N__53294\ : std_logic;
signal \N__53291\ : std_logic;
signal \N__53288\ : std_logic;
signal \N__53283\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53266\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53249\ : std_logic;
signal \N__53246\ : std_logic;
signal \N__53243\ : std_logic;
signal \N__53240\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53228\ : std_logic;
signal \N__53225\ : std_logic;
signal \N__53224\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53215\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53211\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53205\ : std_logic;
signal \N__53204\ : std_logic;
signal \N__53201\ : std_logic;
signal \N__53198\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53189\ : std_logic;
signal \N__53186\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53178\ : std_logic;
signal \N__53173\ : std_logic;
signal \N__53170\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53164\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53156\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53133\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53126\ : std_logic;
signal \N__53123\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53117\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53111\ : std_logic;
signal \N__53108\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53102\ : std_logic;
signal \N__53099\ : std_logic;
signal \N__53094\ : std_logic;
signal \N__53091\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53081\ : std_logic;
signal \N__53080\ : std_logic;
signal \N__53073\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53054\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53040\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53021\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53004\ : std_logic;
signal \N__53001\ : std_logic;
signal \N__52998\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52985\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52974\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52961\ : std_logic;
signal \N__52956\ : std_logic;
signal \N__52955\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52947\ : std_logic;
signal \N__52944\ : std_logic;
signal \N__52941\ : std_logic;
signal \N__52938\ : std_logic;
signal \N__52935\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52923\ : std_logic;
signal \N__52920\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52914\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52904\ : std_logic;
signal \N__52899\ : std_logic;
signal \N__52896\ : std_logic;
signal \N__52893\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52878\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52865\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52839\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52821\ : std_logic;
signal \N__52820\ : std_logic;
signal \N__52815\ : std_logic;
signal \N__52812\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52806\ : std_logic;
signal \N__52803\ : std_logic;
signal \N__52800\ : std_logic;
signal \N__52797\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52776\ : std_logic;
signal \N__52773\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52766\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52760\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52736\ : std_logic;
signal \N__52733\ : std_logic;
signal \N__52730\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52724\ : std_logic;
signal \N__52721\ : std_logic;
signal \N__52718\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52709\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52705\ : std_logic;
signal \N__52702\ : std_logic;
signal \N__52699\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52693\ : std_logic;
signal \N__52690\ : std_logic;
signal \N__52687\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52680\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52676\ : std_logic;
signal \N__52673\ : std_logic;
signal \N__52670\ : std_logic;
signal \N__52667\ : std_logic;
signal \N__52664\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52656\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52643\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52614\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52608\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52598\ : std_logic;
signal \N__52597\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52565\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52529\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52502\ : std_logic;
signal \N__52501\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52488\ : std_logic;
signal \N__52485\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52472\ : std_logic;
signal \N__52469\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52467\ : std_logic;
signal \N__52464\ : std_logic;
signal \N__52461\ : std_logic;
signal \N__52458\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52403\ : std_logic;
signal \N__52400\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52379\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52374\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52368\ : std_logic;
signal \N__52365\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52341\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52324\ : std_logic;
signal \N__52317\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52308\ : std_logic;
signal \N__52307\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52295\ : std_logic;
signal \N__52292\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52274\ : std_logic;
signal \N__52273\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52259\ : std_logic;
signal \N__52256\ : std_logic;
signal \N__52253\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52197\ : std_logic;
signal \N__52194\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52185\ : std_logic;
signal \N__52182\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52173\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52166\ : std_logic;
signal \N__52163\ : std_logic;
signal \N__52160\ : std_logic;
signal \N__52157\ : std_logic;
signal \N__52154\ : std_logic;
signal \N__52149\ : std_logic;
signal \N__52146\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52128\ : std_logic;
signal \N__52127\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52115\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52101\ : std_logic;
signal \N__52098\ : std_logic;
signal \N__52095\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52082\ : std_logic;
signal \N__52079\ : std_logic;
signal \N__52076\ : std_logic;
signal \N__52071\ : std_logic;
signal \N__52068\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52056\ : std_logic;
signal \N__52053\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52032\ : std_logic;
signal \N__52029\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52022\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52011\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51990\ : std_logic;
signal \N__51987\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51981\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51977\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51968\ : std_logic;
signal \N__51965\ : std_logic;
signal \N__51962\ : std_logic;
signal \N__51959\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51941\ : std_logic;
signal \N__51938\ : std_logic;
signal \N__51935\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51929\ : std_logic;
signal \N__51926\ : std_logic;
signal \N__51923\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51912\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51902\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51876\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51869\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51834\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51806\ : std_logic;
signal \N__51803\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51780\ : std_logic;
signal \N__51779\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51737\ : std_logic;
signal \N__51734\ : std_logic;
signal \N__51731\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51701\ : std_logic;
signal \N__51698\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51692\ : std_logic;
signal \N__51689\ : std_logic;
signal \N__51686\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51662\ : std_logic;
signal \N__51659\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51627\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51621\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51611\ : std_logic;
signal \N__51608\ : std_logic;
signal \N__51603\ : std_logic;
signal \N__51600\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51591\ : std_logic;
signal \N__51588\ : std_logic;
signal \N__51585\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51576\ : std_logic;
signal \N__51575\ : std_logic;
signal \N__51572\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51558\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51549\ : std_logic;
signal \N__51548\ : std_logic;
signal \N__51545\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51537\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51524\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51506\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51500\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51468\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51462\ : std_logic;
signal \N__51459\ : std_logic;
signal \N__51456\ : std_logic;
signal \N__51453\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51427\ : std_logic;
signal \N__51426\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51416\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51404\ : std_logic;
signal \N__51401\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51381\ : std_logic;
signal \N__51378\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51366\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51350\ : std_logic;
signal \N__51347\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51334\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51318\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51249\ : std_logic;
signal \N__51246\ : std_logic;
signal \N__51243\ : std_logic;
signal \N__51240\ : std_logic;
signal \N__51237\ : std_logic;
signal \N__51234\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51215\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51195\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51180\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51173\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51162\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51155\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51147\ : std_logic;
signal \N__51144\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51138\ : std_logic;
signal \N__51135\ : std_logic;
signal \N__51132\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51116\ : std_logic;
signal \N__51113\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51099\ : std_logic;
signal \N__51096\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51078\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51072\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51046\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51023\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50997\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50992\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50916\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50838\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50832\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50738\ : std_logic;
signal \N__50735\ : std_logic;
signal \N__50732\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50728\ : std_logic;
signal \N__50725\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50700\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50683\ : std_logic;
signal \N__50680\ : std_logic;
signal \N__50677\ : std_logic;
signal \N__50674\ : std_logic;
signal \N__50671\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50608\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50519\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50193\ : std_logic;
signal \N__50190\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50064\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50024\ : std_logic;
signal \N__50021\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49725\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49556\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49376\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45325\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \Pc2drone_pll_inst.clk_system_pll\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pid_alt.O_3_10\ : std_logic;
signal \pid_alt.O_3_5\ : std_logic;
signal \pid_alt.O_3_14\ : std_logic;
signal \pid_alt.O_3_15\ : std_logic;
signal \pid_alt.O_3_16\ : std_logic;
signal \pid_alt.O_3_17\ : std_logic;
signal \pid_alt.O_3_18\ : std_logic;
signal \pid_alt.O_3_19\ : std_logic;
signal \pid_alt.O_3_20\ : std_logic;
signal \pid_alt.O_3_21\ : std_logic;
signal \pid_alt.O_3_22\ : std_logic;
signal \pid_alt.O_3_23\ : std_logic;
signal \pid_alt.O_3_6\ : std_logic;
signal \pid_alt.O_3_24\ : std_logic;
signal \pid_alt.O_3_7\ : std_logic;
signal \pid_alt.O_3_9\ : std_logic;
signal alt_kd_7 : std_logic;
signal alt_kd_2 : std_logic;
signal alt_kd_1 : std_logic;
signal alt_kd_5 : std_logic;
signal alt_ki_6 : std_logic;
signal alt_ki_7 : std_logic;
signal alt_ki_1 : std_logic;
signal alt_ki_3 : std_logic;
signal alt_ki_4 : std_logic;
signal alt_ki_5 : std_logic;
signal \pid_alt.O_4_9\ : std_logic;
signal \pid_alt.O_4_24\ : std_logic;
signal \pid_alt.O_4_23\ : std_logic;
signal \pid_alt.O_4_22\ : std_logic;
signal \pid_alt.O_4_10\ : std_logic;
signal \pid_alt.O_4_14\ : std_logic;
signal \pid_alt.O_4_11\ : std_logic;
signal \pid_alt.O_4_17\ : std_logic;
signal \pid_alt.O_4_16\ : std_logic;
signal \pid_alt.O_4_20\ : std_logic;
signal \pid_alt.O_4_18\ : std_logic;
signal \pid_alt.O_4_19\ : std_logic;
signal \pid_alt.O_4_6\ : std_logic;
signal \pid_alt.O_4_21\ : std_logic;
signal \pid_alt.O_4_13\ : std_logic;
signal \pid_alt.O_4_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_\ : std_logic;
signal \pid_alt.N_1666_i_1\ : std_logic;
signal \pid_alt.N_3_1\ : std_logic;
signal \pid_alt.N_1668_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2\ : std_logic;
signal \pid_alt.N_1674_0_cascade_\ : std_logic;
signal \pid_alt.N_1666_i_0\ : std_logic;
signal \pid_alt.N_3_0\ : std_logic;
signal \pid_alt.N_1668_0\ : std_logic;
signal \pid_alt.N_5\ : std_logic;
signal \pid_alt.N_1672_0\ : std_logic;
signal \pid_front.O_0_16\ : std_logic;
signal \pid_front.O_0_17\ : std_logic;
signal \pid_front.O_0_18\ : std_logic;
signal \pid_front.O_0_19\ : std_logic;
signal \pid_front.O_0_12\ : std_logic;
signal \pid_front.O_0_7\ : std_logic;
signal \pid_front.O_0_22\ : std_logic;
signal \pid_front.O_0_23\ : std_logic;
signal \pid_front.O_0_24\ : std_logic;
signal \pid_front.O_0_21\ : std_logic;
signal \pid_front.O_0_20\ : std_logic;
signal \pid_front.O_0_14\ : std_logic;
signal \pid_front.O_0_10\ : std_logic;
signal \pid_front.O_0_13\ : std_logic;
signal \pid_alt.O_5_6\ : std_logic;
signal \pid_alt.O_5_5\ : std_logic;
signal \pid_front.O_0_8\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8\ : std_logic;
signal \pid_alt.O_5_7\ : std_logic;
signal \pid_alt.O_5_8\ : std_logic;
signal \pid_alt.O_4_8\ : std_logic;
signal \pid_alt.O_5_11\ : std_logic;
signal \pid_alt.O_5_22\ : std_logic;
signal \pid_alt.O_5_15\ : std_logic;
signal \pid_alt.O_5_17\ : std_logic;
signal \pid_alt.O_5_20\ : std_logic;
signal \pid_alt.O_5_18\ : std_logic;
signal \pid_alt.O_5_21\ : std_logic;
signal \pid_alt.O_5_19\ : std_logic;
signal \pid_alt.O_5_14\ : std_logic;
signal \pid_alt.O_5_23\ : std_logic;
signal \pid_alt.O_5_16\ : std_logic;
signal \pid_alt.O_5_12\ : std_logic;
signal \pid_alt.O_5_13\ : std_logic;
signal \pid_alt.O_5_24\ : std_logic;
signal alt_kd_6 : std_logic;
signal alt_kd_4 : std_logic;
signal alt_kd_3 : std_logic;
signal alt_kd_0 : std_logic;
signal alt_ki_0 : std_logic;
signal alt_ki_2 : std_logic;
signal \Commands_frame_decoder.state_RNIQRI31Z0Z_10\ : std_logic;
signal \pid_alt.g0_4_0\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\ : std_logic;
signal \pid_alt.O_4_5\ : std_logic;
signal \pid_alt.O_3_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_5\ : std_logic;
signal \pid_alt.error_d_regZ0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_6\ : std_logic;
signal \pid_alt.error_d_regZ0Z_6\ : std_logic;
signal \pid_alt.error_p_regZ0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_2\ : std_logic;
signal \pid_alt.error_d_regZ0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_\ : std_logic;
signal \pid_alt.O_5_4\ : std_logic;
signal \pid_alt.error_p_regZ0Z_0\ : std_logic;
signal \pid_alt.N_1666_i\ : std_logic;
signal \pid_alt.error_p_regZ0Z_1\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_1\ : std_logic;
signal \pid_alt.N_1666_i_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_1\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_axb_2_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11\ : std_logic;
signal \pid_alt.error_d_regZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\ : std_logic;
signal \pid_alt.error_d_regZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_12\ : std_logic;
signal \pid_alt.error_p_regZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\ : std_logic;
signal \pid_alt.error_p_regZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_18\ : std_logic;
signal \pid_alt.error_d_regZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\ : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal \pid_alt.error_1\ : std_logic;
signal \pid_alt.error_cry_0\ : std_logic;
signal \pid_alt.error_2\ : std_logic;
signal \pid_alt.error_cry_1\ : std_logic;
signal \pid_alt.error_3\ : std_logic;
signal \pid_alt.error_cry_2\ : std_logic;
signal alt_command_0 : std_logic;
signal \pid_alt.error_4\ : std_logic;
signal \pid_alt.error_cry_3\ : std_logic;
signal alt_command_1 : std_logic;
signal \pid_alt.error_5\ : std_logic;
signal \pid_alt.error_cry_4\ : std_logic;
signal alt_command_2 : std_logic;
signal \pid_alt.error_6\ : std_logic;
signal \pid_alt.error_cry_5\ : std_logic;
signal alt_command_3 : std_logic;
signal \pid_alt.error_7\ : std_logic;
signal \pid_alt.error_cry_6\ : std_logic;
signal \pid_alt.error_cry_7\ : std_logic;
signal alt_command_4 : std_logic;
signal \pid_alt.error_8\ : std_logic;
signal \bfn_2_20_0_\ : std_logic;
signal alt_command_5 : std_logic;
signal \pid_alt.error_9\ : std_logic;
signal \pid_alt.error_cry_8\ : std_logic;
signal alt_command_6 : std_logic;
signal \pid_alt.error_10\ : std_logic;
signal \pid_alt.error_cry_9\ : std_logic;
signal alt_command_7 : std_logic;
signal \pid_alt.error_11\ : std_logic;
signal \pid_alt.error_cry_10\ : std_logic;
signal \pid_alt.error_12\ : std_logic;
signal \pid_alt.error_cry_11\ : std_logic;
signal \pid_alt.error_13\ : std_logic;
signal \pid_alt.error_cry_12\ : std_logic;
signal \pid_alt.error_14\ : std_logic;
signal \pid_alt.error_cry_13\ : std_logic;
signal \pid_alt.error_cry_14\ : std_logic;
signal \pid_alt.error_15\ : std_logic;
signal alt_kp_1 : std_logic;
signal drone_altitude_i_10 : std_logic;
signal alt_kp_0 : std_logic;
signal alt_kp_6 : std_logic;
signal \pid_alt.O_5_9\ : std_logic;
signal \pid_alt.error_p_regZ0Z_5\ : std_logic;
signal \pid_alt.O_5_10\ : std_logic;
signal \pid_alt.error_p_regZ0Z_6\ : std_logic;
signal alt_kp_7 : std_logic;
signal alt_kp_3 : std_logic;
signal \pid_alt.O_3_8\ : std_logic;
signal \Commands_frame_decoder.state_RNIRSI31Z0Z_11\ : std_logic;
signal \pid_alt.O_3_11\ : std_logic;
signal \pid_alt.O_3_12\ : std_logic;
signal \pid_alt.O_3_13\ : std_logic;
signal \pid_alt.O_4_4\ : std_logic;
signal \pid_alt.O_4_7\ : std_logic;
signal \pid_alt.O_4_15\ : std_logic;
signal \pid_alt.N_664_0_g\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8lt7_0\ : std_logic;
signal \pid_alt.error_d_regZ0Z_0\ : std_logic;
signal \pid_alt.error_p_regZ0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_3\ : std_logic;
signal \pid_alt.error_d_regZ0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\ : std_logic;
signal \pid_alt.error_p_regZ0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \pid_alt.error_i_regZ0Z_1\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_0\ : std_logic;
signal \pid_alt.error_i_regZ0Z_2\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_1\ : std_logic;
signal \pid_alt.error_i_regZ0Z_3\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_2\ : std_logic;
signal \pid_alt.error_i_regZ0Z_4\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_3\ : std_logic;
signal \pid_alt.error_i_regZ0Z_5\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_4\ : std_logic;
signal \pid_alt.error_i_regZ0Z_6\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_5\ : std_logic;
signal \pid_alt.error_i_regZ0Z_7\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_6\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_7\ : std_logic;
signal \pid_alt.error_i_regZ0Z_8\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \pid_alt.error_i_regZ0Z_9\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_8\ : std_logic;
signal \pid_alt.error_i_regZ0Z_10\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_9\ : std_logic;
signal \pid_alt.error_i_regZ0Z_11\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_10\ : std_logic;
signal \pid_alt.error_i_regZ0Z_12\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_11\ : std_logic;
signal \pid_alt.error_i_regZ0Z_13\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_12\ : std_logic;
signal \pid_alt.error_i_regZ0Z_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_13\ : std_logic;
signal \pid_alt.error_i_regZ0Z_15\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_15\ : std_logic;
signal \pid_alt.error_i_regZ0Z_16\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \pid_alt.error_i_regZ0Z_17\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_16\ : std_logic;
signal \pid_alt.error_i_regZ0Z_18\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_17\ : std_logic;
signal \pid_alt.error_i_regZ0Z_19\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_18\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19\ : std_logic;
signal \pid_alt.error_i_regZ0Z_20\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\ : std_logic;
signal \pid_alt.un1_pid_prereg_0\ : std_logic;
signal \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_2\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_5\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_6\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_7\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_8\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_12\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_13\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_14\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_15\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_18\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_20\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_21\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_22\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_23\ : std_logic;
signal \pid_alt.error_p_regZ0Z_13\ : std_logic;
signal \pid_alt.error_d_regZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_10\ : std_logic;
signal alt_kp_2 : std_logic;
signal alt_kp_5 : std_logic;
signal \Commands_frame_decoder.stateZ0Z_2\ : std_logic;
signal \pid_alt.error_i_regZ0Z_0\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_18\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_19\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_20\ : std_logic;
signal \pid_alt.m7_e_4_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_16\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_17\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_14\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_15\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_3\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_1\ : std_logic;
signal \pid_alt.N_9_0_cascade_\ : std_logic;
signal \pid_alt.N_62_mux_cascade_\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_0\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_4\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3Z0Z_5\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_2\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_10\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_11\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_6\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_7\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_8\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_9\ : std_logic;
signal \pid_alt.m35_e_2\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11\ : std_logic;
signal \pid_alt.error_p_regZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_10\ : std_logic;
signal \pid_alt.error_d_regZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\ : std_logic;
signal drone_altitude_i_11 : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\ : std_logic;
signal \pid_alt.error_d_regZ0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_9\ : std_logic;
signal \pid_alt.error_p_regZ0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\ : std_logic;
signal \pid_alt.error_p_regZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_14\ : std_logic;
signal \pid_alt.error_d_regZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_8\ : std_logic;
signal \pid_alt.error_p_regZ0Z_8\ : std_logic;
signal \pid_alt.error_d_regZ0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\ : std_logic;
signal \pid_alt.error_d_regZ0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_7\ : std_logic;
signal \pid_alt.error_p_regZ0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\ : std_logic;
signal \pid_alt.error_d_regZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_16\ : std_logic;
signal \pid_alt.error_p_regZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\ : std_logic;
signal \pid_alt.un1_pid_prereg_236_1_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_19\ : std_logic;
signal \pid_alt.error_d_regZ0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\ : std_logic;
signal \pid_alt.error_p_regZ0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_20\ : std_logic;
signal \pid_alt.error_d_regZ0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_236_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20_cascade_\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_416_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_382\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_0_2_2\ : std_logic;
signal \Commands_frame_decoder.N_376_2\ : std_logic;
signal \Commands_frame_decoder.N_377\ : std_logic;
signal \Commands_frame_decoder.N_376_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_379\ : std_logic;
signal \Commands_frame_decoder.N_416\ : std_logic;
signal \Commands_frame_decoder.N_379_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.N_412\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_8\ : std_logic;
signal \Commands_frame_decoder.state_RNIF38SZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_9\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_3\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_2\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_7\ : std_logic;
signal \pid_alt.m21_e_0_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm7lto4\ : std_logic;
signal \pid_alt.m35_e_3\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_9\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_8\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_11\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_6\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_1\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_0\ : std_logic;
signal \pid_alt.m21_e_8_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm7lto12\ : std_logic;
signal \pid_alt.m21_e_2\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_10\ : std_logic;
signal \pid_alt.state_0_g_0\ : std_logic;
signal \pid_alt.m21_e_9\ : std_logic;
signal \pid_alt.m21_e_10\ : std_logic;
signal \pid_alt.N_9_0\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNIO7B05Z0Z_21_cascade_\ : std_logic;
signal \pid_alt.un1_reset_1_0_i_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_21\ : std_logic;
signal \pid_alt.error_i_acumm7lto13\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_13\ : std_logic;
signal \pid_alt.N_72_i_0\ : std_logic;
signal \pid_alt.un1_reset_1_cascade_\ : std_logic;
signal \pid_alt.source_pid_9_0_tz_6_cascade_\ : std_logic;
signal \pid_alt.source_pid_9_0_tz_6\ : std_logic;
signal \pid_alt.pid_preregZ0Z_2\ : std_logic;
signal \pid_alt.pid_preregZ0Z_3\ : std_logic;
signal \pid_alt.pid_preregZ0Z_1\ : std_logic;
signal \pid_alt.N_44_cascade_\ : std_logic;
signal \pid_alt.N_46\ : std_logic;
signal \pid_alt.pid_preregZ0Z_0\ : std_logic;
signal \pid_alt.N_46_cascade_\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_1_7\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_1_4\ : std_logic;
signal \pid_alt.pid_preregZ0Z_11\ : std_logic;
signal \pid_alt.pid_preregZ0Z_9\ : std_logic;
signal \pid_alt.pid_preregZ0Z_10\ : std_logic;
signal \pid_alt.pid_preregZ0Z_8\ : std_logic;
signal \pid_alt.pid_preregZ0Z_7\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_6\ : std_logic;
signal \pid_alt.N_90_cascade_\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_0_2\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_\ : std_logic;
signal \pid_alt.N_43\ : std_logic;
signal \pid_alt.N_48\ : std_logic;
signal \pid_alt.pid_preregZ0Z_15\ : std_logic;
signal \pid_alt.pid_preregZ0Z_23\ : std_logic;
signal \pid_alt.pid_preregZ0Z_21\ : std_logic;
signal \pid_alt.pid_preregZ0Z_18\ : std_logic;
signal \pid_alt.pid_preregZ0Z_22\ : std_logic;
signal \pid_alt.pid_preregZ0Z_20\ : std_logic;
signal \pid_alt.pid_preregZ0Z_17\ : std_logic;
signal \pid_alt.pid_preregZ0Z_19\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_2_6\ : std_logic;
signal \pid_alt.pid_preregZ0Z_14\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_16\ : std_logic;
signal \pid_alt.N_90\ : std_logic;
signal \pid_alt.N_305_cascade_\ : std_logic;
signal \pid_alt.source_pid_9_0_0_4_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_4\ : std_logic;
signal \pid_alt.N_44\ : std_logic;
signal \pid_alt.pid_preregZ0Z_5\ : std_logic;
signal \pid_alt.pid_preregZ0Z_13\ : std_logic;
signal \pid_alt.pid_preregZ0Z_24\ : std_logic;
signal \pid_alt.N_305\ : std_logic;
signal \pid_alt.pid_preregZ0Z_12\ : std_logic;
signal \pid_alt.N_72_i_1\ : std_logic;
signal \pid_alt.un1_reset_0_i\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_17\ : std_logic;
signal \pid_alt.error_p_regZ0Z_17\ : std_logic;
signal \pid_alt.error_d_regZ0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_4\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_1\ : std_logic;
signal \uart_pc.timer_CountZ1Z_1\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_3\ : std_logic;
signal \uart_pc.N_144_1_cascade_\ : std_logic;
signal \uart_pc.un1_state_2_0_a3_0\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_2\ : std_logic;
signal \uart_pc.timer_CountZ1Z_2\ : std_logic;
signal \uart_pc.N_126_li_cascade_\ : std_logic;
signal \uart_pc.N_143\ : std_logic;
signal \uart_pc.N_143_cascade_\ : std_logic;
signal \uart_pc.timer_CountZ0Z_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_0_2_0\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\ : std_logic;
signal \uart_pc.data_rdyc_1\ : std_logic;
signal \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_378\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_i_1_1\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\ : std_logic;
signal xy_kp_4 : std_logic;
signal \Commands_frame_decoder.stateZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_10\ : std_logic;
signal alt_kp_4 : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa\ : std_logic;
signal \pid_front.O_0_6\ : std_logic;
signal \pid_front.O_0_4\ : std_logic;
signal \pid_front.O_0_9\ : std_logic;
signal \pid_front.O_0_15\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_11\ : std_logic;
signal drone_altitude_15 : std_logic;
signal drone_altitude_i_4 : std_logic;
signal drone_altitude_i_5 : std_logic;
signal drone_altitude_i_6 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_9\ : std_logic;
signal drone_altitude_i_9 : std_logic;
signal drone_altitude_i_8 : std_logic;
signal drone_altitude_i_7 : std_logic;
signal \pid_alt.drone_altitude_i_0\ : std_logic;
signal \pid_alt.error_axbZ0Z_13\ : std_logic;
signal \pid_alt.error_axbZ0Z_14\ : std_logic;
signal \pid_alt.error_axbZ0Z_12\ : std_logic;
signal uart_input_drone_c : std_logic;
signal \uart_drone_sync.aux_0__0__0_0\ : std_logic;
signal \uart_drone_sync.aux_1__0__0_0\ : std_logic;
signal \uart_drone_sync.aux_2__0__0_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \Commands_frame_decoder.un1_state57_iZ0\ : std_logic;
signal \uart_pc.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_1\ : std_logic;
signal \uart_pc.N_126_li\ : std_logic;
signal \uart_pc.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_0\ : std_logic;
signal \uart_pc.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_pc.stateZ0Z_4\ : std_logic;
signal \uart_pc.un1_state_4_0_cascade_\ : std_logic;
signal \uart_pc.timer_CountZ0Z_4\ : std_logic;
signal \uart_pc.timer_CountZ1Z_3\ : std_logic;
signal \uart_pc.N_144_1\ : std_logic;
signal \uart_pc.N_145_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_2\ : std_logic;
signal \uart_pc_sync.aux_3__0_Z0Z_0\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_1_cascade_\ : std_logic;
signal \uart_pc.data_AuxZ1Z_0\ : std_logic;
signal \uart_pc.data_AuxZ1Z_1\ : std_logic;
signal \uart_pc.data_AuxZ1Z_2\ : std_logic;
signal \uart_pc.data_AuxZ0Z_3\ : std_logic;
signal \uart_pc.data_AuxZ0Z_4\ : std_logic;
signal \uart_pc.data_AuxZ0Z_5\ : std_logic;
signal \uart_pc.data_AuxZ0Z_6\ : std_logic;
signal \uart_pc.un1_state_2_0\ : std_logic;
signal \debug_CH2_18A_c\ : std_logic;
signal \uart_pc.data_AuxZ0Z_7\ : std_logic;
signal \uart_pc.state_RNIEAGSZ0Z_4\ : std_logic;
signal \uart_pc.stateZ0Z_3\ : std_logic;
signal \uart_pc.CO0_cascade_\ : std_logic;
signal \uart_pc.un1_state_4_0\ : std_logic;
signal \uart_pc.un1_state_7_0\ : std_logic;
signal \uart_pc.data_Auxce_0_0_4\ : std_logic;
signal \uart_pc.data_Auxce_0_5\ : std_logic;
signal \uart_pc.data_Auxce_0_6\ : std_logic;
signal \uart_pc.N_152\ : std_logic;
signal \uart_pc.data_Auxce_0_0_0\ : std_logic;
signal \uart_pc.data_Auxce_0_1\ : std_logic;
signal \uart_pc.data_Auxce_0_0_2\ : std_logic;
signal \uart_pc.bit_CountZ0Z_2\ : std_logic;
signal \uart_pc.bit_CountZ0Z_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_1\ : std_logic;
signal \uart_pc.data_Auxce_0_3\ : std_logic;
signal xy_kp_6 : std_logic;
signal xy_kp_5 : std_logic;
signal drone_altitude_0 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_4\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_5\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_6\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_7\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_8\ : std_logic;
signal drone_altitude_14 : std_logic;
signal drone_altitude_13 : std_logic;
signal drone_altitude_12 : std_logic;
signal \dron_frame_decoder_1.N_513_0\ : std_logic;
signal \pid_front.error_p_regZ0Z_9\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_9\ : std_logic;
signal \pid_front.N_1459_i\ : std_logic;
signal \pid_front.O_0_11\ : std_logic;
signal \pid_front.N_1451_i_cascade_\ : std_logic;
signal \pid_front.error_d_reg_esr_RNINKUFZ0Z_7_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_70_0\ : std_logic;
signal \pid_front.un1_pid_prereg_23\ : std_logic;
signal \pid_front.un1_pid_prereg_23_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_30_cascade_\ : std_logic;
signal \pid_front.error_p_regZ0Z_15\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_15\ : std_logic;
signal \pid_front.un1_pid_prereg_29\ : std_logic;
signal \pid_front.un1_pid_prereg_29_cascade_\ : std_logic;
signal \pid_front.error_p_regZ0Z_14\ : std_logic;
signal \pid_front.un1_pid_prereg_24\ : std_logic;
signal \pid_front.state_0_0\ : std_logic;
signal uart_input_pc_c : std_logic;
signal \uart_pc_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \uart_drone_sync.aux_3__0__0_0\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxa_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxa\ : std_logic;
signal \uart_pc_sync.aux_1__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \Commands_frame_decoder.WDT_RNII19A1Z0Z_4_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT8lto15_N_5L7_1\ : std_logic;
signal \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \Commands_frame_decoder.WDT8_0\ : std_logic;
signal \uart_drone.N_126_li_cascade_\ : std_logic;
signal \uart_drone.N_143_cascade_\ : std_logic;
signal \uart_drone.timer_CountZ1Z_1\ : std_logic;
signal \uart_drone.timer_CountZ0Z_0\ : std_logic;
signal \uart_drone.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_3\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_4\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_2\ : std_logic;
signal \uart_drone.N_143\ : std_logic;
signal \uart_drone.timer_CountZ1Z_2\ : std_logic;
signal \Commands_frame_decoder.preinitZ0\ : std_logic;
signal \uart_drone.data_rdyc_1\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_0\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.count_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_13\ : std_logic;
signal uart_pc_data_rdy : std_logic;
signal \dron_frame_decoder_1.state_ns_0_a3_0_1Z0Z_1_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_220\ : std_logic;
signal \dron_frame_decoder_1.N_220_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_224\ : std_logic;
signal \dron_frame_decoder_1.N_198_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_200\ : std_logic;
signal xy_kp_0 : std_logic;
signal xy_kp_1 : std_logic;
signal xy_kp_2 : std_logic;
signal xy_kp_3 : std_logic;
signal xy_kp_7 : std_logic;
signal \Commands_frame_decoder.state_RNIG48SZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_0\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_a2_0_0_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\ : std_logic;
signal \dron_frame_decoder_1.state_RNI6P6KZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_9\ : std_logic;
signal drone_altitude_1 : std_logic;
signal \pid_alt.error_axbZ0Z_1\ : std_logic;
signal \pid_front.error_p_regZ0Z_8\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_8\ : std_logic;
signal \pid_front.un1_pid_prereg_80_0\ : std_logic;
signal \pid_front.N_1455_i\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_57_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_48_cascade_\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_19\ : std_logic;
signal \pid_front.error_p_regZ0Z_19\ : std_logic;
signal \pid_front.un1_pid_prereg_56\ : std_logic;
signal \pid_front.un1_pid_prereg_56_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_48\ : std_logic;
signal \pid_front.N_1471_i\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIA93NZ0Z_12\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_12\ : std_logic;
signal \pid_front.error_p_regZ0Z_12\ : std_logic;
signal \pid_front.un1_pid_prereg_107_0_cascade_\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11\ : std_logic;
signal \uart_drone.N_145_cascade_\ : std_logic;
signal \uart_drone.un1_state_4_0_cascade_\ : std_logic;
signal \uart_drone.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_2\ : std_logic;
signal \uart_drone.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_drone.N_126_li\ : std_logic;
signal \uart_drone.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_4\ : std_logic;
signal \uart_drone.stateZ0Z_0\ : std_logic;
signal \uart_drone.stateZ0Z_1\ : std_logic;
signal \reset_module_System.reset6_15_cascade_\ : std_logic;
signal \reset_module_System.count_1_1_cascade_\ : std_logic;
signal \reset_module_System.reset6_3_cascade_\ : std_logic;
signal \reset_module_System.reset6_13\ : std_logic;
signal \reset_module_System.reset6_17_cascade_\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \reset_module_System.reset6_19_cascade_\ : std_logic;
signal \uart_drone.data_Auxce_0_0_0\ : std_logic;
signal \uart_drone.data_Auxce_0_0_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_3\ : std_logic;
signal \uart_drone.data_Auxce_0_5\ : std_logic;
signal \uart_drone.data_Auxce_0_6\ : std_logic;
signal \debug_CH0_16A_c\ : std_logic;
signal \uart_drone.un1_state_2_0\ : std_logic;
signal \uart_drone.state_RNIOU0NZ0Z_4\ : std_logic;
signal \uart_drone.data_AuxZ0Z_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_1\ : std_logic;
signal \uart_drone.data_AuxZ0Z_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_5\ : std_logic;
signal \uart_drone.data_AuxZ0Z_4\ : std_logic;
signal \uart_drone.data_AuxZ0Z_6\ : std_logic;
signal \uart_drone.data_AuxZ0Z_7\ : std_logic;
signal \uart_drone.data_rdyc_1_0\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2\ : std_logic;
signal \uart_drone.data_Auxce_0_0_4\ : std_logic;
signal \dron_frame_decoder_1.N_263_5\ : std_logic;
signal \dron_frame_decoder_1.N_263_5_cascade_\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\ : std_logic;
signal \dron_frame_decoder_1.N_219_4\ : std_logic;
signal \dron_frame_decoder_1.N_219_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_1_3\ : std_logic;
signal scaler_4_data_5 : std_logic;
signal \pid_front.O_0_5\ : std_logic;
signal \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_10\ : std_logic;
signal \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13_cascade_\ : std_logic;
signal \pid_front.pid_prereg_esr_RNICUKFAZ0Z_6_cascade_\ : std_logic;
signal \pid_front.un1_reset_0_i_cascade_\ : std_logic;
signal \pid_front.un1_reset_0_i_rn_0\ : std_logic;
signal \pid_front.m32_1_cascade_\ : std_logic;
signal \pid_front.un1_reset_0_i_sn\ : std_logic;
signal \pid_alt.error_i_acumm7lto5\ : std_logic;
signal \pid_alt.N_62_mux\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_5\ : std_logic;
signal \pid_alt.un1_reset_1_0_i\ : std_logic;
signal \pid_front.un1_pid_prereg_57\ : std_logic;
signal \pid_front.error_p_regZ0Z_18\ : std_logic;
signal \pid_front.un1_pid_prereg_18\ : std_logic;
signal \pid_front.error_p_regZ0Z_13\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_13\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13\ : std_logic;
signal \pid_front.pid_prereg_esr_RNI6FQ75Z0Z_23\ : std_logic;
signal \pid_front.un1_pid_prereg_42\ : std_logic;
signal \pid_front.un1_pid_prereg_47\ : std_logic;
signal \pid_front.un1_pid_prereg_42_cascade_\ : std_logic;
signal \pid_front.error_p_regZ0Z_16\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_16\ : std_logic;
signal \pid_front.un1_pid_prereg_35\ : std_logic;
signal \pid_front.un1_pid_prereg_36_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_30\ : std_logic;
signal \pid_front.error_p_regZ0Z_17\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_17\ : std_logic;
signal \pid_front.un1_pid_prereg_41\ : std_logic;
signal \pid_front.un1_pid_prereg_41_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_36\ : std_logic;
signal \pid_front.error_p_regZ0Z_11\ : std_logic;
signal \uart_drone.un1_state_7_0\ : std_logic;
signal \uart_drone.CO0\ : std_logic;
signal \uart_drone.stateZ0Z_3\ : std_logic;
signal \uart_drone.un1_state_4_0\ : std_logic;
signal \uart_drone.timer_CountZ1Z_3\ : std_logic;
signal \uart_drone.timer_CountZ0Z_4\ : std_logic;
signal \uart_drone.N_144_1\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \uart_drone.data_Auxce_0_1\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.reset6_11\ : std_logic;
signal \dron_frame_decoder_1.WDT10_0_i\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_0\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_1\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_2\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_3\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_4\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_5\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_7\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_8\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_9\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_10\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_11\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_12\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_14\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_14\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_15\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_9\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNIIVJ1Z0Z_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_13\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_10\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_11\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_8\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_12\ : std_logic;
signal \dron_frame_decoder_1.WDT10lto13_1\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.N_218\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3\ : std_logic;
signal throttle_order_5 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_13\ : std_logic;
signal throttle_order_13 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\ : std_logic;
signal throttle_order_10 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_13\ : std_logic;
signal \pid_alt.error_axbZ0Z_2\ : std_logic;
signal drone_altitude_2 : std_logic;
signal \pid_alt.error_axbZ0Z_3\ : std_logic;
signal drone_altitude_3 : std_logic;
signal \dron_frame_decoder_1.N_521_0\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_i_0\ : std_logic;
signal \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12_cascade_\ : std_logic;
signal \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10_cascade_\ : std_logic;
signal \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5_cascade_\ : std_logic;
signal \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5\ : std_logic;
signal \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10\ : std_logic;
signal \pid_front.error_p_regZ0Z_7\ : std_logic;
signal \pid_front.un1_pid_prereg_60_0_cascade_\ : std_logic;
signal \pid_front.N_1447_i_cascade_\ : std_logic;
signal \pid_front.error_p_regZ0Z_6\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_6\ : std_logic;
signal \pid_front.un1_pid_prereg_50_0_cascade_\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_7\ : std_logic;
signal \pid_front.m26_e_5_cascade_\ : std_logic;
signal \pid_front.m26_e_1_cascade_\ : std_logic;
signal \pid_front.m26_e_5\ : std_logic;
signal \pid_front.pid_prereg_esr_RNIGSMQ1Z0Z_10\ : std_logic;
signal \pid_front.m18_s_5\ : std_logic;
signal \pid_front.m18_s_4\ : std_logic;
signal \pid_front.m9_e_4_cascade_\ : std_logic;
signal \pid_front.m9_e_5\ : std_logic;
signal \pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20\ : std_logic;
signal \pid_front.pid_prereg_esr_RNIVDO51Z0Z_10\ : std_logic;
signal \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12\ : std_logic;
signal \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13\ : std_logic;
signal \pid_front.state_0_1\ : std_logic;
signal \pid_front.un1_reset_0_i\ : std_logic;
signal \pid_front.state_RNIVIRQZ0Z_0_cascade_\ : std_logic;
signal \pid_front.error_p_regZ0Z_10\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI653NZ0Z_10_cascade_\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_10\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI653NZ0Z_10\ : std_logic;
signal \pid_front.N_1463_i\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIM6G7Z0Z_9\ : std_logic;
signal \uart_drone.N_152\ : std_logic;
signal \pid_side.state_0_0\ : std_logic;
signal \uart_drone.bit_CountZ0Z_2\ : std_logic;
signal \uart_drone.bit_CountZ0Z_1\ : std_logic;
signal \uart_drone.bit_CountZ0Z_0\ : std_logic;
signal \uart_drone.data_Auxce_0_3\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \frame_decoder_CH4data_1\ : std_logic;
signal \frame_decoder_OFF4data_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH4data_2\ : std_logic;
signal \frame_decoder_OFF4data_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH4data_3\ : std_logic;
signal \frame_decoder_OFF4data_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH4data_4\ : std_logic;
signal \frame_decoder_OFF4data_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH4data_5\ : std_logic;
signal \frame_decoder_OFF4data_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_OFF4data_6\ : std_logic;
signal \frame_decoder_CH4data_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8\ : std_logic;
signal \frame_decoder_OFF4data_7\ : std_logic;
signal \frame_decoder_CH4data_7\ : std_logic;
signal \scaler_4.N_1849_i_l_ofxZ0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\ : std_logic;
signal throttle_order_6 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\ : std_logic;
signal throttle_order_3 : std_logic;
signal throttle_order_9 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_3_THRU_CO\ : std_logic;
signal throttle_order_4 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\ : std_logic;
signal throttle_order_8 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\ : std_logic;
signal throttle_order_12 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_1_THRU_CO\ : std_logic;
signal throttle_order_0 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\ : std_logic;
signal throttle_order_7 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\ : std_logic;
signal \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\ : std_logic;
signal \pid_front.error_p_regZ0Z_3\ : std_logic;
signal \pid_front.un1_pid_prereg_2_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_0\ : std_logic;
signal \pid_front.un1_pid_prereg_2\ : std_logic;
signal \pid_front.un1_pid_prereg_0_cascade_\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_3\ : std_logic;
signal \drone_H_disp_front_1\ : std_logic;
signal \dron_frame_decoder_1.N_489_0\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_0\ : std_logic;
signal \pid_front.pid_preregZ0Z_2\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_1\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIH7Q01Z0Z_1\ : std_logic;
signal \pid_front.pid_preregZ0Z_3\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_0_0\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIJCSGZ0Z_2\ : std_logic;
signal \pid_front.error_p_reg_esr_RNICVO11Z0Z_2\ : std_logic;
signal \pid_front.pid_preregZ0Z_4\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_1_0\ : std_logic;
signal \pid_front.pid_preregZ0Z_5\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_2\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIH8R01Z0Z_5\ : std_logic;
signal \pid_front.pid_preregZ0Z_6\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_3\ : std_logic;
signal \pid_front.error_d_reg_esr_RNIIFUFZ0Z_6\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI94TVZ0Z_6\ : std_logic;
signal \pid_front.pid_preregZ0Z_7\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_4\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_5\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIJETVZ0Z_7\ : std_logic;
signal \pid_front.error_d_reg_esr_RNINKUFZ0Z_7\ : std_logic;
signal \pid_front.pid_preregZ0Z_8\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \pid_front.error_d_reg_esr_RNISPUFZ0Z_8\ : std_logic;
signal \pid_front.error_p_reg_esr_RNITOTVZ0Z_8\ : std_logic;
signal \pid_front.pid_preregZ0Z_9\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_6\ : std_logic;
signal \pid_front.error_d_reg_esr_RNISPQT1Z0Z_10\ : std_logic;
signal \pid_front.error_d_reg_esr_RNI1VUFZ0Z_9\ : std_logic;
signal \pid_front.pid_preregZ0Z_10\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_7\ : std_logic;
signal \pid_front.error_d_reg_esr_RNI9NAB3Z0Z_10\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10\ : std_logic;
signal \pid_front.pid_preregZ0Z_11\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_8\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIESET1Z0Z_10\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI1E6A4Z0Z_12\ : std_logic;
signal \pid_front.pid_preregZ0Z_12\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_9\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12\ : std_logic;
signal \pid_front.error_d_reg_esr_RNIBO6A4Z0Z_12\ : std_logic;
signal \pid_front.pid_preregZ0Z_13\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_10\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIO6FT1Z0Z_12\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIN47A4Z0Z_12\ : std_logic;
signal \pid_front.pid_preregZ0Z_14\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_11\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI42GP4Z0Z_13\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13\ : std_logic;
signal \pid_front.pid_preregZ0Z_15\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_12\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_13\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI54OC2Z0Z_14\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIGEGP4Z0Z_14\ : std_logic;
signal \pid_front.pid_preregZ0Z_16\ : std_logic;
signal \bfn_12_23_0_\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIBAOC2Z0Z_15\ : std_logic;
signal \pid_front.error_p_reg_esr_RNISQGP4Z0Z_15\ : std_logic;
signal \pid_front.pid_preregZ0Z_17\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_14\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIHGOC2Z0Z_16\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI87HP4Z0Z_16\ : std_logic;
signal \pid_front.pid_preregZ0Z_18\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_15\ : std_logic;
signal \pid_front.error_p_reg_esr_RNINMOC2Z0Z_17\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIKJHP4Z0Z_17\ : std_logic;
signal \pid_front.pid_preregZ0Z_19\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_16\ : std_logic;
signal \pid_front.error_p_reg_esr_RNITSOC2Z0Z_18\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI57KP4Z0Z_18\ : std_logic;
signal \pid_front.pid_preregZ0Z_20\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_17\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI8ARC2Z0Z_19\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIOUOP4Z0Z_19\ : std_logic;
signal \pid_front.pid_preregZ0Z_21\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_18\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI09RP4Z0Z_20\ : std_logic;
signal \pid_front.pid_preregZ0Z_22\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_19\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_20\ : std_logic;
signal \pid_front.pid_preregZ0Z_23\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\ : std_logic;
signal \pid_front.un1_pid_prereg_axb_21\ : std_logic;
signal front_command_7 : std_logic;
signal \pid_front.error_p_regZ0Z_20\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_13\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8_c_RNIS918\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_9\ : std_logic;
signal scaler_4_data_14 : std_logic;
signal \scaler_4.debug_CH3_20A_c_0\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\ : std_logic;
signal scaler_4_data_7 : std_logic;
signal \ppm_encoder_1.N_134_0_cascade_\ : std_logic;
signal ppm_output_c : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\ : std_logic;
signal throttle_order_2 : std_logic;
signal scaler_4_data_6 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_4_THRU_CO\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_0\ : std_logic;
signal front_order_2 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_1_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_2\ : std_logic;
signal front_order_4 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_3_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_3\ : std_logic;
signal front_order_5 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_4_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_4\ : std_logic;
signal front_order_6 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_5_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7\ : std_logic;
signal front_order_8 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal front_order_9 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8\ : std_logic;
signal front_order_10 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9\ : std_logic;
signal front_order_11 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_13\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_13\ : std_logic;
signal \ppm_encoder_1.N_299\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_13\ : std_logic;
signal front_order_13 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_13\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_7\ : std_logic;
signal \pid_front.error_p_regZ0Z_2\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_2\ : std_logic;
signal \pid_front.error_d_reg_esr_RNIOBP11Z0Z_5\ : std_logic;
signal \pid_front.un1_pid_prereg_40_0\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4\ : std_logic;
signal \pid_front.error_p_regZ0Z_5\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_\ : std_logic;
signal \pid_front.error_d_reg_esr_RNIVOSGZ0Z_5\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_5\ : std_logic;
signal \pid_front.error_p_regZ0Z_4\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_4\ : std_logic;
signal \pid_front.un1_pid_prereg_17\ : std_logic;
signal \pid_front.un1_pid_prereg_17_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg_3\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIPISGZ0Z_3\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI4KF7Z0Z_0_cascade_\ : std_logic;
signal \pid_front.error_d_reg_esr_RNINGRVZ0Z_1\ : std_logic;
signal \pid_front.error_p_regZ0Z_1\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1_cascade_\ : std_logic;
signal \pid_front.un1_pid_prereg\ : std_logic;
signal \drone_H_disp_front_3\ : std_logic;
signal \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIUQTFZ0Z_1\ : std_logic;
signal \pid_alt.error_d_regZ0Z_15\ : std_logic;
signal \pid_alt.error_p_regZ0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_5\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_4\ : std_logic;
signal \pid_front.error_p_regZ0Z_0\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_0\ : std_logic;
signal \pid_front.N_1427_i\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_6\ : std_logic;
signal \drone_H_disp_front_2\ : std_logic;
signal \drone_H_disp_front_0\ : std_logic;
signal \pid_front.error_axb_0\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \pid_front.error_axbZ0Z_1\ : std_logic;
signal \pid_front.error_1\ : std_logic;
signal \pid_front.error_cry_0\ : std_logic;
signal \pid_front.error_axbZ0Z_2\ : std_logic;
signal \pid_front.error_2\ : std_logic;
signal \pid_front.error_cry_1\ : std_logic;
signal \pid_front.error_axbZ0Z_3\ : std_logic;
signal \pid_front.error_3\ : std_logic;
signal \pid_front.error_cry_2\ : std_logic;
signal \drone_H_disp_front_i_4\ : std_logic;
signal front_command_0 : std_logic;
signal \pid_front.error_4\ : std_logic;
signal \pid_front.error_cry_3\ : std_logic;
signal \drone_H_disp_front_i_5\ : std_logic;
signal front_command_1 : std_logic;
signal \pid_front.error_5\ : std_logic;
signal \pid_front.error_cry_0_0\ : std_logic;
signal \drone_H_disp_front_i_6\ : std_logic;
signal front_command_2 : std_logic;
signal \pid_front.error_6\ : std_logic;
signal \pid_front.error_cry_1_0\ : std_logic;
signal \drone_H_disp_front_i_7\ : std_logic;
signal front_command_3 : std_logic;
signal \pid_front.error_7\ : std_logic;
signal \pid_front.error_cry_2_0\ : std_logic;
signal \pid_front.error_cry_3_0\ : std_logic;
signal \drone_H_disp_front_i_8\ : std_logic;
signal front_command_4 : std_logic;
signal \pid_front.error_8\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal front_command_5 : std_logic;
signal \pid_front.error_9\ : std_logic;
signal \pid_front.error_cry_4\ : std_logic;
signal \drone_H_disp_front_i_10\ : std_logic;
signal front_command_6 : std_logic;
signal \pid_front.error_10\ : std_logic;
signal \pid_front.error_cry_5\ : std_logic;
signal \pid_front.error_axbZ0Z_7\ : std_logic;
signal \pid_front.error_11\ : std_logic;
signal \pid_front.error_cry_6\ : std_logic;
signal \pid_front.error_axb_8_l_ofx_0\ : std_logic;
signal \pid_front.error_12\ : std_logic;
signal \pid_front.error_cry_7\ : std_logic;
signal \drone_H_disp_front_i_12\ : std_logic;
signal \pid_front.error_13\ : std_logic;
signal \pid_front.error_cry_8\ : std_logic;
signal \drone_H_disp_front_i_13\ : std_logic;
signal \pid_front.error_14\ : std_logic;
signal \pid_front.error_cry_9\ : std_logic;
signal \pid_front.error_cry_10\ : std_logic;
signal \pid_front.error_15\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_10\ : std_logic;
signal \drone_H_disp_front_11\ : std_logic;
signal \drone_H_disp_front_12\ : std_logic;
signal \drone_H_disp_front_14\ : std_logic;
signal \drone_H_disp_front_15\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_8\ : std_logic;
signal \pid_alt.state_0_0\ : std_logic;
signal \pid_alt.state_1_0_0\ : std_logic;
signal scaler_4_data_9 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\ : std_logic;
signal scaler_4_data_8 : std_logic;
signal scaler_4_data_10 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\ : std_logic;
signal scaler_4_data_13 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\ : std_logic;
signal \pid_alt.N_72_i\ : std_logic;
signal \pid_alt.stateZ0Z_0\ : std_logic;
signal scaler_4_data_11 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\ : std_logic;
signal scaler_4_data_12 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_298_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_12\ : std_logic;
signal front_order_12 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_12\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_11\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_297_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_11\ : std_logic;
signal throttle_order_11 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_9\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_9\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_295\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_6\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_6\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_6\ : std_logic;
signal \ppm_encoder_1.N_292_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_5_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_7\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_7\ : std_logic;
signal \ppm_encoder_1.N_293_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\ : std_logic;
signal front_order_7 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_8\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_8\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_8\ : std_logic;
signal \ppm_encoder_1.N_294_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_14\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_14\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_14\ : std_logic;
signal \ppm_encoder_1.N_300_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_14\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_10_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_10\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_7\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_10\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_10\ : std_logic;
signal \ppm_encoder_1.N_296_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_10\ : std_logic;
signal \drone_H_disp_front_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_2150_i\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_7\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_15\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_17\ : std_logic;
signal \ppm_encoder_1.N_419_g\ : std_logic;
signal \debug_CH3_20A_c\ : std_logic;
signal uart_drone_data_rdy : std_logic;
signal \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_313_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_12\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_12\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\ : std_logic;
signal \scaler_4.un2_source_data_0\ : std_logic;
signal \frame_decoder_OFF4data_0\ : std_logic;
signal \frame_decoder_CH4data_0\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1_c_RNOZ0\ : std_logic;
signal side_order_2 : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\ : std_logic;
signal \ppm_encoder_1.N_221_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_5\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.throttle_m_1\ : std_logic;
signal \ppm_encoder_1.N_287_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\ : std_logic;
signal side_order_1 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_0_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_0_THRU_CO\ : std_logic;
signal front_order_1 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\ : std_logic;
signal throttle_order_1 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_1\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIUINC6Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_2\ : std_logic;
signal \ppm_encoder_1.elevator_RNIFISN6Z0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_3\ : std_logic;
signal \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_4\ : std_logic;
signal \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_5\ : std_logic;
signal \ppm_encoder_1.throttle_RNILVOO6Z0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_7\ : std_logic;
signal \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_8\ : std_logic;
signal \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_9\ : std_logic;
signal \ppm_encoder_1.elevator_RNIC22D6Z0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_10\ : std_logic;
signal \ppm_encoder_1.elevator_RNIH72D6Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_11\ : std_logic;
signal \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_12\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_15\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_18\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_0\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_4\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_12\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_4\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_7\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_2\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\ : std_logic;
signal \ppm_encoder_1.N_232_cascade_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_14\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_13\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_6\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_5\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_4\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_12\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_8\ : std_logic;
signal \ppm_encoder_1.N_139_17\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\ : std_logic;
signal \ppm_encoder_1.N_139_17_cascade_\ : std_logic;
signal \ppm_encoder_1.N_139\ : std_logic;
signal \pid_front.un1_pid_prereg_92\ : std_logic;
signal \pid_front.un1_pid_prereg_93\ : std_logic;
signal \pid_front.error_p_reg_esr_RNIGKTC2Z0Z_20\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_16\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_16\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_17\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_15\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_16\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_20\ : std_logic;
signal side_order_10 : std_logic;
signal side_order_11 : std_logic;
signal side_order_6 : std_logic;
signal side_order_7 : std_logic;
signal side_order_8 : std_logic;
signal side_order_9 : std_logic;
signal side_order_0 : std_logic;
signal side_order_5 : std_logic;
signal side_order_4 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_5\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_5\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_6\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_2_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.N_221\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_0_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_232\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_0\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_3\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_3_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIT3R05Z0Z_3\ : std_logic;
signal \ppm_encoder_1.N_289\ : std_logic;
signal side_order_3 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_2_THRU_CO\ : std_logic;
signal front_order_3 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_18\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_14\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_16\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_16\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_11_mux\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_3\ : std_logic;
signal \ppm_encoder_1.N_2150_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_10\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_9\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_11\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_17\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_17\ : std_logic;
signal \pid_side.m32_1\ : std_logic;
signal reset_system : std_logic;
signal \pid_side.m26_e_5_cascade_\ : std_logic;
signal \pid_side.N_11_0_cascade_\ : std_logic;
signal \pid_side.pid_prereg_esr_RNILRSP2Z0Z_5\ : std_logic;
signal \pid_side.m26_e_5\ : std_logic;
signal \pid_side.pid_prereg_esr_RNIGJDR1Z0Z_10_cascade_\ : std_logic;
signal \pid_side.m18_s_4\ : std_logic;
signal \pid_side.pid_prereg_esr_RNIQBAH2Z0Z_23_cascade_\ : std_logic;
signal \pid_side.un1_reset_0_i_sn\ : std_logic;
signal \pid_side.i19_mux_cascade_\ : std_logic;
signal \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12\ : std_logic;
signal \pid_side.N_11_0\ : std_logic;
signal \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12_cascade_\ : std_logic;
signal \pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10\ : std_logic;
signal \pid_side.N_82_mux\ : std_logic;
signal side_order_12 : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_2_sqmuxa_0\ : std_logic;
signal front_order_0 : std_logic;
signal pid_altitude_dv : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_6\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_0_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_5\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_7\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_8\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_8\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_9\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_9\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\ : std_logic;
signal scaler_4_data_4 : std_logic;
signal \ppm_encoder_1.rudderZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pid_altitude_dv_0\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_314_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_10\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_7\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_11\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_12\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_12\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_2\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_2\ : std_logic;
signal \ppm_encoder_1.N_288\ : std_logic;
signal \ppm_encoder_1.N_290\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_153_d\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_15\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_11\ : std_logic;
signal \pid_alt.state_RNIFCSD1Z0Z_0\ : std_logic;
signal \pid_alt.N_664_0\ : std_logic;
signal \pid_side.pid_preregZ0Z_0\ : std_logic;
signal \pid_side.pid_preregZ0Z_1\ : std_logic;
signal \debug_CH1_0A_c\ : std_logic;
signal \pid_side.stateZ0Z_0\ : std_logic;
signal \pid_side.m18_s_5\ : std_logic;
signal \pid_side.stateZ0Z_1\ : std_logic;
signal \pid_side.un1_reset_0_i_rn_0\ : std_logic;
signal \pid_side.m26_e_1\ : std_logic;
signal \pid_side.m9_e_4\ : std_logic;
signal \pid_side.m9_e_5_cascade_\ : std_logic;
signal \pid_side.pid_prereg_esr_RNIFB07Z0Z_20\ : std_logic;
signal \pid_side.pid_prereg_esr_RNIFB07Z0Z_20_cascade_\ : std_logic;
signal side_order_13 : std_logic;
signal \pid_side.state_0_1\ : std_logic;
signal \pid_side.un1_reset_0_i\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_13\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_11\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_8\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_11\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_16\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_16\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_18\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_53_d\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_18\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_5\ : std_logic;
signal \pid_front.un1_pid_prereg_axb_0\ : std_logic;
signal \pid_front.pid_preregZ0Z_0\ : std_logic;
signal \pid_front.error_d_reg_prevZ0Z_18\ : std_logic;
signal \pid_front.state_0_g_0\ : std_logic;
signal \pid_front.O_6\ : std_logic;
signal \pid_front.error_d_regZ0Z_2\ : std_logic;
signal \GB_BUFFER_reset_system_g_THRU_CO\ : std_logic;
signal \bfn_20_9_0_\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_0_THRU_CO\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_0\ : std_logic;
signal \pid_side.pid_preregZ0Z_2\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_1\ : std_logic;
signal \pid_side.pid_preregZ0Z_3\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_0_0\ : std_logic;
signal \pid_side.pid_preregZ0Z_4\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_1_0\ : std_logic;
signal \pid_side.pid_preregZ0Z_5\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_2\ : std_logic;
signal \pid_side.pid_preregZ0Z_6\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_3\ : std_logic;
signal \pid_side.pid_preregZ0Z_7\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_4\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_5\ : std_logic;
signal \pid_side.pid_preregZ0Z_8\ : std_logic;
signal \bfn_20_10_0_\ : std_logic;
signal \pid_side.pid_preregZ0Z_9\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_6\ : std_logic;
signal \pid_side.pid_preregZ0Z_10\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_7\ : std_logic;
signal \pid_side.pid_preregZ0Z_11\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_8\ : std_logic;
signal \pid_side.pid_preregZ0Z_12\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_9\ : std_logic;
signal \pid_side.pid_preregZ0Z_13\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_10\ : std_logic;
signal \pid_side.pid_preregZ0Z_14\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_11\ : std_logic;
signal \pid_side.pid_preregZ0Z_15\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_12\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_13\ : std_logic;
signal \pid_side.pid_preregZ0Z_16\ : std_logic;
signal \bfn_20_11_0_\ : std_logic;
signal \pid_side.pid_preregZ0Z_17\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_14\ : std_logic;
signal \pid_side.pid_preregZ0Z_18\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_15\ : std_logic;
signal \pid_side.pid_preregZ0Z_19\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_16\ : std_logic;
signal \pid_side.pid_preregZ0Z_20\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_17\ : std_logic;
signal \pid_side.pid_preregZ0Z_21\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_18\ : std_logic;
signal \pid_side.pid_preregZ0Z_22\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_19\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_20\ : std_logic;
signal \pid_side.pid_preregZ0Z_23\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNILHF23Z0Z_18\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIJV5H1Z0Z_15\ : std_logic;
signal \pid_side.un1_pid_prereg_30_cascade_\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI0PB23Z0Z_14\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI4UC23Z0Z_17\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI5I6H1Z0Z_18\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIP56H1Z0Z_16\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_16\ : std_logic;
signal \pid_side.un1_pid_prereg_35\ : std_logic;
signal \pid_side.un1_pid_prereg_36_cascade_\ : std_logic;
signal \pid_side.un1_pid_prereg_30\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIC5C23Z0Z_15\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI89K23Z0Z_19\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIGJM23Z0Z_20\ : std_logic;
signal \pid_side.un1_pid_prereg_axb_21\ : std_logic;
signal \ppm_encoder_1.N_286\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIGV8H1Z0Z_19\ : std_logic;
signal \drone_H_disp_side_1\ : std_logic;
signal uart_drone_data_2 : std_logic;
signal \drone_H_disp_side_2\ : std_logic;
signal \drone_H_disp_side_3\ : std_logic;
signal \dron_frame_decoder_1.N_505_0\ : std_logic;
signal \drone_H_disp_front_i_9\ : std_logic;
signal uart_drone_data_1 : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_9\ : std_logic;
signal \dron_frame_decoder_1.N_481_0\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_4\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_6\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_7\ : std_logic;
signal \pid_front.stateZ0Z_1\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_0_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_axb_1\ : std_logic;
signal \pid_front.stateZ0Z_0\ : std_logic;
signal \pid_front.pid_preregZ0Z_1\ : std_logic;
signal side_command_7 : std_logic;
signal \pid_front.O_7\ : std_logic;
signal \pid_front.error_d_regZ0Z_3\ : std_logic;
signal \pid_side.error_p_reg_esr_RNI5QI23Z0Z_5\ : std_logic;
signal \pid_side.un1_pid_prereg_axb_1\ : std_logic;
signal \pid_side.error_p_reg_esr_RNISH6JZ0Z_0_cascade_\ : std_logic;
signal \pid_side.error_d_reg_esr_RNIFP9R2Z0Z_1\ : std_logic;
signal \pid_side.N_1546_i\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_1\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1_cascade_\ : std_logic;
signal \pid_side.un1_pid_prereg\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_0\ : std_logic;
signal \pid_side.un1_pid_prereg_axb_0\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIAVKD1Z0Z_1\ : std_logic;
signal \pid_side.un1_pid_prereg_18_cascade_\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13_cascade_\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_13\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI4NA21Z0Z_12\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIDP5H1Z0Z_14\ : std_logic;
signal \pid_side.error_d_reg_esr_RNIKMFP2Z0Z_10\ : std_logic;
signal \pid_side.N_1582_i\ : std_logic;
signal \pid_side.N_1582_i_cascade_\ : std_logic;
signal \pid_side.error_d_reg_esr_RNI104E2Z0Z_10\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIKCB23Z0Z_13\ : std_logic;
signal \pid_side.un1_pid_prereg_23\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13\ : std_logic;
signal \pid_side.un1_pid_prereg_18\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIBAGJ2Z0Z_12\ : std_logic;
signal \pid_side.un1_pid_prereg_29\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIO9BH1Z0Z_20\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNILJFJ2Z0Z_12\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10_cascade_\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11_cascade_\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIQCA21Z0Z_10\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12\ : std_logic;
signal \pid_side.N_1590_i_cascade_\ : std_logic;
signal \pid_side.error_d_reg_esr_RNIVTFJ2Z0Z_12\ : std_logic;
signal \pid_side.un1_pid_prereg_107_0\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_12\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNI2VN9Z0Z_12\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_11\ : std_logic;
signal \pid_side.O_2_15\ : std_logic;
signal \pid_side.error_p_regZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_291\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\ : std_logic;
signal \pid_side.un1_pid_prereg_56\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_19\ : std_logic;
signal \pid_side.un1_pid_prereg_57\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\ : std_logic;
signal \drone_H_disp_side_0\ : std_logic;
signal \pid_side.error_axb_0\ : std_logic;
signal \bfn_21_17_0_\ : std_logic;
signal \pid_side.error_axbZ0Z_1\ : std_logic;
signal \pid_side.error_1\ : std_logic;
signal \pid_side.error_cry_0\ : std_logic;
signal \pid_side.error_axbZ0Z_2\ : std_logic;
signal \pid_side.error_2\ : std_logic;
signal \pid_side.error_cry_1\ : std_logic;
signal \pid_side.error_axbZ0Z_3\ : std_logic;
signal \pid_side.error_3\ : std_logic;
signal \pid_side.error_cry_2\ : std_logic;
signal \drone_H_disp_side_i_4\ : std_logic;
signal side_command_0 : std_logic;
signal \pid_side.error_4\ : std_logic;
signal \pid_side.error_cry_3\ : std_logic;
signal \drone_H_disp_side_i_5\ : std_logic;
signal side_command_1 : std_logic;
signal \pid_side.error_5\ : std_logic;
signal \pid_side.error_cry_0_0\ : std_logic;
signal \drone_H_disp_side_i_6\ : std_logic;
signal side_command_2 : std_logic;
signal \pid_side.error_6\ : std_logic;
signal \pid_side.error_cry_1_0\ : std_logic;
signal \drone_H_disp_side_i_7\ : std_logic;
signal side_command_3 : std_logic;
signal \pid_side.error_7\ : std_logic;
signal \pid_side.error_cry_2_0\ : std_logic;
signal \pid_side.error_cry_3_0\ : std_logic;
signal \drone_H_disp_side_i_8\ : std_logic;
signal side_command_4 : std_logic;
signal \pid_side.error_8\ : std_logic;
signal \bfn_21_18_0_\ : std_logic;
signal \drone_H_disp_side_i_9\ : std_logic;
signal side_command_5 : std_logic;
signal \pid_side.error_9\ : std_logic;
signal \pid_side.error_cry_4\ : std_logic;
signal \drone_H_disp_side_i_10\ : std_logic;
signal side_command_6 : std_logic;
signal \pid_side.error_10\ : std_logic;
signal \pid_side.error_cry_5\ : std_logic;
signal \pid_side.error_axbZ0Z_7\ : std_logic;
signal \pid_side.error_11\ : std_logic;
signal \pid_side.error_cry_6\ : std_logic;
signal \pid_side.error_axb_8_l_ofxZ0\ : std_logic;
signal \pid_side.error_12\ : std_logic;
signal \pid_side.error_cry_7\ : std_logic;
signal \drone_H_disp_side_i_12\ : std_logic;
signal \pid_side.error_13\ : std_logic;
signal \pid_side.error_cry_8\ : std_logic;
signal \drone_H_disp_side_i_13\ : std_logic;
signal \pid_side.error_14\ : std_logic;
signal \pid_side.error_cry_9\ : std_logic;
signal \pid_side.error_cry_10\ : std_logic;
signal \pid_side.error_15\ : std_logic;
signal uart_drone_data_3 : std_logic;
signal \drone_H_disp_side_11\ : std_logic;
signal uart_drone_data_4 : std_logic;
signal \drone_H_disp_side_12\ : std_logic;
signal uart_drone_data_5 : std_logic;
signal \drone_H_disp_side_13\ : std_logic;
signal uart_drone_data_7 : std_logic;
signal \drone_H_disp_side_15\ : std_logic;
signal uart_drone_data_0 : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_8\ : std_logic;
signal \pid_front.O_10\ : std_logic;
signal \pid_front.error_d_regZ0Z_6\ : std_logic;
signal \pid_side.error_d_reg_esr_RNI76TK1Z0Z_5\ : std_logic;
signal \pid_side.un1_pid_prereg_40_0_cascade_\ : std_logic;
signal \pid_side.error_d_reg_esr_RNI86Q93Z0Z_5\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4\ : std_logic;
signal \pid_side.un1_pid_prereg_17_cascade_\ : std_logic;
signal \pid_side.error_p_reg_esr_RNI10TK1Z0Z_3\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_4\ : std_logic;
signal \pid_side.un1_pid_prereg_17\ : std_logic;
signal \pid_side.error_p_reg_esr_RNISPP93Z0Z_2\ : std_logic;
signal \pid_side.O_2_9\ : std_logic;
signal \pid_side.O_2_4\ : std_logic;
signal \pid_side.error_p_regZ0Z_0\ : std_logic;
signal \pid_side.state_RNINK4UZ0Z_0\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIE47JZ0Z_9\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_15\ : std_logic;
signal \pid_side.un1_pid_prereg_24\ : std_logic;
signal \pid_side.un1_pid_prereg_48\ : std_logic;
signal \pid_side.un1_pid_prereg_36\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIOHC23Z0Z_16\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_18\ : std_logic;
signal \pid_side.un1_pid_prereg_47\ : std_logic;
signal \pid_side.un1_pid_prereg_47_cascade_\ : std_logic;
signal \pid_side.error_d_reg_prev_esr_RNIVB6H1Z0Z_17\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_10\ : std_logic;
signal \pid_side.O_1_4\ : std_logic;
signal \pid_side.error_d_regZ0Z_0\ : std_logic;
signal \pid_side.O_1_8\ : std_logic;
signal \pid_side.error_d_regZ0Z_4\ : std_logic;
signal \pid_side.O_1_5\ : std_logic;
signal \pid_side.error_d_regZ0Z_1\ : std_logic;
signal uart_pc_data_4 : std_logic;
signal xy_kd_4 : std_logic;
signal uart_drone_data_6 : std_logic;
signal \drone_H_disp_side_14\ : std_logic;
signal \dron_frame_decoder_1.N_497_0\ : std_logic;
signal \pid_front.O_9\ : std_logic;
signal \pid_front.error_d_regZ0Z_5\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1\ : std_logic;
signal \pid_side.error_p_reg_esr_RNI5PH23Z0Z_1\ : std_logic;
signal \pid_side.un1_pid_prereg_2\ : std_logic;
signal \pid_side.un1_pid_prereg_2_cascade_\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIRPSK1Z0Z_2\ : std_logic;
signal \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2\ : std_logic;
signal \pid_side.un1_pid_prereg_0\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_3\ : std_logic;
signal \pid_side.un1_pid_prereg_3\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_2\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_14\ : std_logic;
signal \pid_side.error_p_regZ0Z_5\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_5\ : std_logic;
signal \pid_side.N_1566_i_cascade_\ : std_logic;
signal \pid_side.N_1578_i_cascade_\ : std_logic;
signal \pid_side.error_d_reg_esr_RNID3MD1Z0Z_9\ : std_logic;
signal \pid_side.N_1574_i_cascade_\ : std_logic;
signal \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8\ : std_logic;
signal \pid_side.un1_pid_prereg_80_0\ : std_logic;
signal \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8_cascade_\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIL1CR2Z0Z_8\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_8\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_9\ : std_logic;
signal \pid_side.un1_pid_prereg_41\ : std_logic;
signal \pid_side.un1_pid_prereg_42\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_17\ : std_logic;
signal \pid_side.O_1_13\ : std_logic;
signal \pid_side.error_d_regZ0Z_9\ : std_logic;
signal \pid_side.un1_pid_prereg_93\ : std_logic;
signal \pid_side.un1_pid_prereg_92\ : std_logic;
signal \pid_front.O_12\ : std_logic;
signal \pid_front.error_d_regZ0Z_8\ : std_logic;
signal \pid_front.O_16\ : std_logic;
signal \pid_front.error_d_regZ0Z_12\ : std_logic;
signal \pid_front.O_14\ : std_logic;
signal \pid_front.error_d_regZ0Z_10\ : std_logic;
signal \pid_side.O_2_8\ : std_logic;
signal \pid_side.error_p_regZ0Z_4\ : std_logic;
signal \pid_side.O_2_5\ : std_logic;
signal \pid_side.error_p_regZ0Z_1\ : std_logic;
signal \pid_side.O_2_7\ : std_logic;
signal \pid_side.error_p_regZ0Z_3\ : std_logic;
signal \pid_side.O_2_22\ : std_logic;
signal \pid_side.error_p_regZ0Z_18\ : std_logic;
signal \pid_side.O_2_6\ : std_logic;
signal \pid_side.error_p_regZ0Z_2\ : std_logic;
signal \pid_side.O_2_20\ : std_logic;
signal \pid_side.error_p_regZ0Z_16\ : std_logic;
signal \pid_side.O_2_21\ : std_logic;
signal \pid_side.error_p_regZ0Z_17\ : std_logic;
signal \pid_side.O_1_6\ : std_logic;
signal \pid_side.error_d_regZ0Z_2\ : std_logic;
signal \pid_side.O_2_17\ : std_logic;
signal \pid_side.error_p_regZ0Z_13\ : std_logic;
signal \pid_side.O_2_12\ : std_logic;
signal \pid_side.error_p_regZ0Z_8\ : std_logic;
signal \pid_side.O_2_24\ : std_logic;
signal \pid_side.error_p_regZ0Z_20\ : std_logic;
signal \pid_side.O_2_18\ : std_logic;
signal \pid_side.error_p_regZ0Z_14\ : std_logic;
signal \pid_side.O_2_14\ : std_logic;
signal \pid_side.error_p_regZ0Z_10\ : std_logic;
signal \pid_side.O_2_19\ : std_logic;
signal \pid_side.error_p_regZ0Z_15\ : std_logic;
signal \pid_side.O_2_10\ : std_logic;
signal \pid_side.O_2_13\ : std_logic;
signal \pid_side.error_p_regZ0Z_9\ : std_logic;
signal \pid_side.O_2_11\ : std_logic;
signal \pid_side.O_2_23\ : std_logic;
signal \pid_side.error_p_regZ0Z_19\ : std_logic;
signal \pid_side.O_2_16\ : std_logic;
signal \pid_side.error_p_regZ0Z_12\ : std_logic;
signal \pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6\ : std_logic;
signal \pid_side.un1_pid_prereg_60_0_cascade_\ : std_logic;
signal \pid_side.error_p_reg_esr_RNI1DBR2Z0Z_6\ : std_logic;
signal \pid_side.N_1570_i_cascade_\ : std_logic;
signal \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7\ : std_logic;
signal \pid_side.un1_pid_prereg_70_0\ : std_logic;
signal \pid_side.error_p_regZ0Z_7\ : std_logic;
signal \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7_cascade_\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_7\ : std_logic;
signal \pid_side.error_p_reg_esr_RNIBNBR2Z0Z_7\ : std_logic;
signal \pid_side.error_p_regZ0Z_6\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_6\ : std_logic;
signal \pid_side.un1_pid_prereg_50_0\ : std_logic;
signal \pid_side.O_1_15\ : std_logic;
signal \pid_side.error_d_regZ0Z_11\ : std_logic;
signal \pid_side.O_1_21\ : std_logic;
signal \pid_side.error_d_regZ0Z_17\ : std_logic;
signal \pid_side.O_1_19\ : std_logic;
signal \pid_side.error_d_regZ0Z_15\ : std_logic;
signal \pid_side.O_1_12\ : std_logic;
signal \pid_side.error_d_regZ0Z_8\ : std_logic;
signal \pid_side.O_1_9\ : std_logic;
signal \pid_side.error_d_regZ0Z_5\ : std_logic;
signal \pid_side.O_1_16\ : std_logic;
signal \pid_side.error_d_regZ0Z_12\ : std_logic;
signal \pid_side.O_1_18\ : std_logic;
signal \pid_side.error_d_regZ0Z_14\ : std_logic;
signal \pid_side.O_1_7\ : std_logic;
signal \pid_side.error_d_regZ0Z_3\ : std_logic;
signal \pid_side.O_1_17\ : std_logic;
signal \pid_side.error_d_regZ0Z_13\ : std_logic;
signal \pid_side.O_1_14\ : std_logic;
signal \pid_side.error_d_regZ0Z_10\ : std_logic;
signal \pid_side.O_1_23\ : std_logic;
signal \pid_side.error_d_regZ0Z_19\ : std_logic;
signal \pid_side.O_1_24\ : std_logic;
signal \pid_side.O_1_10\ : std_logic;
signal \pid_side.error_d_regZ0Z_6\ : std_logic;
signal \pid_side.O_1_22\ : std_logic;
signal \pid_side.error_d_regZ0Z_18\ : std_logic;
signal \pid_side.O_1_11\ : std_logic;
signal \pid_side.error_d_regZ0Z_7\ : std_logic;
signal \pid_side.O_1_20\ : std_logic;
signal \pid_side.error_d_regZ0Z_16\ : std_logic;
signal \pid_side.N_599_0\ : std_logic;
signal uart_pc_data_0 : std_logic;
signal xy_kd_0 : std_logic;
signal uart_pc_data_1 : std_logic;
signal xy_kd_1 : std_logic;
signal uart_pc_data_2 : std_logic;
signal xy_kd_2 : std_logic;
signal uart_pc_data_5 : std_logic;
signal xy_kd_5 : std_logic;
signal uart_pc_data_6 : std_logic;
signal xy_kd_6 : std_logic;
signal uart_pc_data_7 : std_logic;
signal xy_kd_7 : std_logic;
signal uart_pc_data_3 : std_logic;
signal xy_kd_3 : std_logic;
signal \Commands_frame_decoder.state_RNITUI31Z0Z_13\ : std_logic;
signal \pid_side.error_d_regZ0Z_20\ : std_logic;
signal \pid_side.error_d_reg_prevZ0Z_20\ : std_logic;
signal \pid_side.state_0_g_0\ : std_logic;
signal reset_system_g : std_logic;
signal \pid_front.O_4\ : std_logic;
signal \pid_front.error_d_regZ0Z_0\ : std_logic;
signal \pid_front.O_5\ : std_logic;
signal \pid_front.error_d_regZ0Z_1\ : std_logic;
signal \pid_front.O_17\ : std_logic;
signal \pid_front.error_d_regZ0Z_13\ : std_logic;
signal \pid_front.O_15\ : std_logic;
signal \pid_front.error_d_regZ0Z_11\ : std_logic;
signal \pid_front.O_13\ : std_logic;
signal \pid_front.error_d_regZ0Z_9\ : std_logic;
signal \pid_front.O_20\ : std_logic;
signal \pid_front.error_d_regZ0Z_16\ : std_logic;
signal \pid_front.O_21\ : std_logic;
signal \pid_front.error_d_regZ0Z_17\ : std_logic;
signal \pid_front.O_22\ : std_logic;
signal \pid_front.error_d_regZ0Z_18\ : std_logic;
signal \pid_front.O_23\ : std_logic;
signal \pid_front.error_d_regZ0Z_19\ : std_logic;
signal \pid_front.O_24\ : std_logic;
signal \pid_front.error_d_regZ0Z_20\ : std_logic;
signal \pid_front.O_18\ : std_logic;
signal \pid_front.error_d_regZ0Z_14\ : std_logic;
signal \pid_front.O_8\ : std_logic;
signal \pid_front.error_d_regZ0Z_4\ : std_logic;
signal \pid_front.O_11\ : std_logic;
signal \pid_front.error_d_regZ0Z_7\ : std_logic;
signal \pid_front.O_19\ : std_logic;
signal \pid_front.error_d_regZ0Z_15\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_system_pll_g : std_logic;
signal \pid_front.N_543_0\ : std_logic;
signal \N_665_g\ : std_logic;

signal clk_system_wire : std_logic;
signal uart_input_pc_wire : std_logic;
signal \debug_CH2_18A_wire\ : std_logic;
signal \debug_CH0_16A_wire\ : std_logic;
signal \debug_CH1_0A_wire\ : std_logic;
signal \debug_CH5_31B_wire\ : std_logic;
signal \debug_CH4_2A_wire\ : std_logic;
signal ppm_output_wire : std_logic;
signal \debug_CH3_20A_wire\ : std_logic;
signal \debug_CH6_5B_wire\ : std_logic;
signal uart_input_drone_wire : std_logic;
signal \Pc2drone_pll_inst.Pc2drone_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_side.un2_error_1_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_1_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_1_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_1_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_1_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_front.un2_error_1_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_1_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_1_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_1_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_1_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    clk_system_wire <= clk_system;
    uart_input_pc_wire <= uart_input_pc;
    debug_CH2_18A <= \debug_CH2_18A_wire\;
    debug_CH0_16A <= \debug_CH0_16A_wire\;
    debug_CH1_0A <= \debug_CH1_0A_wire\;
    debug_CH5_31B <= \debug_CH5_31B_wire\;
    debug_CH4_2A <= \debug_CH4_2A_wire\;
    ppm_output <= ppm_output_wire;
    debug_CH3_20A <= \debug_CH3_20A_wire\;
    debug_CH6_5B <= \debug_CH6_5B_wire\;
    uart_input_drone_wire <= uart_input_drone;
    \Pc2drone_pll_inst.Pc2drone_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pid_alt.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_A_wire\ <= \N__24010\&\N__24062\&\N__24100\&\N__24152\&\N__24205\&\N__23542\&\N__23605\&\N__23668\&\N__23731\&\N__23794\&\N__23848\&\N__23908\&\N__23338\&\N__23386\&\N__23422\&\N__30685\;
    \pid_alt.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24312\&\N__23946\&\N__25680\&\N__29316\&\N__24303\&\N__25692\&\N__23976\&\N__23958\;
    \pid_alt.O_5_24\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_5_23\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_5_22\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_5_21\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_5_20\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_5_19\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_5_18\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_5_17\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_5_16\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_5_15\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_5_14\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_5_13\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_5_12\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_5_11\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_5_10\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_5_9\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_5_8\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_5_7\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_5_6\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_5_5\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_5_4\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ <= \N__24017\&\N__24058\&\N__24107\&\N__24151\&\N__24206\&\N__23543\&\N__23606\&\N__23669\&\N__23732\&\N__23795\&\N__23849\&\N__23909\&\N__23345\&\N__23387\&\N__23429\&\N__30686\;
    \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22083\&\N__22095\&\N__22041\&\N__22050\&\N__22059\&\N__22632\&\N__22071\&\N__22644\;
    \pid_alt.O_4_24\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_4_23\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_4_22\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_4_21\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_4_20\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_4_19\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_4_18\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_4_17\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_4_16\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_4_15\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_4_14\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_4_13\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_4_12\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_4_11\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_4_10\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_4_9\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_4_8\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_4_7\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_4_6\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_4_5\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_4_4\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\ <= \N__24021\&\N__24063\&\N__24111\&\N__24159\&\N__24207\&\N__23550\&\N__23610\&\N__23676\&\N__23733\&\N__23796\&\N__23856\&\N__23916\&\N__23352\&\N__23394\&\N__23436\&\N__30693\;
    \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21969\&\N__22686\&\N__22101\&\N__22677\&\N__22668\&\N__21963\&\N__21957\&\N__22656\;
    \pid_alt.O_3_24\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_3_23\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_3_22\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_3_21\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_3_20\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_3_19\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_3_18\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_3_17\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_3_16\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_3_15\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_3_14\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_3_13\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_3_12\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_3_11\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_3_10\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_3_9\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_3_8\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_3_7\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_3_6\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_3_5\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_3_4\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(4);
    \pid_front.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_front.un2_error_mulonly_0_24_0_A_wire\ <= \N__39453\&\N__39498\&\N__38960\&\N__39003\&\N__39051\&\N__39099\&\N__39159\&\N__39210\&\N__39270\&\N__39326\&\N__38634\&\N__38691\&\N__38751\&\N__38802\&\N__38853\&\N__38912\;
    \pid_front.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_front.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__31967\&\N__30758\&\N__30722\&\N__29423\&\N__32006\&\N__32033\&\N__32076\&\N__32111\;
    \pid_front.O_0_24\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(24);
    \pid_front.O_0_23\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(23);
    \pid_front.O_0_22\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(22);
    \pid_front.O_0_21\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(21);
    \pid_front.O_0_20\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(20);
    \pid_front.O_0_19\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(19);
    \pid_front.O_0_18\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_front.O_0_17\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_front.O_0_16\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_front.O_0_15\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_front.O_0_14\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_front.O_0_13\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_front.O_0_12\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_front.O_0_11\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_front.O_0_10\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_front.O_0_9\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_front.O_0_8\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_front.O_0_7\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_front.O_0_6\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_front.O_0_5\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_front.O_0_4\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(4);
    \pid_side.un2_error_1_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_side.un2_error_1_mulonly_0_24_0_A_wire\ <= \N__52736\&\N__52769\&\N__51869\&\N__51905\&\N__51941\&\N__51977\&\N__52028\&\N__52082\&\N__52127\&\N__52166\&\N__51575\&\N__51620\&\N__51665\&\N__51704\&\N__51740\&\N__51779\;
    \pid_side.un2_error_1_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_side.un2_error_1_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__55388\&\N__55595\&\N__55766\&\N__53249\&\N__55223\&\N__55943\&\N__56153\&\N__56324\;
    \pid_side.O_1_24\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(24);
    \pid_side.O_1_23\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(23);
    \pid_side.O_1_22\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(22);
    \pid_side.O_1_21\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(21);
    \pid_side.O_1_20\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(20);
    \pid_side.O_1_19\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(19);
    \pid_side.O_1_18\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(18);
    \pid_side.O_1_17\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(17);
    \pid_side.O_1_16\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(16);
    \pid_side.O_1_15\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(15);
    \pid_side.O_1_14\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(14);
    \pid_side.O_1_13\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(13);
    \pid_side.O_1_12\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(12);
    \pid_side.O_1_11\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(11);
    \pid_side.O_1_10\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(10);
    \pid_side.O_1_9\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(9);
    \pid_side.O_1_8\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(8);
    \pid_side.O_1_7\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(7);
    \pid_side.O_1_6\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(6);
    \pid_side.O_1_5\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(5);
    \pid_side.O_1_4\ <= \pid_side.un2_error_1_mulonly_0_24_0_O_wire\(4);
    \pid_side.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_side.un2_error_mulonly_0_24_0_A_wire\ <= \N__52740\&\N__52770\&\N__51873\&\N__51909\&\N__51945\&\N__51981\&\N__52032\&\N__52086\&\N__52131\&\N__52173\&\N__51582\&\N__51627\&\N__51672\&\N__51708\&\N__51744\&\N__51786\;
    \pid_side.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_side.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__31971\&\N__30762\&\N__30729\&\N__29433\&\N__32010\&\N__32043\&\N__32075\&\N__32115\;
    \pid_side.O_2_24\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(24);
    \pid_side.O_2_23\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(23);
    \pid_side.O_2_22\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(22);
    \pid_side.O_2_21\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(21);
    \pid_side.O_2_20\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(20);
    \pid_side.O_2_19\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(19);
    \pid_side.O_2_18\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_side.O_2_17\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_side.O_2_16\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_side.O_2_15\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_side.O_2_14\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_side.O_2_13\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_side.O_2_12\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_side.O_2_11\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_side.O_2_10\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_side.O_2_9\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_side.O_2_8\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_side.O_2_7\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_side.O_2_6\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_side.O_2_5\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_side.O_2_4\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(4);
    \pid_front.un2_error_1_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_front.un2_error_1_mulonly_0_24_0_A_wire\ <= \N__39452\&\N__39494\&\N__38961\&\N__38993\&\N__39047\&\N__39095\&\N__39155\&\N__39206\&\N__39266\&\N__39327\&\N__38630\&\N__38684\&\N__38747\&\N__38795\&\N__38849\&\N__38916\;
    \pid_front.un2_error_1_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_front.un2_error_1_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__55395\&\N__55605\&\N__55773\&\N__53253\&\N__55230\&\N__55950\&\N__56163\&\N__56334\;
    \pid_front.O_24\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(24);
    \pid_front.O_23\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(23);
    \pid_front.O_22\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(22);
    \pid_front.O_21\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(21);
    \pid_front.O_20\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(20);
    \pid_front.O_19\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(19);
    \pid_front.O_18\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(18);
    \pid_front.O_17\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(17);
    \pid_front.O_16\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(16);
    \pid_front.O_15\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(15);
    \pid_front.O_14\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(14);
    \pid_front.O_13\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(13);
    \pid_front.O_12\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(12);
    \pid_front.O_11\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(11);
    \pid_front.O_10\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(10);
    \pid_front.O_9\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(9);
    \pid_front.O_8\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(8);
    \pid_front.O_7\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(7);
    \pid_front.O_6\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(6);
    \pid_front.O_5\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(5);
    \pid_front.O_4\ <= \pid_front.un2_error_1_mulonly_0_24_0_O_wire\(4);

    \Pc2drone_pll_inst.Pc2drone_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => OPEN,
            SDI => \GNDG0\,
            BYPASS => \GNDG0\,
            RESETB => \N__42457\,
            PLLOUTCORE => \Pc2drone_pll_inst.clk_system_pll\,
            LOCK => OPEN,
            SDO => OPEN,
            SCLK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            EXTFEEDBACK => \GNDG0\,
            DYNAMICDELAY => \Pc2drone_pll_inst.Pc2drone_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__59697\
        );

    \pid_alt.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42363\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42326\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un2_error_1_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42230\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42229\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un2_error_2_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42287\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42286\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\
        );

    \pid_front.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42288\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42237\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_front.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_front.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_front.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_front.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_front.un2_error_mulonly_0_24_0_O_wire\
        );

    \pid_side.un2_error_1_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42458\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42432\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_side.un2_error_1_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_side.un2_error_1_mulonly_0_24_0_A_wire\,
            C => \pid_side.un2_error_1_mulonly_0_24_0_C_wire\,
            B => \pid_side.un2_error_1_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_side.un2_error_1_mulonly_0_24_0_O_wire\
        );

    \pid_side.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42228\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42392\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_side.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_side.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_side.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_side.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_side.un2_error_mulonly_0_24_0_O_wire\
        );

    \pid_front.un2_error_1_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__42459\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__42285\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_front.un2_error_1_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_front.un2_error_1_mulonly_0_24_0_A_wire\,
            C => \pid_front.un2_error_1_mulonly_0_24_0_C_wire\,
            B => \pid_front.un2_error_1_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_front.un2_error_1_mulonly_0_24_0_O_wire\
        );

    \Pc2drone_pll_inst.Pc2drone_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__59697\,
            PACKAGEPIN => clk_system_wire
        );

    \uart_input_pc_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59683\,
            DIN => \N__59682\,
            DOUT => \N__59681\,
            PACKAGEPIN => uart_input_pc_wire
        );

    \uart_input_pc_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__59683\,
            PADOUT => \N__59682\,
            PADIN => \N__59681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_pc_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH2_18A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59674\,
            DIN => \N__59673\,
            DOUT => \N__59672\,
            PACKAGEPIN => \debug_CH2_18A_wire\
        );

    \debug_CH2_18A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59674\,
            PADOUT => \N__59673\,
            PADIN => \N__59672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30354\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH0_16A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59665\,
            DIN => \N__59664\,
            DOUT => \N__59663\,
            PACKAGEPIN => \debug_CH0_16A_wire\
        );

    \debug_CH0_16A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59665\,
            PADOUT => \N__59664\,
            PADIN => \N__59663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32904\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH1_0A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59656\,
            DIN => \N__59655\,
            DOUT => \N__59654\,
            PACKAGEPIN => \debug_CH1_0A_wire\
        );

    \debug_CH1_0A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59656\,
            PADOUT => \N__59655\,
            PADIN => \N__59654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__47715\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH5_31B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59647\,
            DIN => \N__59646\,
            DOUT => \N__59645\,
            PACKAGEPIN => \debug_CH5_31B_wire\
        );

    \debug_CH5_31B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59647\,
            PADOUT => \N__59646\,
            PADIN => \N__59645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH4_2A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59638\,
            DIN => \N__59637\,
            DOUT => \N__59636\,
            PACKAGEPIN => \debug_CH4_2A_wire\
        );

    \debug_CH4_2A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59638\,
            PADOUT => \N__59637\,
            PADIN => \N__59636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ppm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59629\,
            DIN => \N__59628\,
            DOUT => \N__59627\,
            PACKAGEPIN => ppm_output_wire
        );

    \ppm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59629\,
            PADOUT => \N__59628\,
            PADIN => \N__59627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37641\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH3_20A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59620\,
            DIN => \N__59619\,
            DOUT => \N__59618\,
            PACKAGEPIN => \debug_CH3_20A_wire\
        );

    \debug_CH3_20A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59620\,
            PADOUT => \N__59619\,
            PADIN => \N__59618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__41031\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH6_5B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59611\,
            DIN => \N__59610\,
            DOUT => \N__59609\,
            PACKAGEPIN => \debug_CH6_5B_wire\
        );

    \debug_CH6_5B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__59611\,
            PADOUT => \N__59610\,
            PADIN => \N__59609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_drone_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59602\,
            DIN => \N__59601\,
            DOUT => \N__59600\,
            PACKAGEPIN => uart_input_drone_wire
        );

    \uart_input_drone_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__59602\,
            PADOUT => \N__59601\,
            PADIN => \N__59600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_drone_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__14335\ : InMux
    port map (
            O => \N__59583\,
            I => \N__59580\
        );

    \I__14334\ : LocalMux
    port map (
            O => \N__59580\,
            I => \N__59577\
        );

    \I__14333\ : Odrv4
    port map (
            O => \N__59577\,
            I => \pid_front.O_22\
        );

    \I__14332\ : InMux
    port map (
            O => \N__59574\,
            I => \N__59569\
        );

    \I__14331\ : InMux
    port map (
            O => \N__59573\,
            I => \N__59566\
        );

    \I__14330\ : InMux
    port map (
            O => \N__59572\,
            I => \N__59563\
        );

    \I__14329\ : LocalMux
    port map (
            O => \N__59569\,
            I => \N__59560\
        );

    \I__14328\ : LocalMux
    port map (
            O => \N__59566\,
            I => \N__59557\
        );

    \I__14327\ : LocalMux
    port map (
            O => \N__59563\,
            I => \N__59554\
        );

    \I__14326\ : Span12Mux_h
    port map (
            O => \N__59560\,
            I => \N__59551\
        );

    \I__14325\ : Span12Mux_v
    port map (
            O => \N__59557\,
            I => \N__59546\
        );

    \I__14324\ : Span12Mux_h
    port map (
            O => \N__59554\,
            I => \N__59546\
        );

    \I__14323\ : Span12Mux_h
    port map (
            O => \N__59551\,
            I => \N__59543\
        );

    \I__14322\ : Odrv12
    port map (
            O => \N__59546\,
            I => \pid_front.error_d_regZ0Z_18\
        );

    \I__14321\ : Odrv12
    port map (
            O => \N__59543\,
            I => \pid_front.error_d_regZ0Z_18\
        );

    \I__14320\ : InMux
    port map (
            O => \N__59538\,
            I => \N__59535\
        );

    \I__14319\ : LocalMux
    port map (
            O => \N__59535\,
            I => \N__59532\
        );

    \I__14318\ : Odrv4
    port map (
            O => \N__59532\,
            I => \pid_front.O_23\
        );

    \I__14317\ : InMux
    port map (
            O => \N__59529\,
            I => \N__59520\
        );

    \I__14316\ : InMux
    port map (
            O => \N__59528\,
            I => \N__59520\
        );

    \I__14315\ : InMux
    port map (
            O => \N__59527\,
            I => \N__59520\
        );

    \I__14314\ : LocalMux
    port map (
            O => \N__59520\,
            I => \N__59517\
        );

    \I__14313\ : Span12Mux_h
    port map (
            O => \N__59517\,
            I => \N__59514\
        );

    \I__14312\ : Odrv12
    port map (
            O => \N__59514\,
            I => \pid_front.error_d_regZ0Z_19\
        );

    \I__14311\ : InMux
    port map (
            O => \N__59511\,
            I => \N__59508\
        );

    \I__14310\ : LocalMux
    port map (
            O => \N__59508\,
            I => \N__59505\
        );

    \I__14309\ : Odrv4
    port map (
            O => \N__59505\,
            I => \pid_front.O_24\
        );

    \I__14308\ : InMux
    port map (
            O => \N__59502\,
            I => \N__59497\
        );

    \I__14307\ : InMux
    port map (
            O => \N__59501\,
            I => \N__59492\
        );

    \I__14306\ : InMux
    port map (
            O => \N__59500\,
            I => \N__59492\
        );

    \I__14305\ : LocalMux
    port map (
            O => \N__59497\,
            I => \N__59487\
        );

    \I__14304\ : LocalMux
    port map (
            O => \N__59492\,
            I => \N__59487\
        );

    \I__14303\ : Span4Mux_h
    port map (
            O => \N__59487\,
            I => \N__59484\
        );

    \I__14302\ : Span4Mux_h
    port map (
            O => \N__59484\,
            I => \N__59481\
        );

    \I__14301\ : Span4Mux_h
    port map (
            O => \N__59481\,
            I => \N__59478\
        );

    \I__14300\ : Odrv4
    port map (
            O => \N__59478\,
            I => \pid_front.error_d_regZ0Z_20\
        );

    \I__14299\ : InMux
    port map (
            O => \N__59475\,
            I => \N__59472\
        );

    \I__14298\ : LocalMux
    port map (
            O => \N__59472\,
            I => \N__59469\
        );

    \I__14297\ : Odrv4
    port map (
            O => \N__59469\,
            I => \pid_front.O_18\
        );

    \I__14296\ : InMux
    port map (
            O => \N__59466\,
            I => \N__59463\
        );

    \I__14295\ : LocalMux
    port map (
            O => \N__59463\,
            I => \N__59460\
        );

    \I__14294\ : Span4Mux_v
    port map (
            O => \N__59460\,
            I => \N__59455\
        );

    \I__14293\ : InMux
    port map (
            O => \N__59459\,
            I => \N__59452\
        );

    \I__14292\ : InMux
    port map (
            O => \N__59458\,
            I => \N__59449\
        );

    \I__14291\ : Span4Mux_h
    port map (
            O => \N__59455\,
            I => \N__59446\
        );

    \I__14290\ : LocalMux
    port map (
            O => \N__59452\,
            I => \N__59443\
        );

    \I__14289\ : LocalMux
    port map (
            O => \N__59449\,
            I => \N__59436\
        );

    \I__14288\ : Sp12to4
    port map (
            O => \N__59446\,
            I => \N__59436\
        );

    \I__14287\ : Span12Mux_h
    port map (
            O => \N__59443\,
            I => \N__59436\
        );

    \I__14286\ : Odrv12
    port map (
            O => \N__59436\,
            I => \pid_front.error_d_regZ0Z_14\
        );

    \I__14285\ : InMux
    port map (
            O => \N__59433\,
            I => \N__59430\
        );

    \I__14284\ : LocalMux
    port map (
            O => \N__59430\,
            I => \pid_front.O_8\
        );

    \I__14283\ : InMux
    port map (
            O => \N__59427\,
            I => \N__59418\
        );

    \I__14282\ : InMux
    port map (
            O => \N__59426\,
            I => \N__59418\
        );

    \I__14281\ : InMux
    port map (
            O => \N__59425\,
            I => \N__59418\
        );

    \I__14280\ : LocalMux
    port map (
            O => \N__59418\,
            I => \N__59415\
        );

    \I__14279\ : Span4Mux_h
    port map (
            O => \N__59415\,
            I => \N__59412\
        );

    \I__14278\ : Span4Mux_h
    port map (
            O => \N__59412\,
            I => \N__59409\
        );

    \I__14277\ : Span4Mux_h
    port map (
            O => \N__59409\,
            I => \N__59406\
        );

    \I__14276\ : Odrv4
    port map (
            O => \N__59406\,
            I => \pid_front.error_d_regZ0Z_4\
        );

    \I__14275\ : InMux
    port map (
            O => \N__59403\,
            I => \N__59400\
        );

    \I__14274\ : LocalMux
    port map (
            O => \N__59400\,
            I => \pid_front.O_11\
        );

    \I__14273\ : InMux
    port map (
            O => \N__59397\,
            I => \N__59392\
        );

    \I__14272\ : InMux
    port map (
            O => \N__59396\,
            I => \N__59387\
        );

    \I__14271\ : InMux
    port map (
            O => \N__59395\,
            I => \N__59387\
        );

    \I__14270\ : LocalMux
    port map (
            O => \N__59392\,
            I => \N__59382\
        );

    \I__14269\ : LocalMux
    port map (
            O => \N__59387\,
            I => \N__59382\
        );

    \I__14268\ : Span4Mux_h
    port map (
            O => \N__59382\,
            I => \N__59379\
        );

    \I__14267\ : Span4Mux_h
    port map (
            O => \N__59379\,
            I => \N__59376\
        );

    \I__14266\ : Span4Mux_h
    port map (
            O => \N__59376\,
            I => \N__59373\
        );

    \I__14265\ : Span4Mux_h
    port map (
            O => \N__59373\,
            I => \N__59370\
        );

    \I__14264\ : Odrv4
    port map (
            O => \N__59370\,
            I => \pid_front.error_d_regZ0Z_7\
        );

    \I__14263\ : InMux
    port map (
            O => \N__59367\,
            I => \N__59364\
        );

    \I__14262\ : LocalMux
    port map (
            O => \N__59364\,
            I => \pid_front.O_19\
        );

    \I__14261\ : InMux
    port map (
            O => \N__59361\,
            I => \N__59352\
        );

    \I__14260\ : InMux
    port map (
            O => \N__59360\,
            I => \N__59352\
        );

    \I__14259\ : InMux
    port map (
            O => \N__59359\,
            I => \N__59352\
        );

    \I__14258\ : LocalMux
    port map (
            O => \N__59352\,
            I => \N__59349\
        );

    \I__14257\ : Span4Mux_v
    port map (
            O => \N__59349\,
            I => \N__59346\
        );

    \I__14256\ : Sp12to4
    port map (
            O => \N__59346\,
            I => \N__59343\
        );

    \I__14255\ : Span12Mux_h
    port map (
            O => \N__59343\,
            I => \N__59340\
        );

    \I__14254\ : Odrv12
    port map (
            O => \N__59340\,
            I => \pid_front.error_d_regZ0Z_15\
        );

    \I__14253\ : ClkMux
    port map (
            O => \N__59337\,
            I => \N__58545\
        );

    \I__14252\ : ClkMux
    port map (
            O => \N__59336\,
            I => \N__58545\
        );

    \I__14251\ : ClkMux
    port map (
            O => \N__59335\,
            I => \N__58545\
        );

    \I__14250\ : ClkMux
    port map (
            O => \N__59334\,
            I => \N__58545\
        );

    \I__14249\ : ClkMux
    port map (
            O => \N__59333\,
            I => \N__58545\
        );

    \I__14248\ : ClkMux
    port map (
            O => \N__59332\,
            I => \N__58545\
        );

    \I__14247\ : ClkMux
    port map (
            O => \N__59331\,
            I => \N__58545\
        );

    \I__14246\ : ClkMux
    port map (
            O => \N__59330\,
            I => \N__58545\
        );

    \I__14245\ : ClkMux
    port map (
            O => \N__59329\,
            I => \N__58545\
        );

    \I__14244\ : ClkMux
    port map (
            O => \N__59328\,
            I => \N__58545\
        );

    \I__14243\ : ClkMux
    port map (
            O => \N__59327\,
            I => \N__58545\
        );

    \I__14242\ : ClkMux
    port map (
            O => \N__59326\,
            I => \N__58545\
        );

    \I__14241\ : ClkMux
    port map (
            O => \N__59325\,
            I => \N__58545\
        );

    \I__14240\ : ClkMux
    port map (
            O => \N__59324\,
            I => \N__58545\
        );

    \I__14239\ : ClkMux
    port map (
            O => \N__59323\,
            I => \N__58545\
        );

    \I__14238\ : ClkMux
    port map (
            O => \N__59322\,
            I => \N__58545\
        );

    \I__14237\ : ClkMux
    port map (
            O => \N__59321\,
            I => \N__58545\
        );

    \I__14236\ : ClkMux
    port map (
            O => \N__59320\,
            I => \N__58545\
        );

    \I__14235\ : ClkMux
    port map (
            O => \N__59319\,
            I => \N__58545\
        );

    \I__14234\ : ClkMux
    port map (
            O => \N__59318\,
            I => \N__58545\
        );

    \I__14233\ : ClkMux
    port map (
            O => \N__59317\,
            I => \N__58545\
        );

    \I__14232\ : ClkMux
    port map (
            O => \N__59316\,
            I => \N__58545\
        );

    \I__14231\ : ClkMux
    port map (
            O => \N__59315\,
            I => \N__58545\
        );

    \I__14230\ : ClkMux
    port map (
            O => \N__59314\,
            I => \N__58545\
        );

    \I__14229\ : ClkMux
    port map (
            O => \N__59313\,
            I => \N__58545\
        );

    \I__14228\ : ClkMux
    port map (
            O => \N__59312\,
            I => \N__58545\
        );

    \I__14227\ : ClkMux
    port map (
            O => \N__59311\,
            I => \N__58545\
        );

    \I__14226\ : ClkMux
    port map (
            O => \N__59310\,
            I => \N__58545\
        );

    \I__14225\ : ClkMux
    port map (
            O => \N__59309\,
            I => \N__58545\
        );

    \I__14224\ : ClkMux
    port map (
            O => \N__59308\,
            I => \N__58545\
        );

    \I__14223\ : ClkMux
    port map (
            O => \N__59307\,
            I => \N__58545\
        );

    \I__14222\ : ClkMux
    port map (
            O => \N__59306\,
            I => \N__58545\
        );

    \I__14221\ : ClkMux
    port map (
            O => \N__59305\,
            I => \N__58545\
        );

    \I__14220\ : ClkMux
    port map (
            O => \N__59304\,
            I => \N__58545\
        );

    \I__14219\ : ClkMux
    port map (
            O => \N__59303\,
            I => \N__58545\
        );

    \I__14218\ : ClkMux
    port map (
            O => \N__59302\,
            I => \N__58545\
        );

    \I__14217\ : ClkMux
    port map (
            O => \N__59301\,
            I => \N__58545\
        );

    \I__14216\ : ClkMux
    port map (
            O => \N__59300\,
            I => \N__58545\
        );

    \I__14215\ : ClkMux
    port map (
            O => \N__59299\,
            I => \N__58545\
        );

    \I__14214\ : ClkMux
    port map (
            O => \N__59298\,
            I => \N__58545\
        );

    \I__14213\ : ClkMux
    port map (
            O => \N__59297\,
            I => \N__58545\
        );

    \I__14212\ : ClkMux
    port map (
            O => \N__59296\,
            I => \N__58545\
        );

    \I__14211\ : ClkMux
    port map (
            O => \N__59295\,
            I => \N__58545\
        );

    \I__14210\ : ClkMux
    port map (
            O => \N__59294\,
            I => \N__58545\
        );

    \I__14209\ : ClkMux
    port map (
            O => \N__59293\,
            I => \N__58545\
        );

    \I__14208\ : ClkMux
    port map (
            O => \N__59292\,
            I => \N__58545\
        );

    \I__14207\ : ClkMux
    port map (
            O => \N__59291\,
            I => \N__58545\
        );

    \I__14206\ : ClkMux
    port map (
            O => \N__59290\,
            I => \N__58545\
        );

    \I__14205\ : ClkMux
    port map (
            O => \N__59289\,
            I => \N__58545\
        );

    \I__14204\ : ClkMux
    port map (
            O => \N__59288\,
            I => \N__58545\
        );

    \I__14203\ : ClkMux
    port map (
            O => \N__59287\,
            I => \N__58545\
        );

    \I__14202\ : ClkMux
    port map (
            O => \N__59286\,
            I => \N__58545\
        );

    \I__14201\ : ClkMux
    port map (
            O => \N__59285\,
            I => \N__58545\
        );

    \I__14200\ : ClkMux
    port map (
            O => \N__59284\,
            I => \N__58545\
        );

    \I__14199\ : ClkMux
    port map (
            O => \N__59283\,
            I => \N__58545\
        );

    \I__14198\ : ClkMux
    port map (
            O => \N__59282\,
            I => \N__58545\
        );

    \I__14197\ : ClkMux
    port map (
            O => \N__59281\,
            I => \N__58545\
        );

    \I__14196\ : ClkMux
    port map (
            O => \N__59280\,
            I => \N__58545\
        );

    \I__14195\ : ClkMux
    port map (
            O => \N__59279\,
            I => \N__58545\
        );

    \I__14194\ : ClkMux
    port map (
            O => \N__59278\,
            I => \N__58545\
        );

    \I__14193\ : ClkMux
    port map (
            O => \N__59277\,
            I => \N__58545\
        );

    \I__14192\ : ClkMux
    port map (
            O => \N__59276\,
            I => \N__58545\
        );

    \I__14191\ : ClkMux
    port map (
            O => \N__59275\,
            I => \N__58545\
        );

    \I__14190\ : ClkMux
    port map (
            O => \N__59274\,
            I => \N__58545\
        );

    \I__14189\ : ClkMux
    port map (
            O => \N__59273\,
            I => \N__58545\
        );

    \I__14188\ : ClkMux
    port map (
            O => \N__59272\,
            I => \N__58545\
        );

    \I__14187\ : ClkMux
    port map (
            O => \N__59271\,
            I => \N__58545\
        );

    \I__14186\ : ClkMux
    port map (
            O => \N__59270\,
            I => \N__58545\
        );

    \I__14185\ : ClkMux
    port map (
            O => \N__59269\,
            I => \N__58545\
        );

    \I__14184\ : ClkMux
    port map (
            O => \N__59268\,
            I => \N__58545\
        );

    \I__14183\ : ClkMux
    port map (
            O => \N__59267\,
            I => \N__58545\
        );

    \I__14182\ : ClkMux
    port map (
            O => \N__59266\,
            I => \N__58545\
        );

    \I__14181\ : ClkMux
    port map (
            O => \N__59265\,
            I => \N__58545\
        );

    \I__14180\ : ClkMux
    port map (
            O => \N__59264\,
            I => \N__58545\
        );

    \I__14179\ : ClkMux
    port map (
            O => \N__59263\,
            I => \N__58545\
        );

    \I__14178\ : ClkMux
    port map (
            O => \N__59262\,
            I => \N__58545\
        );

    \I__14177\ : ClkMux
    port map (
            O => \N__59261\,
            I => \N__58545\
        );

    \I__14176\ : ClkMux
    port map (
            O => \N__59260\,
            I => \N__58545\
        );

    \I__14175\ : ClkMux
    port map (
            O => \N__59259\,
            I => \N__58545\
        );

    \I__14174\ : ClkMux
    port map (
            O => \N__59258\,
            I => \N__58545\
        );

    \I__14173\ : ClkMux
    port map (
            O => \N__59257\,
            I => \N__58545\
        );

    \I__14172\ : ClkMux
    port map (
            O => \N__59256\,
            I => \N__58545\
        );

    \I__14171\ : ClkMux
    port map (
            O => \N__59255\,
            I => \N__58545\
        );

    \I__14170\ : ClkMux
    port map (
            O => \N__59254\,
            I => \N__58545\
        );

    \I__14169\ : ClkMux
    port map (
            O => \N__59253\,
            I => \N__58545\
        );

    \I__14168\ : ClkMux
    port map (
            O => \N__59252\,
            I => \N__58545\
        );

    \I__14167\ : ClkMux
    port map (
            O => \N__59251\,
            I => \N__58545\
        );

    \I__14166\ : ClkMux
    port map (
            O => \N__59250\,
            I => \N__58545\
        );

    \I__14165\ : ClkMux
    port map (
            O => \N__59249\,
            I => \N__58545\
        );

    \I__14164\ : ClkMux
    port map (
            O => \N__59248\,
            I => \N__58545\
        );

    \I__14163\ : ClkMux
    port map (
            O => \N__59247\,
            I => \N__58545\
        );

    \I__14162\ : ClkMux
    port map (
            O => \N__59246\,
            I => \N__58545\
        );

    \I__14161\ : ClkMux
    port map (
            O => \N__59245\,
            I => \N__58545\
        );

    \I__14160\ : ClkMux
    port map (
            O => \N__59244\,
            I => \N__58545\
        );

    \I__14159\ : ClkMux
    port map (
            O => \N__59243\,
            I => \N__58545\
        );

    \I__14158\ : ClkMux
    port map (
            O => \N__59242\,
            I => \N__58545\
        );

    \I__14157\ : ClkMux
    port map (
            O => \N__59241\,
            I => \N__58545\
        );

    \I__14156\ : ClkMux
    port map (
            O => \N__59240\,
            I => \N__58545\
        );

    \I__14155\ : ClkMux
    port map (
            O => \N__59239\,
            I => \N__58545\
        );

    \I__14154\ : ClkMux
    port map (
            O => \N__59238\,
            I => \N__58545\
        );

    \I__14153\ : ClkMux
    port map (
            O => \N__59237\,
            I => \N__58545\
        );

    \I__14152\ : ClkMux
    port map (
            O => \N__59236\,
            I => \N__58545\
        );

    \I__14151\ : ClkMux
    port map (
            O => \N__59235\,
            I => \N__58545\
        );

    \I__14150\ : ClkMux
    port map (
            O => \N__59234\,
            I => \N__58545\
        );

    \I__14149\ : ClkMux
    port map (
            O => \N__59233\,
            I => \N__58545\
        );

    \I__14148\ : ClkMux
    port map (
            O => \N__59232\,
            I => \N__58545\
        );

    \I__14147\ : ClkMux
    port map (
            O => \N__59231\,
            I => \N__58545\
        );

    \I__14146\ : ClkMux
    port map (
            O => \N__59230\,
            I => \N__58545\
        );

    \I__14145\ : ClkMux
    port map (
            O => \N__59229\,
            I => \N__58545\
        );

    \I__14144\ : ClkMux
    port map (
            O => \N__59228\,
            I => \N__58545\
        );

    \I__14143\ : ClkMux
    port map (
            O => \N__59227\,
            I => \N__58545\
        );

    \I__14142\ : ClkMux
    port map (
            O => \N__59226\,
            I => \N__58545\
        );

    \I__14141\ : ClkMux
    port map (
            O => \N__59225\,
            I => \N__58545\
        );

    \I__14140\ : ClkMux
    port map (
            O => \N__59224\,
            I => \N__58545\
        );

    \I__14139\ : ClkMux
    port map (
            O => \N__59223\,
            I => \N__58545\
        );

    \I__14138\ : ClkMux
    port map (
            O => \N__59222\,
            I => \N__58545\
        );

    \I__14137\ : ClkMux
    port map (
            O => \N__59221\,
            I => \N__58545\
        );

    \I__14136\ : ClkMux
    port map (
            O => \N__59220\,
            I => \N__58545\
        );

    \I__14135\ : ClkMux
    port map (
            O => \N__59219\,
            I => \N__58545\
        );

    \I__14134\ : ClkMux
    port map (
            O => \N__59218\,
            I => \N__58545\
        );

    \I__14133\ : ClkMux
    port map (
            O => \N__59217\,
            I => \N__58545\
        );

    \I__14132\ : ClkMux
    port map (
            O => \N__59216\,
            I => \N__58545\
        );

    \I__14131\ : ClkMux
    port map (
            O => \N__59215\,
            I => \N__58545\
        );

    \I__14130\ : ClkMux
    port map (
            O => \N__59214\,
            I => \N__58545\
        );

    \I__14129\ : ClkMux
    port map (
            O => \N__59213\,
            I => \N__58545\
        );

    \I__14128\ : ClkMux
    port map (
            O => \N__59212\,
            I => \N__58545\
        );

    \I__14127\ : ClkMux
    port map (
            O => \N__59211\,
            I => \N__58545\
        );

    \I__14126\ : ClkMux
    port map (
            O => \N__59210\,
            I => \N__58545\
        );

    \I__14125\ : ClkMux
    port map (
            O => \N__59209\,
            I => \N__58545\
        );

    \I__14124\ : ClkMux
    port map (
            O => \N__59208\,
            I => \N__58545\
        );

    \I__14123\ : ClkMux
    port map (
            O => \N__59207\,
            I => \N__58545\
        );

    \I__14122\ : ClkMux
    port map (
            O => \N__59206\,
            I => \N__58545\
        );

    \I__14121\ : ClkMux
    port map (
            O => \N__59205\,
            I => \N__58545\
        );

    \I__14120\ : ClkMux
    port map (
            O => \N__59204\,
            I => \N__58545\
        );

    \I__14119\ : ClkMux
    port map (
            O => \N__59203\,
            I => \N__58545\
        );

    \I__14118\ : ClkMux
    port map (
            O => \N__59202\,
            I => \N__58545\
        );

    \I__14117\ : ClkMux
    port map (
            O => \N__59201\,
            I => \N__58545\
        );

    \I__14116\ : ClkMux
    port map (
            O => \N__59200\,
            I => \N__58545\
        );

    \I__14115\ : ClkMux
    port map (
            O => \N__59199\,
            I => \N__58545\
        );

    \I__14114\ : ClkMux
    port map (
            O => \N__59198\,
            I => \N__58545\
        );

    \I__14113\ : ClkMux
    port map (
            O => \N__59197\,
            I => \N__58545\
        );

    \I__14112\ : ClkMux
    port map (
            O => \N__59196\,
            I => \N__58545\
        );

    \I__14111\ : ClkMux
    port map (
            O => \N__59195\,
            I => \N__58545\
        );

    \I__14110\ : ClkMux
    port map (
            O => \N__59194\,
            I => \N__58545\
        );

    \I__14109\ : ClkMux
    port map (
            O => \N__59193\,
            I => \N__58545\
        );

    \I__14108\ : ClkMux
    port map (
            O => \N__59192\,
            I => \N__58545\
        );

    \I__14107\ : ClkMux
    port map (
            O => \N__59191\,
            I => \N__58545\
        );

    \I__14106\ : ClkMux
    port map (
            O => \N__59190\,
            I => \N__58545\
        );

    \I__14105\ : ClkMux
    port map (
            O => \N__59189\,
            I => \N__58545\
        );

    \I__14104\ : ClkMux
    port map (
            O => \N__59188\,
            I => \N__58545\
        );

    \I__14103\ : ClkMux
    port map (
            O => \N__59187\,
            I => \N__58545\
        );

    \I__14102\ : ClkMux
    port map (
            O => \N__59186\,
            I => \N__58545\
        );

    \I__14101\ : ClkMux
    port map (
            O => \N__59185\,
            I => \N__58545\
        );

    \I__14100\ : ClkMux
    port map (
            O => \N__59184\,
            I => \N__58545\
        );

    \I__14099\ : ClkMux
    port map (
            O => \N__59183\,
            I => \N__58545\
        );

    \I__14098\ : ClkMux
    port map (
            O => \N__59182\,
            I => \N__58545\
        );

    \I__14097\ : ClkMux
    port map (
            O => \N__59181\,
            I => \N__58545\
        );

    \I__14096\ : ClkMux
    port map (
            O => \N__59180\,
            I => \N__58545\
        );

    \I__14095\ : ClkMux
    port map (
            O => \N__59179\,
            I => \N__58545\
        );

    \I__14094\ : ClkMux
    port map (
            O => \N__59178\,
            I => \N__58545\
        );

    \I__14093\ : ClkMux
    port map (
            O => \N__59177\,
            I => \N__58545\
        );

    \I__14092\ : ClkMux
    port map (
            O => \N__59176\,
            I => \N__58545\
        );

    \I__14091\ : ClkMux
    port map (
            O => \N__59175\,
            I => \N__58545\
        );

    \I__14090\ : ClkMux
    port map (
            O => \N__59174\,
            I => \N__58545\
        );

    \I__14089\ : ClkMux
    port map (
            O => \N__59173\,
            I => \N__58545\
        );

    \I__14088\ : ClkMux
    port map (
            O => \N__59172\,
            I => \N__58545\
        );

    \I__14087\ : ClkMux
    port map (
            O => \N__59171\,
            I => \N__58545\
        );

    \I__14086\ : ClkMux
    port map (
            O => \N__59170\,
            I => \N__58545\
        );

    \I__14085\ : ClkMux
    port map (
            O => \N__59169\,
            I => \N__58545\
        );

    \I__14084\ : ClkMux
    port map (
            O => \N__59168\,
            I => \N__58545\
        );

    \I__14083\ : ClkMux
    port map (
            O => \N__59167\,
            I => \N__58545\
        );

    \I__14082\ : ClkMux
    port map (
            O => \N__59166\,
            I => \N__58545\
        );

    \I__14081\ : ClkMux
    port map (
            O => \N__59165\,
            I => \N__58545\
        );

    \I__14080\ : ClkMux
    port map (
            O => \N__59164\,
            I => \N__58545\
        );

    \I__14079\ : ClkMux
    port map (
            O => \N__59163\,
            I => \N__58545\
        );

    \I__14078\ : ClkMux
    port map (
            O => \N__59162\,
            I => \N__58545\
        );

    \I__14077\ : ClkMux
    port map (
            O => \N__59161\,
            I => \N__58545\
        );

    \I__14076\ : ClkMux
    port map (
            O => \N__59160\,
            I => \N__58545\
        );

    \I__14075\ : ClkMux
    port map (
            O => \N__59159\,
            I => \N__58545\
        );

    \I__14074\ : ClkMux
    port map (
            O => \N__59158\,
            I => \N__58545\
        );

    \I__14073\ : ClkMux
    port map (
            O => \N__59157\,
            I => \N__58545\
        );

    \I__14072\ : ClkMux
    port map (
            O => \N__59156\,
            I => \N__58545\
        );

    \I__14071\ : ClkMux
    port map (
            O => \N__59155\,
            I => \N__58545\
        );

    \I__14070\ : ClkMux
    port map (
            O => \N__59154\,
            I => \N__58545\
        );

    \I__14069\ : ClkMux
    port map (
            O => \N__59153\,
            I => \N__58545\
        );

    \I__14068\ : ClkMux
    port map (
            O => \N__59152\,
            I => \N__58545\
        );

    \I__14067\ : ClkMux
    port map (
            O => \N__59151\,
            I => \N__58545\
        );

    \I__14066\ : ClkMux
    port map (
            O => \N__59150\,
            I => \N__58545\
        );

    \I__14065\ : ClkMux
    port map (
            O => \N__59149\,
            I => \N__58545\
        );

    \I__14064\ : ClkMux
    port map (
            O => \N__59148\,
            I => \N__58545\
        );

    \I__14063\ : ClkMux
    port map (
            O => \N__59147\,
            I => \N__58545\
        );

    \I__14062\ : ClkMux
    port map (
            O => \N__59146\,
            I => \N__58545\
        );

    \I__14061\ : ClkMux
    port map (
            O => \N__59145\,
            I => \N__58545\
        );

    \I__14060\ : ClkMux
    port map (
            O => \N__59144\,
            I => \N__58545\
        );

    \I__14059\ : ClkMux
    port map (
            O => \N__59143\,
            I => \N__58545\
        );

    \I__14058\ : ClkMux
    port map (
            O => \N__59142\,
            I => \N__58545\
        );

    \I__14057\ : ClkMux
    port map (
            O => \N__59141\,
            I => \N__58545\
        );

    \I__14056\ : ClkMux
    port map (
            O => \N__59140\,
            I => \N__58545\
        );

    \I__14055\ : ClkMux
    port map (
            O => \N__59139\,
            I => \N__58545\
        );

    \I__14054\ : ClkMux
    port map (
            O => \N__59138\,
            I => \N__58545\
        );

    \I__14053\ : ClkMux
    port map (
            O => \N__59137\,
            I => \N__58545\
        );

    \I__14052\ : ClkMux
    port map (
            O => \N__59136\,
            I => \N__58545\
        );

    \I__14051\ : ClkMux
    port map (
            O => \N__59135\,
            I => \N__58545\
        );

    \I__14050\ : ClkMux
    port map (
            O => \N__59134\,
            I => \N__58545\
        );

    \I__14049\ : ClkMux
    port map (
            O => \N__59133\,
            I => \N__58545\
        );

    \I__14048\ : ClkMux
    port map (
            O => \N__59132\,
            I => \N__58545\
        );

    \I__14047\ : ClkMux
    port map (
            O => \N__59131\,
            I => \N__58545\
        );

    \I__14046\ : ClkMux
    port map (
            O => \N__59130\,
            I => \N__58545\
        );

    \I__14045\ : ClkMux
    port map (
            O => \N__59129\,
            I => \N__58545\
        );

    \I__14044\ : ClkMux
    port map (
            O => \N__59128\,
            I => \N__58545\
        );

    \I__14043\ : ClkMux
    port map (
            O => \N__59127\,
            I => \N__58545\
        );

    \I__14042\ : ClkMux
    port map (
            O => \N__59126\,
            I => \N__58545\
        );

    \I__14041\ : ClkMux
    port map (
            O => \N__59125\,
            I => \N__58545\
        );

    \I__14040\ : ClkMux
    port map (
            O => \N__59124\,
            I => \N__58545\
        );

    \I__14039\ : ClkMux
    port map (
            O => \N__59123\,
            I => \N__58545\
        );

    \I__14038\ : ClkMux
    port map (
            O => \N__59122\,
            I => \N__58545\
        );

    \I__14037\ : ClkMux
    port map (
            O => \N__59121\,
            I => \N__58545\
        );

    \I__14036\ : ClkMux
    port map (
            O => \N__59120\,
            I => \N__58545\
        );

    \I__14035\ : ClkMux
    port map (
            O => \N__59119\,
            I => \N__58545\
        );

    \I__14034\ : ClkMux
    port map (
            O => \N__59118\,
            I => \N__58545\
        );

    \I__14033\ : ClkMux
    port map (
            O => \N__59117\,
            I => \N__58545\
        );

    \I__14032\ : ClkMux
    port map (
            O => \N__59116\,
            I => \N__58545\
        );

    \I__14031\ : ClkMux
    port map (
            O => \N__59115\,
            I => \N__58545\
        );

    \I__14030\ : ClkMux
    port map (
            O => \N__59114\,
            I => \N__58545\
        );

    \I__14029\ : ClkMux
    port map (
            O => \N__59113\,
            I => \N__58545\
        );

    \I__14028\ : ClkMux
    port map (
            O => \N__59112\,
            I => \N__58545\
        );

    \I__14027\ : ClkMux
    port map (
            O => \N__59111\,
            I => \N__58545\
        );

    \I__14026\ : ClkMux
    port map (
            O => \N__59110\,
            I => \N__58545\
        );

    \I__14025\ : ClkMux
    port map (
            O => \N__59109\,
            I => \N__58545\
        );

    \I__14024\ : ClkMux
    port map (
            O => \N__59108\,
            I => \N__58545\
        );

    \I__14023\ : ClkMux
    port map (
            O => \N__59107\,
            I => \N__58545\
        );

    \I__14022\ : ClkMux
    port map (
            O => \N__59106\,
            I => \N__58545\
        );

    \I__14021\ : ClkMux
    port map (
            O => \N__59105\,
            I => \N__58545\
        );

    \I__14020\ : ClkMux
    port map (
            O => \N__59104\,
            I => \N__58545\
        );

    \I__14019\ : ClkMux
    port map (
            O => \N__59103\,
            I => \N__58545\
        );

    \I__14018\ : ClkMux
    port map (
            O => \N__59102\,
            I => \N__58545\
        );

    \I__14017\ : ClkMux
    port map (
            O => \N__59101\,
            I => \N__58545\
        );

    \I__14016\ : ClkMux
    port map (
            O => \N__59100\,
            I => \N__58545\
        );

    \I__14015\ : ClkMux
    port map (
            O => \N__59099\,
            I => \N__58545\
        );

    \I__14014\ : ClkMux
    port map (
            O => \N__59098\,
            I => \N__58545\
        );

    \I__14013\ : ClkMux
    port map (
            O => \N__59097\,
            I => \N__58545\
        );

    \I__14012\ : ClkMux
    port map (
            O => \N__59096\,
            I => \N__58545\
        );

    \I__14011\ : ClkMux
    port map (
            O => \N__59095\,
            I => \N__58545\
        );

    \I__14010\ : ClkMux
    port map (
            O => \N__59094\,
            I => \N__58545\
        );

    \I__14009\ : ClkMux
    port map (
            O => \N__59093\,
            I => \N__58545\
        );

    \I__14008\ : ClkMux
    port map (
            O => \N__59092\,
            I => \N__58545\
        );

    \I__14007\ : ClkMux
    port map (
            O => \N__59091\,
            I => \N__58545\
        );

    \I__14006\ : ClkMux
    port map (
            O => \N__59090\,
            I => \N__58545\
        );

    \I__14005\ : ClkMux
    port map (
            O => \N__59089\,
            I => \N__58545\
        );

    \I__14004\ : ClkMux
    port map (
            O => \N__59088\,
            I => \N__58545\
        );

    \I__14003\ : ClkMux
    port map (
            O => \N__59087\,
            I => \N__58545\
        );

    \I__14002\ : ClkMux
    port map (
            O => \N__59086\,
            I => \N__58545\
        );

    \I__14001\ : ClkMux
    port map (
            O => \N__59085\,
            I => \N__58545\
        );

    \I__14000\ : ClkMux
    port map (
            O => \N__59084\,
            I => \N__58545\
        );

    \I__13999\ : ClkMux
    port map (
            O => \N__59083\,
            I => \N__58545\
        );

    \I__13998\ : ClkMux
    port map (
            O => \N__59082\,
            I => \N__58545\
        );

    \I__13997\ : ClkMux
    port map (
            O => \N__59081\,
            I => \N__58545\
        );

    \I__13996\ : ClkMux
    port map (
            O => \N__59080\,
            I => \N__58545\
        );

    \I__13995\ : ClkMux
    port map (
            O => \N__59079\,
            I => \N__58545\
        );

    \I__13994\ : ClkMux
    port map (
            O => \N__59078\,
            I => \N__58545\
        );

    \I__13993\ : ClkMux
    port map (
            O => \N__59077\,
            I => \N__58545\
        );

    \I__13992\ : ClkMux
    port map (
            O => \N__59076\,
            I => \N__58545\
        );

    \I__13991\ : ClkMux
    port map (
            O => \N__59075\,
            I => \N__58545\
        );

    \I__13990\ : ClkMux
    port map (
            O => \N__59074\,
            I => \N__58545\
        );

    \I__13989\ : GlobalMux
    port map (
            O => \N__58545\,
            I => \N__58542\
        );

    \I__13988\ : gio2CtrlBuf
    port map (
            O => \N__58542\,
            I => clk_system_pll_g
        );

    \I__13987\ : CEMux
    port map (
            O => \N__58539\,
            I => \N__58531\
        );

    \I__13986\ : CEMux
    port map (
            O => \N__58538\,
            I => \N__58528\
        );

    \I__13985\ : CEMux
    port map (
            O => \N__58537\,
            I => \N__58525\
        );

    \I__13984\ : CEMux
    port map (
            O => \N__58536\,
            I => \N__58520\
        );

    \I__13983\ : CEMux
    port map (
            O => \N__58535\,
            I => \N__58517\
        );

    \I__13982\ : CEMux
    port map (
            O => \N__58534\,
            I => \N__58514\
        );

    \I__13981\ : LocalMux
    port map (
            O => \N__58531\,
            I => \N__58511\
        );

    \I__13980\ : LocalMux
    port map (
            O => \N__58528\,
            I => \N__58508\
        );

    \I__13979\ : LocalMux
    port map (
            O => \N__58525\,
            I => \N__58504\
        );

    \I__13978\ : CEMux
    port map (
            O => \N__58524\,
            I => \N__58499\
        );

    \I__13977\ : CEMux
    port map (
            O => \N__58523\,
            I => \N__58496\
        );

    \I__13976\ : LocalMux
    port map (
            O => \N__58520\,
            I => \N__58491\
        );

    \I__13975\ : LocalMux
    port map (
            O => \N__58517\,
            I => \N__58486\
        );

    \I__13974\ : LocalMux
    port map (
            O => \N__58514\,
            I => \N__58486\
        );

    \I__13973\ : Span4Mux_v
    port map (
            O => \N__58511\,
            I => \N__58483\
        );

    \I__13972\ : Span4Mux_s3_h
    port map (
            O => \N__58508\,
            I => \N__58480\
        );

    \I__13971\ : CEMux
    port map (
            O => \N__58507\,
            I => \N__58477\
        );

    \I__13970\ : Span4Mux_s3_h
    port map (
            O => \N__58504\,
            I => \N__58474\
        );

    \I__13969\ : CEMux
    port map (
            O => \N__58503\,
            I => \N__58471\
        );

    \I__13968\ : CEMux
    port map (
            O => \N__58502\,
            I => \N__58468\
        );

    \I__13967\ : LocalMux
    port map (
            O => \N__58499\,
            I => \N__58465\
        );

    \I__13966\ : LocalMux
    port map (
            O => \N__58496\,
            I => \N__58462\
        );

    \I__13965\ : CEMux
    port map (
            O => \N__58495\,
            I => \N__58459\
        );

    \I__13964\ : CEMux
    port map (
            O => \N__58494\,
            I => \N__58456\
        );

    \I__13963\ : Span4Mux_s1_h
    port map (
            O => \N__58491\,
            I => \N__58450\
        );

    \I__13962\ : Span4Mux_v
    port map (
            O => \N__58486\,
            I => \N__58450\
        );

    \I__13961\ : Span4Mux_v
    port map (
            O => \N__58483\,
            I => \N__58446\
        );

    \I__13960\ : Span4Mux_v
    port map (
            O => \N__58480\,
            I => \N__58443\
        );

    \I__13959\ : LocalMux
    port map (
            O => \N__58477\,
            I => \N__58440\
        );

    \I__13958\ : Span4Mux_h
    port map (
            O => \N__58474\,
            I => \N__58435\
        );

    \I__13957\ : LocalMux
    port map (
            O => \N__58471\,
            I => \N__58435\
        );

    \I__13956\ : LocalMux
    port map (
            O => \N__58468\,
            I => \N__58432\
        );

    \I__13955\ : Span4Mux_s2_h
    port map (
            O => \N__58465\,
            I => \N__58423\
        );

    \I__13954\ : Span4Mux_s2_h
    port map (
            O => \N__58462\,
            I => \N__58423\
        );

    \I__13953\ : LocalMux
    port map (
            O => \N__58459\,
            I => \N__58423\
        );

    \I__13952\ : LocalMux
    port map (
            O => \N__58456\,
            I => \N__58423\
        );

    \I__13951\ : CEMux
    port map (
            O => \N__58455\,
            I => \N__58420\
        );

    \I__13950\ : Span4Mux_h
    port map (
            O => \N__58450\,
            I => \N__58417\
        );

    \I__13949\ : CEMux
    port map (
            O => \N__58449\,
            I => \N__58414\
        );

    \I__13948\ : Span4Mux_h
    port map (
            O => \N__58446\,
            I => \N__58411\
        );

    \I__13947\ : Span4Mux_h
    port map (
            O => \N__58443\,
            I => \N__58408\
        );

    \I__13946\ : Span4Mux_h
    port map (
            O => \N__58440\,
            I => \N__58405\
        );

    \I__13945\ : Span4Mux_h
    port map (
            O => \N__58435\,
            I => \N__58402\
        );

    \I__13944\ : Span4Mux_h
    port map (
            O => \N__58432\,
            I => \N__58395\
        );

    \I__13943\ : Span4Mux_h
    port map (
            O => \N__58423\,
            I => \N__58395\
        );

    \I__13942\ : LocalMux
    port map (
            O => \N__58420\,
            I => \N__58395\
        );

    \I__13941\ : Span4Mux_h
    port map (
            O => \N__58417\,
            I => \N__58392\
        );

    \I__13940\ : LocalMux
    port map (
            O => \N__58414\,
            I => \N__58389\
        );

    \I__13939\ : Span4Mux_h
    port map (
            O => \N__58411\,
            I => \N__58386\
        );

    \I__13938\ : Span4Mux_h
    port map (
            O => \N__58408\,
            I => \N__58383\
        );

    \I__13937\ : Span4Mux_v
    port map (
            O => \N__58405\,
            I => \N__58378\
        );

    \I__13936\ : Span4Mux_v
    port map (
            O => \N__58402\,
            I => \N__58378\
        );

    \I__13935\ : Span4Mux_h
    port map (
            O => \N__58395\,
            I => \N__58375\
        );

    \I__13934\ : Span4Mux_h
    port map (
            O => \N__58392\,
            I => \N__58370\
        );

    \I__13933\ : Span4Mux_h
    port map (
            O => \N__58389\,
            I => \N__58370\
        );

    \I__13932\ : Odrv4
    port map (
            O => \N__58386\,
            I => \pid_front.N_543_0\
        );

    \I__13931\ : Odrv4
    port map (
            O => \N__58383\,
            I => \pid_front.N_543_0\
        );

    \I__13930\ : Odrv4
    port map (
            O => \N__58378\,
            I => \pid_front.N_543_0\
        );

    \I__13929\ : Odrv4
    port map (
            O => \N__58375\,
            I => \pid_front.N_543_0\
        );

    \I__13928\ : Odrv4
    port map (
            O => \N__58370\,
            I => \pid_front.N_543_0\
        );

    \I__13927\ : InMux
    port map (
            O => \N__58359\,
            I => \N__58314\
        );

    \I__13926\ : InMux
    port map (
            O => \N__58358\,
            I => \N__58314\
        );

    \I__13925\ : InMux
    port map (
            O => \N__58357\,
            I => \N__58305\
        );

    \I__13924\ : InMux
    port map (
            O => \N__58356\,
            I => \N__58305\
        );

    \I__13923\ : InMux
    port map (
            O => \N__58355\,
            I => \N__58305\
        );

    \I__13922\ : InMux
    port map (
            O => \N__58354\,
            I => \N__58305\
        );

    \I__13921\ : InMux
    port map (
            O => \N__58353\,
            I => \N__58300\
        );

    \I__13920\ : InMux
    port map (
            O => \N__58352\,
            I => \N__58300\
        );

    \I__13919\ : InMux
    port map (
            O => \N__58351\,
            I => \N__58295\
        );

    \I__13918\ : InMux
    port map (
            O => \N__58350\,
            I => \N__58295\
        );

    \I__13917\ : InMux
    port map (
            O => \N__58349\,
            I => \N__58286\
        );

    \I__13916\ : InMux
    port map (
            O => \N__58348\,
            I => \N__58286\
        );

    \I__13915\ : InMux
    port map (
            O => \N__58347\,
            I => \N__58286\
        );

    \I__13914\ : InMux
    port map (
            O => \N__58346\,
            I => \N__58286\
        );

    \I__13913\ : InMux
    port map (
            O => \N__58345\,
            I => \N__58281\
        );

    \I__13912\ : InMux
    port map (
            O => \N__58344\,
            I => \N__58281\
        );

    \I__13911\ : InMux
    port map (
            O => \N__58343\,
            I => \N__58276\
        );

    \I__13910\ : InMux
    port map (
            O => \N__58342\,
            I => \N__58276\
        );

    \I__13909\ : InMux
    port map (
            O => \N__58341\,
            I => \N__58265\
        );

    \I__13908\ : InMux
    port map (
            O => \N__58340\,
            I => \N__58265\
        );

    \I__13907\ : InMux
    port map (
            O => \N__58339\,
            I => \N__58265\
        );

    \I__13906\ : InMux
    port map (
            O => \N__58338\,
            I => \N__58265\
        );

    \I__13905\ : InMux
    port map (
            O => \N__58337\,
            I => \N__58265\
        );

    \I__13904\ : InMux
    port map (
            O => \N__58336\,
            I => \N__58262\
        );

    \I__13903\ : InMux
    port map (
            O => \N__58335\,
            I => \N__58257\
        );

    \I__13902\ : InMux
    port map (
            O => \N__58334\,
            I => \N__58257\
        );

    \I__13901\ : InMux
    port map (
            O => \N__58333\,
            I => \N__58252\
        );

    \I__13900\ : InMux
    port map (
            O => \N__58332\,
            I => \N__58252\
        );

    \I__13899\ : InMux
    port map (
            O => \N__58331\,
            I => \N__58247\
        );

    \I__13898\ : InMux
    port map (
            O => \N__58330\,
            I => \N__58247\
        );

    \I__13897\ : InMux
    port map (
            O => \N__58329\,
            I => \N__58232\
        );

    \I__13896\ : InMux
    port map (
            O => \N__58328\,
            I => \N__58232\
        );

    \I__13895\ : InMux
    port map (
            O => \N__58327\,
            I => \N__58232\
        );

    \I__13894\ : InMux
    port map (
            O => \N__58326\,
            I => \N__58232\
        );

    \I__13893\ : InMux
    port map (
            O => \N__58325\,
            I => \N__58232\
        );

    \I__13892\ : InMux
    port map (
            O => \N__58324\,
            I => \N__58232\
        );

    \I__13891\ : InMux
    port map (
            O => \N__58323\,
            I => \N__58232\
        );

    \I__13890\ : InMux
    port map (
            O => \N__58322\,
            I => \N__58229\
        );

    \I__13889\ : InMux
    port map (
            O => \N__58321\,
            I => \N__58226\
        );

    \I__13888\ : InMux
    port map (
            O => \N__58320\,
            I => \N__58223\
        );

    \I__13887\ : InMux
    port map (
            O => \N__58319\,
            I => \N__58220\
        );

    \I__13886\ : LocalMux
    port map (
            O => \N__58314\,
            I => \N__58176\
        );

    \I__13885\ : LocalMux
    port map (
            O => \N__58305\,
            I => \N__58173\
        );

    \I__13884\ : LocalMux
    port map (
            O => \N__58300\,
            I => \N__58170\
        );

    \I__13883\ : LocalMux
    port map (
            O => \N__58295\,
            I => \N__58167\
        );

    \I__13882\ : LocalMux
    port map (
            O => \N__58286\,
            I => \N__58164\
        );

    \I__13881\ : LocalMux
    port map (
            O => \N__58281\,
            I => \N__58161\
        );

    \I__13880\ : LocalMux
    port map (
            O => \N__58276\,
            I => \N__58158\
        );

    \I__13879\ : LocalMux
    port map (
            O => \N__58265\,
            I => \N__58155\
        );

    \I__13878\ : LocalMux
    port map (
            O => \N__58262\,
            I => \N__58152\
        );

    \I__13877\ : LocalMux
    port map (
            O => \N__58257\,
            I => \N__58149\
        );

    \I__13876\ : LocalMux
    port map (
            O => \N__58252\,
            I => \N__58146\
        );

    \I__13875\ : LocalMux
    port map (
            O => \N__58247\,
            I => \N__58143\
        );

    \I__13874\ : LocalMux
    port map (
            O => \N__58232\,
            I => \N__58140\
        );

    \I__13873\ : LocalMux
    port map (
            O => \N__58229\,
            I => \N__58137\
        );

    \I__13872\ : LocalMux
    port map (
            O => \N__58226\,
            I => \N__58134\
        );

    \I__13871\ : LocalMux
    port map (
            O => \N__58223\,
            I => \N__58131\
        );

    \I__13870\ : LocalMux
    port map (
            O => \N__58220\,
            I => \N__58128\
        );

    \I__13869\ : SRMux
    port map (
            O => \N__58219\,
            I => \N__58011\
        );

    \I__13868\ : SRMux
    port map (
            O => \N__58218\,
            I => \N__58011\
        );

    \I__13867\ : SRMux
    port map (
            O => \N__58217\,
            I => \N__58011\
        );

    \I__13866\ : SRMux
    port map (
            O => \N__58216\,
            I => \N__58011\
        );

    \I__13865\ : SRMux
    port map (
            O => \N__58215\,
            I => \N__58011\
        );

    \I__13864\ : SRMux
    port map (
            O => \N__58214\,
            I => \N__58011\
        );

    \I__13863\ : SRMux
    port map (
            O => \N__58213\,
            I => \N__58011\
        );

    \I__13862\ : SRMux
    port map (
            O => \N__58212\,
            I => \N__58011\
        );

    \I__13861\ : SRMux
    port map (
            O => \N__58211\,
            I => \N__58011\
        );

    \I__13860\ : SRMux
    port map (
            O => \N__58210\,
            I => \N__58011\
        );

    \I__13859\ : SRMux
    port map (
            O => \N__58209\,
            I => \N__58011\
        );

    \I__13858\ : SRMux
    port map (
            O => \N__58208\,
            I => \N__58011\
        );

    \I__13857\ : SRMux
    port map (
            O => \N__58207\,
            I => \N__58011\
        );

    \I__13856\ : SRMux
    port map (
            O => \N__58206\,
            I => \N__58011\
        );

    \I__13855\ : SRMux
    port map (
            O => \N__58205\,
            I => \N__58011\
        );

    \I__13854\ : SRMux
    port map (
            O => \N__58204\,
            I => \N__58011\
        );

    \I__13853\ : SRMux
    port map (
            O => \N__58203\,
            I => \N__58011\
        );

    \I__13852\ : SRMux
    port map (
            O => \N__58202\,
            I => \N__58011\
        );

    \I__13851\ : SRMux
    port map (
            O => \N__58201\,
            I => \N__58011\
        );

    \I__13850\ : SRMux
    port map (
            O => \N__58200\,
            I => \N__58011\
        );

    \I__13849\ : SRMux
    port map (
            O => \N__58199\,
            I => \N__58011\
        );

    \I__13848\ : SRMux
    port map (
            O => \N__58198\,
            I => \N__58011\
        );

    \I__13847\ : SRMux
    port map (
            O => \N__58197\,
            I => \N__58011\
        );

    \I__13846\ : SRMux
    port map (
            O => \N__58196\,
            I => \N__58011\
        );

    \I__13845\ : SRMux
    port map (
            O => \N__58195\,
            I => \N__58011\
        );

    \I__13844\ : SRMux
    port map (
            O => \N__58194\,
            I => \N__58011\
        );

    \I__13843\ : SRMux
    port map (
            O => \N__58193\,
            I => \N__58011\
        );

    \I__13842\ : SRMux
    port map (
            O => \N__58192\,
            I => \N__58011\
        );

    \I__13841\ : SRMux
    port map (
            O => \N__58191\,
            I => \N__58011\
        );

    \I__13840\ : SRMux
    port map (
            O => \N__58190\,
            I => \N__58011\
        );

    \I__13839\ : SRMux
    port map (
            O => \N__58189\,
            I => \N__58011\
        );

    \I__13838\ : SRMux
    port map (
            O => \N__58188\,
            I => \N__58011\
        );

    \I__13837\ : SRMux
    port map (
            O => \N__58187\,
            I => \N__58011\
        );

    \I__13836\ : SRMux
    port map (
            O => \N__58186\,
            I => \N__58011\
        );

    \I__13835\ : SRMux
    port map (
            O => \N__58185\,
            I => \N__58011\
        );

    \I__13834\ : SRMux
    port map (
            O => \N__58184\,
            I => \N__58011\
        );

    \I__13833\ : SRMux
    port map (
            O => \N__58183\,
            I => \N__58011\
        );

    \I__13832\ : SRMux
    port map (
            O => \N__58182\,
            I => \N__58011\
        );

    \I__13831\ : SRMux
    port map (
            O => \N__58181\,
            I => \N__58011\
        );

    \I__13830\ : SRMux
    port map (
            O => \N__58180\,
            I => \N__58011\
        );

    \I__13829\ : SRMux
    port map (
            O => \N__58179\,
            I => \N__58011\
        );

    \I__13828\ : Glb2LocalMux
    port map (
            O => \N__58176\,
            I => \N__58011\
        );

    \I__13827\ : Glb2LocalMux
    port map (
            O => \N__58173\,
            I => \N__58011\
        );

    \I__13826\ : Glb2LocalMux
    port map (
            O => \N__58170\,
            I => \N__58011\
        );

    \I__13825\ : Glb2LocalMux
    port map (
            O => \N__58167\,
            I => \N__58011\
        );

    \I__13824\ : Glb2LocalMux
    port map (
            O => \N__58164\,
            I => \N__58011\
        );

    \I__13823\ : Glb2LocalMux
    port map (
            O => \N__58161\,
            I => \N__58011\
        );

    \I__13822\ : Glb2LocalMux
    port map (
            O => \N__58158\,
            I => \N__58011\
        );

    \I__13821\ : Glb2LocalMux
    port map (
            O => \N__58155\,
            I => \N__58011\
        );

    \I__13820\ : Glb2LocalMux
    port map (
            O => \N__58152\,
            I => \N__58011\
        );

    \I__13819\ : Glb2LocalMux
    port map (
            O => \N__58149\,
            I => \N__58011\
        );

    \I__13818\ : Glb2LocalMux
    port map (
            O => \N__58146\,
            I => \N__58011\
        );

    \I__13817\ : Glb2LocalMux
    port map (
            O => \N__58143\,
            I => \N__58011\
        );

    \I__13816\ : Glb2LocalMux
    port map (
            O => \N__58140\,
            I => \N__58011\
        );

    \I__13815\ : Glb2LocalMux
    port map (
            O => \N__58137\,
            I => \N__58011\
        );

    \I__13814\ : Glb2LocalMux
    port map (
            O => \N__58134\,
            I => \N__58011\
        );

    \I__13813\ : Glb2LocalMux
    port map (
            O => \N__58131\,
            I => \N__58011\
        );

    \I__13812\ : Glb2LocalMux
    port map (
            O => \N__58128\,
            I => \N__58011\
        );

    \I__13811\ : GlobalMux
    port map (
            O => \N__58011\,
            I => \N__58008\
        );

    \I__13810\ : gio2CtrlBuf
    port map (
            O => \N__58008\,
            I => \N_665_g\
        );

    \I__13809\ : InMux
    port map (
            O => \N__58005\,
            I => \N__58001\
        );

    \I__13808\ : InMux
    port map (
            O => \N__58004\,
            I => \N__57998\
        );

    \I__13807\ : LocalMux
    port map (
            O => \N__58001\,
            I => \N__57994\
        );

    \I__13806\ : LocalMux
    port map (
            O => \N__57998\,
            I => \N__57991\
        );

    \I__13805\ : InMux
    port map (
            O => \N__57997\,
            I => \N__57988\
        );

    \I__13804\ : Odrv12
    port map (
            O => \N__57994\,
            I => \pid_side.error_d_regZ0Z_20\
        );

    \I__13803\ : Odrv4
    port map (
            O => \N__57991\,
            I => \pid_side.error_d_regZ0Z_20\
        );

    \I__13802\ : LocalMux
    port map (
            O => \N__57988\,
            I => \pid_side.error_d_regZ0Z_20\
        );

    \I__13801\ : InMux
    port map (
            O => \N__57981\,
            I => \N__57977\
        );

    \I__13800\ : InMux
    port map (
            O => \N__57980\,
            I => \N__57974\
        );

    \I__13799\ : LocalMux
    port map (
            O => \N__57977\,
            I => \N__57969\
        );

    \I__13798\ : LocalMux
    port map (
            O => \N__57974\,
            I => \N__57969\
        );

    \I__13797\ : Odrv4
    port map (
            O => \N__57969\,
            I => \pid_side.error_d_reg_prevZ0Z_20\
        );

    \I__13796\ : CEMux
    port map (
            O => \N__57966\,
            I => \N__57909\
        );

    \I__13795\ : CEMux
    port map (
            O => \N__57965\,
            I => \N__57909\
        );

    \I__13794\ : CEMux
    port map (
            O => \N__57964\,
            I => \N__57909\
        );

    \I__13793\ : CEMux
    port map (
            O => \N__57963\,
            I => \N__57909\
        );

    \I__13792\ : CEMux
    port map (
            O => \N__57962\,
            I => \N__57909\
        );

    \I__13791\ : CEMux
    port map (
            O => \N__57961\,
            I => \N__57909\
        );

    \I__13790\ : CEMux
    port map (
            O => \N__57960\,
            I => \N__57909\
        );

    \I__13789\ : CEMux
    port map (
            O => \N__57959\,
            I => \N__57909\
        );

    \I__13788\ : CEMux
    port map (
            O => \N__57958\,
            I => \N__57909\
        );

    \I__13787\ : CEMux
    port map (
            O => \N__57957\,
            I => \N__57909\
        );

    \I__13786\ : CEMux
    port map (
            O => \N__57956\,
            I => \N__57909\
        );

    \I__13785\ : CEMux
    port map (
            O => \N__57955\,
            I => \N__57909\
        );

    \I__13784\ : CEMux
    port map (
            O => \N__57954\,
            I => \N__57909\
        );

    \I__13783\ : CEMux
    port map (
            O => \N__57953\,
            I => \N__57909\
        );

    \I__13782\ : CEMux
    port map (
            O => \N__57952\,
            I => \N__57909\
        );

    \I__13781\ : CEMux
    port map (
            O => \N__57951\,
            I => \N__57909\
        );

    \I__13780\ : CEMux
    port map (
            O => \N__57950\,
            I => \N__57909\
        );

    \I__13779\ : CEMux
    port map (
            O => \N__57949\,
            I => \N__57909\
        );

    \I__13778\ : CEMux
    port map (
            O => \N__57948\,
            I => \N__57909\
        );

    \I__13777\ : GlobalMux
    port map (
            O => \N__57909\,
            I => \N__57906\
        );

    \I__13776\ : gio2CtrlBuf
    port map (
            O => \N__57906\,
            I => \pid_side.state_0_g_0\
        );

    \I__13775\ : CascadeMux
    port map (
            O => \N__57903\,
            I => \N__57897\
        );

    \I__13774\ : CascadeMux
    port map (
            O => \N__57902\,
            I => \N__57891\
        );

    \I__13773\ : CascadeMux
    port map (
            O => \N__57901\,
            I => \N__57872\
        );

    \I__13772\ : CascadeMux
    port map (
            O => \N__57900\,
            I => \N__57838\
        );

    \I__13771\ : InMux
    port map (
            O => \N__57897\,
            I => \N__57824\
        );

    \I__13770\ : InMux
    port map (
            O => \N__57896\,
            I => \N__57821\
        );

    \I__13769\ : InMux
    port map (
            O => \N__57895\,
            I => \N__57818\
        );

    \I__13768\ : InMux
    port map (
            O => \N__57894\,
            I => \N__57811\
        );

    \I__13767\ : InMux
    port map (
            O => \N__57891\,
            I => \N__57811\
        );

    \I__13766\ : InMux
    port map (
            O => \N__57890\,
            I => \N__57811\
        );

    \I__13765\ : InMux
    port map (
            O => \N__57889\,
            I => \N__57808\
        );

    \I__13764\ : InMux
    port map (
            O => \N__57888\,
            I => \N__57799\
        );

    \I__13763\ : InMux
    port map (
            O => \N__57887\,
            I => \N__57799\
        );

    \I__13762\ : InMux
    port map (
            O => \N__57886\,
            I => \N__57799\
        );

    \I__13761\ : InMux
    port map (
            O => \N__57885\,
            I => \N__57799\
        );

    \I__13760\ : InMux
    port map (
            O => \N__57884\,
            I => \N__57794\
        );

    \I__13759\ : InMux
    port map (
            O => \N__57883\,
            I => \N__57794\
        );

    \I__13758\ : InMux
    port map (
            O => \N__57882\,
            I => \N__57787\
        );

    \I__13757\ : InMux
    port map (
            O => \N__57881\,
            I => \N__57787\
        );

    \I__13756\ : InMux
    port map (
            O => \N__57880\,
            I => \N__57787\
        );

    \I__13755\ : InMux
    port map (
            O => \N__57879\,
            I => \N__57782\
        );

    \I__13754\ : InMux
    port map (
            O => \N__57878\,
            I => \N__57782\
        );

    \I__13753\ : InMux
    port map (
            O => \N__57877\,
            I => \N__57775\
        );

    \I__13752\ : InMux
    port map (
            O => \N__57876\,
            I => \N__57775\
        );

    \I__13751\ : InMux
    port map (
            O => \N__57875\,
            I => \N__57775\
        );

    \I__13750\ : InMux
    port map (
            O => \N__57872\,
            I => \N__57770\
        );

    \I__13749\ : InMux
    port map (
            O => \N__57871\,
            I => \N__57770\
        );

    \I__13748\ : InMux
    port map (
            O => \N__57870\,
            I => \N__57767\
        );

    \I__13747\ : InMux
    port map (
            O => \N__57869\,
            I => \N__57760\
        );

    \I__13746\ : InMux
    port map (
            O => \N__57868\,
            I => \N__57760\
        );

    \I__13745\ : InMux
    port map (
            O => \N__57867\,
            I => \N__57760\
        );

    \I__13744\ : InMux
    port map (
            O => \N__57866\,
            I => \N__57757\
        );

    \I__13743\ : InMux
    port map (
            O => \N__57865\,
            I => \N__57754\
        );

    \I__13742\ : InMux
    port map (
            O => \N__57864\,
            I => \N__57751\
        );

    \I__13741\ : InMux
    port map (
            O => \N__57863\,
            I => \N__57746\
        );

    \I__13740\ : InMux
    port map (
            O => \N__57862\,
            I => \N__57746\
        );

    \I__13739\ : InMux
    port map (
            O => \N__57861\,
            I => \N__57743\
        );

    \I__13738\ : InMux
    port map (
            O => \N__57860\,
            I => \N__57740\
        );

    \I__13737\ : InMux
    port map (
            O => \N__57859\,
            I => \N__57737\
        );

    \I__13736\ : InMux
    port map (
            O => \N__57858\,
            I => \N__57734\
        );

    \I__13735\ : InMux
    port map (
            O => \N__57857\,
            I => \N__57727\
        );

    \I__13734\ : InMux
    port map (
            O => \N__57856\,
            I => \N__57727\
        );

    \I__13733\ : InMux
    port map (
            O => \N__57855\,
            I => \N__57727\
        );

    \I__13732\ : InMux
    port map (
            O => \N__57854\,
            I => \N__57724\
        );

    \I__13731\ : InMux
    port map (
            O => \N__57853\,
            I => \N__57719\
        );

    \I__13730\ : InMux
    port map (
            O => \N__57852\,
            I => \N__57719\
        );

    \I__13729\ : InMux
    port map (
            O => \N__57851\,
            I => \N__57716\
        );

    \I__13728\ : InMux
    port map (
            O => \N__57850\,
            I => \N__57713\
        );

    \I__13727\ : InMux
    port map (
            O => \N__57849\,
            I => \N__57710\
        );

    \I__13726\ : InMux
    port map (
            O => \N__57848\,
            I => \N__57707\
        );

    \I__13725\ : InMux
    port map (
            O => \N__57847\,
            I => \N__57704\
        );

    \I__13724\ : InMux
    port map (
            O => \N__57846\,
            I => \N__57701\
        );

    \I__13723\ : InMux
    port map (
            O => \N__57845\,
            I => \N__57698\
        );

    \I__13722\ : InMux
    port map (
            O => \N__57844\,
            I => \N__57695\
        );

    \I__13721\ : InMux
    port map (
            O => \N__57843\,
            I => \N__57690\
        );

    \I__13720\ : InMux
    port map (
            O => \N__57842\,
            I => \N__57690\
        );

    \I__13719\ : InMux
    port map (
            O => \N__57841\,
            I => \N__57687\
        );

    \I__13718\ : InMux
    port map (
            O => \N__57838\,
            I => \N__57684\
        );

    \I__13717\ : InMux
    port map (
            O => \N__57837\,
            I => \N__57681\
        );

    \I__13716\ : InMux
    port map (
            O => \N__57836\,
            I => \N__57678\
        );

    \I__13715\ : InMux
    port map (
            O => \N__57835\,
            I => \N__57675\
        );

    \I__13714\ : InMux
    port map (
            O => \N__57834\,
            I => \N__57672\
        );

    \I__13713\ : InMux
    port map (
            O => \N__57833\,
            I => \N__57669\
        );

    \I__13712\ : InMux
    port map (
            O => \N__57832\,
            I => \N__57666\
        );

    \I__13711\ : InMux
    port map (
            O => \N__57831\,
            I => \N__57663\
        );

    \I__13710\ : InMux
    port map (
            O => \N__57830\,
            I => \N__57660\
        );

    \I__13709\ : InMux
    port map (
            O => \N__57829\,
            I => \N__57657\
        );

    \I__13708\ : InMux
    port map (
            O => \N__57828\,
            I => \N__57654\
        );

    \I__13707\ : InMux
    port map (
            O => \N__57827\,
            I => \N__57651\
        );

    \I__13706\ : LocalMux
    port map (
            O => \N__57824\,
            I => \N__57493\
        );

    \I__13705\ : LocalMux
    port map (
            O => \N__57821\,
            I => \N__57490\
        );

    \I__13704\ : LocalMux
    port map (
            O => \N__57818\,
            I => \N__57487\
        );

    \I__13703\ : LocalMux
    port map (
            O => \N__57811\,
            I => \N__57484\
        );

    \I__13702\ : LocalMux
    port map (
            O => \N__57808\,
            I => \N__57481\
        );

    \I__13701\ : LocalMux
    port map (
            O => \N__57799\,
            I => \N__57478\
        );

    \I__13700\ : LocalMux
    port map (
            O => \N__57794\,
            I => \N__57475\
        );

    \I__13699\ : LocalMux
    port map (
            O => \N__57787\,
            I => \N__57472\
        );

    \I__13698\ : LocalMux
    port map (
            O => \N__57782\,
            I => \N__57469\
        );

    \I__13697\ : LocalMux
    port map (
            O => \N__57775\,
            I => \N__57466\
        );

    \I__13696\ : LocalMux
    port map (
            O => \N__57770\,
            I => \N__57463\
        );

    \I__13695\ : LocalMux
    port map (
            O => \N__57767\,
            I => \N__57460\
        );

    \I__13694\ : LocalMux
    port map (
            O => \N__57760\,
            I => \N__57457\
        );

    \I__13693\ : LocalMux
    port map (
            O => \N__57757\,
            I => \N__57454\
        );

    \I__13692\ : LocalMux
    port map (
            O => \N__57754\,
            I => \N__57451\
        );

    \I__13691\ : LocalMux
    port map (
            O => \N__57751\,
            I => \N__57448\
        );

    \I__13690\ : LocalMux
    port map (
            O => \N__57746\,
            I => \N__57445\
        );

    \I__13689\ : LocalMux
    port map (
            O => \N__57743\,
            I => \N__57442\
        );

    \I__13688\ : LocalMux
    port map (
            O => \N__57740\,
            I => \N__57439\
        );

    \I__13687\ : LocalMux
    port map (
            O => \N__57737\,
            I => \N__57436\
        );

    \I__13686\ : LocalMux
    port map (
            O => \N__57734\,
            I => \N__57433\
        );

    \I__13685\ : LocalMux
    port map (
            O => \N__57727\,
            I => \N__57430\
        );

    \I__13684\ : LocalMux
    port map (
            O => \N__57724\,
            I => \N__57427\
        );

    \I__13683\ : LocalMux
    port map (
            O => \N__57719\,
            I => \N__57424\
        );

    \I__13682\ : LocalMux
    port map (
            O => \N__57716\,
            I => \N__57421\
        );

    \I__13681\ : LocalMux
    port map (
            O => \N__57713\,
            I => \N__57418\
        );

    \I__13680\ : LocalMux
    port map (
            O => \N__57710\,
            I => \N__57415\
        );

    \I__13679\ : LocalMux
    port map (
            O => \N__57707\,
            I => \N__57412\
        );

    \I__13678\ : LocalMux
    port map (
            O => \N__57704\,
            I => \N__57409\
        );

    \I__13677\ : LocalMux
    port map (
            O => \N__57701\,
            I => \N__57406\
        );

    \I__13676\ : LocalMux
    port map (
            O => \N__57698\,
            I => \N__57403\
        );

    \I__13675\ : LocalMux
    port map (
            O => \N__57695\,
            I => \N__57400\
        );

    \I__13674\ : LocalMux
    port map (
            O => \N__57690\,
            I => \N__57397\
        );

    \I__13673\ : LocalMux
    port map (
            O => \N__57687\,
            I => \N__57394\
        );

    \I__13672\ : LocalMux
    port map (
            O => \N__57684\,
            I => \N__57391\
        );

    \I__13671\ : LocalMux
    port map (
            O => \N__57681\,
            I => \N__57388\
        );

    \I__13670\ : LocalMux
    port map (
            O => \N__57678\,
            I => \N__57385\
        );

    \I__13669\ : LocalMux
    port map (
            O => \N__57675\,
            I => \N__57382\
        );

    \I__13668\ : LocalMux
    port map (
            O => \N__57672\,
            I => \N__57379\
        );

    \I__13667\ : LocalMux
    port map (
            O => \N__57669\,
            I => \N__57376\
        );

    \I__13666\ : LocalMux
    port map (
            O => \N__57666\,
            I => \N__57373\
        );

    \I__13665\ : LocalMux
    port map (
            O => \N__57663\,
            I => \N__57370\
        );

    \I__13664\ : LocalMux
    port map (
            O => \N__57660\,
            I => \N__57367\
        );

    \I__13663\ : LocalMux
    port map (
            O => \N__57657\,
            I => \N__57364\
        );

    \I__13662\ : LocalMux
    port map (
            O => \N__57654\,
            I => \N__57361\
        );

    \I__13661\ : LocalMux
    port map (
            O => \N__57651\,
            I => \N__57358\
        );

    \I__13660\ : SRMux
    port map (
            O => \N__57650\,
            I => \N__56955\
        );

    \I__13659\ : SRMux
    port map (
            O => \N__57649\,
            I => \N__56955\
        );

    \I__13658\ : SRMux
    port map (
            O => \N__57648\,
            I => \N__56955\
        );

    \I__13657\ : SRMux
    port map (
            O => \N__57647\,
            I => \N__56955\
        );

    \I__13656\ : SRMux
    port map (
            O => \N__57646\,
            I => \N__56955\
        );

    \I__13655\ : SRMux
    port map (
            O => \N__57645\,
            I => \N__56955\
        );

    \I__13654\ : SRMux
    port map (
            O => \N__57644\,
            I => \N__56955\
        );

    \I__13653\ : SRMux
    port map (
            O => \N__57643\,
            I => \N__56955\
        );

    \I__13652\ : SRMux
    port map (
            O => \N__57642\,
            I => \N__56955\
        );

    \I__13651\ : SRMux
    port map (
            O => \N__57641\,
            I => \N__56955\
        );

    \I__13650\ : SRMux
    port map (
            O => \N__57640\,
            I => \N__56955\
        );

    \I__13649\ : SRMux
    port map (
            O => \N__57639\,
            I => \N__56955\
        );

    \I__13648\ : SRMux
    port map (
            O => \N__57638\,
            I => \N__56955\
        );

    \I__13647\ : SRMux
    port map (
            O => \N__57637\,
            I => \N__56955\
        );

    \I__13646\ : SRMux
    port map (
            O => \N__57636\,
            I => \N__56955\
        );

    \I__13645\ : SRMux
    port map (
            O => \N__57635\,
            I => \N__56955\
        );

    \I__13644\ : SRMux
    port map (
            O => \N__57634\,
            I => \N__56955\
        );

    \I__13643\ : SRMux
    port map (
            O => \N__57633\,
            I => \N__56955\
        );

    \I__13642\ : SRMux
    port map (
            O => \N__57632\,
            I => \N__56955\
        );

    \I__13641\ : SRMux
    port map (
            O => \N__57631\,
            I => \N__56955\
        );

    \I__13640\ : SRMux
    port map (
            O => \N__57630\,
            I => \N__56955\
        );

    \I__13639\ : SRMux
    port map (
            O => \N__57629\,
            I => \N__56955\
        );

    \I__13638\ : SRMux
    port map (
            O => \N__57628\,
            I => \N__56955\
        );

    \I__13637\ : SRMux
    port map (
            O => \N__57627\,
            I => \N__56955\
        );

    \I__13636\ : SRMux
    port map (
            O => \N__57626\,
            I => \N__56955\
        );

    \I__13635\ : SRMux
    port map (
            O => \N__57625\,
            I => \N__56955\
        );

    \I__13634\ : SRMux
    port map (
            O => \N__57624\,
            I => \N__56955\
        );

    \I__13633\ : SRMux
    port map (
            O => \N__57623\,
            I => \N__56955\
        );

    \I__13632\ : SRMux
    port map (
            O => \N__57622\,
            I => \N__56955\
        );

    \I__13631\ : SRMux
    port map (
            O => \N__57621\,
            I => \N__56955\
        );

    \I__13630\ : SRMux
    port map (
            O => \N__57620\,
            I => \N__56955\
        );

    \I__13629\ : SRMux
    port map (
            O => \N__57619\,
            I => \N__56955\
        );

    \I__13628\ : SRMux
    port map (
            O => \N__57618\,
            I => \N__56955\
        );

    \I__13627\ : SRMux
    port map (
            O => \N__57617\,
            I => \N__56955\
        );

    \I__13626\ : SRMux
    port map (
            O => \N__57616\,
            I => \N__56955\
        );

    \I__13625\ : SRMux
    port map (
            O => \N__57615\,
            I => \N__56955\
        );

    \I__13624\ : SRMux
    port map (
            O => \N__57614\,
            I => \N__56955\
        );

    \I__13623\ : SRMux
    port map (
            O => \N__57613\,
            I => \N__56955\
        );

    \I__13622\ : SRMux
    port map (
            O => \N__57612\,
            I => \N__56955\
        );

    \I__13621\ : SRMux
    port map (
            O => \N__57611\,
            I => \N__56955\
        );

    \I__13620\ : SRMux
    port map (
            O => \N__57610\,
            I => \N__56955\
        );

    \I__13619\ : SRMux
    port map (
            O => \N__57609\,
            I => \N__56955\
        );

    \I__13618\ : SRMux
    port map (
            O => \N__57608\,
            I => \N__56955\
        );

    \I__13617\ : SRMux
    port map (
            O => \N__57607\,
            I => \N__56955\
        );

    \I__13616\ : SRMux
    port map (
            O => \N__57606\,
            I => \N__56955\
        );

    \I__13615\ : SRMux
    port map (
            O => \N__57605\,
            I => \N__56955\
        );

    \I__13614\ : SRMux
    port map (
            O => \N__57604\,
            I => \N__56955\
        );

    \I__13613\ : SRMux
    port map (
            O => \N__57603\,
            I => \N__56955\
        );

    \I__13612\ : SRMux
    port map (
            O => \N__57602\,
            I => \N__56955\
        );

    \I__13611\ : SRMux
    port map (
            O => \N__57601\,
            I => \N__56955\
        );

    \I__13610\ : SRMux
    port map (
            O => \N__57600\,
            I => \N__56955\
        );

    \I__13609\ : SRMux
    port map (
            O => \N__57599\,
            I => \N__56955\
        );

    \I__13608\ : SRMux
    port map (
            O => \N__57598\,
            I => \N__56955\
        );

    \I__13607\ : SRMux
    port map (
            O => \N__57597\,
            I => \N__56955\
        );

    \I__13606\ : SRMux
    port map (
            O => \N__57596\,
            I => \N__56955\
        );

    \I__13605\ : SRMux
    port map (
            O => \N__57595\,
            I => \N__56955\
        );

    \I__13604\ : SRMux
    port map (
            O => \N__57594\,
            I => \N__56955\
        );

    \I__13603\ : SRMux
    port map (
            O => \N__57593\,
            I => \N__56955\
        );

    \I__13602\ : SRMux
    port map (
            O => \N__57592\,
            I => \N__56955\
        );

    \I__13601\ : SRMux
    port map (
            O => \N__57591\,
            I => \N__56955\
        );

    \I__13600\ : SRMux
    port map (
            O => \N__57590\,
            I => \N__56955\
        );

    \I__13599\ : SRMux
    port map (
            O => \N__57589\,
            I => \N__56955\
        );

    \I__13598\ : SRMux
    port map (
            O => \N__57588\,
            I => \N__56955\
        );

    \I__13597\ : SRMux
    port map (
            O => \N__57587\,
            I => \N__56955\
        );

    \I__13596\ : SRMux
    port map (
            O => \N__57586\,
            I => \N__56955\
        );

    \I__13595\ : SRMux
    port map (
            O => \N__57585\,
            I => \N__56955\
        );

    \I__13594\ : SRMux
    port map (
            O => \N__57584\,
            I => \N__56955\
        );

    \I__13593\ : SRMux
    port map (
            O => \N__57583\,
            I => \N__56955\
        );

    \I__13592\ : SRMux
    port map (
            O => \N__57582\,
            I => \N__56955\
        );

    \I__13591\ : SRMux
    port map (
            O => \N__57581\,
            I => \N__56955\
        );

    \I__13590\ : SRMux
    port map (
            O => \N__57580\,
            I => \N__56955\
        );

    \I__13589\ : SRMux
    port map (
            O => \N__57579\,
            I => \N__56955\
        );

    \I__13588\ : SRMux
    port map (
            O => \N__57578\,
            I => \N__56955\
        );

    \I__13587\ : SRMux
    port map (
            O => \N__57577\,
            I => \N__56955\
        );

    \I__13586\ : SRMux
    port map (
            O => \N__57576\,
            I => \N__56955\
        );

    \I__13585\ : SRMux
    port map (
            O => \N__57575\,
            I => \N__56955\
        );

    \I__13584\ : SRMux
    port map (
            O => \N__57574\,
            I => \N__56955\
        );

    \I__13583\ : SRMux
    port map (
            O => \N__57573\,
            I => \N__56955\
        );

    \I__13582\ : SRMux
    port map (
            O => \N__57572\,
            I => \N__56955\
        );

    \I__13581\ : SRMux
    port map (
            O => \N__57571\,
            I => \N__56955\
        );

    \I__13580\ : SRMux
    port map (
            O => \N__57570\,
            I => \N__56955\
        );

    \I__13579\ : SRMux
    port map (
            O => \N__57569\,
            I => \N__56955\
        );

    \I__13578\ : SRMux
    port map (
            O => \N__57568\,
            I => \N__56955\
        );

    \I__13577\ : SRMux
    port map (
            O => \N__57567\,
            I => \N__56955\
        );

    \I__13576\ : SRMux
    port map (
            O => \N__57566\,
            I => \N__56955\
        );

    \I__13575\ : SRMux
    port map (
            O => \N__57565\,
            I => \N__56955\
        );

    \I__13574\ : SRMux
    port map (
            O => \N__57564\,
            I => \N__56955\
        );

    \I__13573\ : SRMux
    port map (
            O => \N__57563\,
            I => \N__56955\
        );

    \I__13572\ : SRMux
    port map (
            O => \N__57562\,
            I => \N__56955\
        );

    \I__13571\ : SRMux
    port map (
            O => \N__57561\,
            I => \N__56955\
        );

    \I__13570\ : SRMux
    port map (
            O => \N__57560\,
            I => \N__56955\
        );

    \I__13569\ : SRMux
    port map (
            O => \N__57559\,
            I => \N__56955\
        );

    \I__13568\ : SRMux
    port map (
            O => \N__57558\,
            I => \N__56955\
        );

    \I__13567\ : SRMux
    port map (
            O => \N__57557\,
            I => \N__56955\
        );

    \I__13566\ : SRMux
    port map (
            O => \N__57556\,
            I => \N__56955\
        );

    \I__13565\ : SRMux
    port map (
            O => \N__57555\,
            I => \N__56955\
        );

    \I__13564\ : SRMux
    port map (
            O => \N__57554\,
            I => \N__56955\
        );

    \I__13563\ : SRMux
    port map (
            O => \N__57553\,
            I => \N__56955\
        );

    \I__13562\ : SRMux
    port map (
            O => \N__57552\,
            I => \N__56955\
        );

    \I__13561\ : SRMux
    port map (
            O => \N__57551\,
            I => \N__56955\
        );

    \I__13560\ : SRMux
    port map (
            O => \N__57550\,
            I => \N__56955\
        );

    \I__13559\ : SRMux
    port map (
            O => \N__57549\,
            I => \N__56955\
        );

    \I__13558\ : SRMux
    port map (
            O => \N__57548\,
            I => \N__56955\
        );

    \I__13557\ : SRMux
    port map (
            O => \N__57547\,
            I => \N__56955\
        );

    \I__13556\ : SRMux
    port map (
            O => \N__57546\,
            I => \N__56955\
        );

    \I__13555\ : SRMux
    port map (
            O => \N__57545\,
            I => \N__56955\
        );

    \I__13554\ : SRMux
    port map (
            O => \N__57544\,
            I => \N__56955\
        );

    \I__13553\ : SRMux
    port map (
            O => \N__57543\,
            I => \N__56955\
        );

    \I__13552\ : SRMux
    port map (
            O => \N__57542\,
            I => \N__56955\
        );

    \I__13551\ : SRMux
    port map (
            O => \N__57541\,
            I => \N__56955\
        );

    \I__13550\ : SRMux
    port map (
            O => \N__57540\,
            I => \N__56955\
        );

    \I__13549\ : SRMux
    port map (
            O => \N__57539\,
            I => \N__56955\
        );

    \I__13548\ : SRMux
    port map (
            O => \N__57538\,
            I => \N__56955\
        );

    \I__13547\ : SRMux
    port map (
            O => \N__57537\,
            I => \N__56955\
        );

    \I__13546\ : SRMux
    port map (
            O => \N__57536\,
            I => \N__56955\
        );

    \I__13545\ : SRMux
    port map (
            O => \N__57535\,
            I => \N__56955\
        );

    \I__13544\ : SRMux
    port map (
            O => \N__57534\,
            I => \N__56955\
        );

    \I__13543\ : SRMux
    port map (
            O => \N__57533\,
            I => \N__56955\
        );

    \I__13542\ : SRMux
    port map (
            O => \N__57532\,
            I => \N__56955\
        );

    \I__13541\ : SRMux
    port map (
            O => \N__57531\,
            I => \N__56955\
        );

    \I__13540\ : SRMux
    port map (
            O => \N__57530\,
            I => \N__56955\
        );

    \I__13539\ : SRMux
    port map (
            O => \N__57529\,
            I => \N__56955\
        );

    \I__13538\ : SRMux
    port map (
            O => \N__57528\,
            I => \N__56955\
        );

    \I__13537\ : SRMux
    port map (
            O => \N__57527\,
            I => \N__56955\
        );

    \I__13536\ : SRMux
    port map (
            O => \N__57526\,
            I => \N__56955\
        );

    \I__13535\ : SRMux
    port map (
            O => \N__57525\,
            I => \N__56955\
        );

    \I__13534\ : SRMux
    port map (
            O => \N__57524\,
            I => \N__56955\
        );

    \I__13533\ : SRMux
    port map (
            O => \N__57523\,
            I => \N__56955\
        );

    \I__13532\ : SRMux
    port map (
            O => \N__57522\,
            I => \N__56955\
        );

    \I__13531\ : SRMux
    port map (
            O => \N__57521\,
            I => \N__56955\
        );

    \I__13530\ : SRMux
    port map (
            O => \N__57520\,
            I => \N__56955\
        );

    \I__13529\ : SRMux
    port map (
            O => \N__57519\,
            I => \N__56955\
        );

    \I__13528\ : SRMux
    port map (
            O => \N__57518\,
            I => \N__56955\
        );

    \I__13527\ : SRMux
    port map (
            O => \N__57517\,
            I => \N__56955\
        );

    \I__13526\ : SRMux
    port map (
            O => \N__57516\,
            I => \N__56955\
        );

    \I__13525\ : SRMux
    port map (
            O => \N__57515\,
            I => \N__56955\
        );

    \I__13524\ : SRMux
    port map (
            O => \N__57514\,
            I => \N__56955\
        );

    \I__13523\ : SRMux
    port map (
            O => \N__57513\,
            I => \N__56955\
        );

    \I__13522\ : SRMux
    port map (
            O => \N__57512\,
            I => \N__56955\
        );

    \I__13521\ : SRMux
    port map (
            O => \N__57511\,
            I => \N__56955\
        );

    \I__13520\ : SRMux
    port map (
            O => \N__57510\,
            I => \N__56955\
        );

    \I__13519\ : SRMux
    port map (
            O => \N__57509\,
            I => \N__56955\
        );

    \I__13518\ : SRMux
    port map (
            O => \N__57508\,
            I => \N__56955\
        );

    \I__13517\ : SRMux
    port map (
            O => \N__57507\,
            I => \N__56955\
        );

    \I__13516\ : SRMux
    port map (
            O => \N__57506\,
            I => \N__56955\
        );

    \I__13515\ : SRMux
    port map (
            O => \N__57505\,
            I => \N__56955\
        );

    \I__13514\ : SRMux
    port map (
            O => \N__57504\,
            I => \N__56955\
        );

    \I__13513\ : SRMux
    port map (
            O => \N__57503\,
            I => \N__56955\
        );

    \I__13512\ : SRMux
    port map (
            O => \N__57502\,
            I => \N__56955\
        );

    \I__13511\ : SRMux
    port map (
            O => \N__57501\,
            I => \N__56955\
        );

    \I__13510\ : SRMux
    port map (
            O => \N__57500\,
            I => \N__56955\
        );

    \I__13509\ : SRMux
    port map (
            O => \N__57499\,
            I => \N__56955\
        );

    \I__13508\ : SRMux
    port map (
            O => \N__57498\,
            I => \N__56955\
        );

    \I__13507\ : SRMux
    port map (
            O => \N__57497\,
            I => \N__56955\
        );

    \I__13506\ : SRMux
    port map (
            O => \N__57496\,
            I => \N__56955\
        );

    \I__13505\ : Glb2LocalMux
    port map (
            O => \N__57493\,
            I => \N__56955\
        );

    \I__13504\ : Glb2LocalMux
    port map (
            O => \N__57490\,
            I => \N__56955\
        );

    \I__13503\ : Glb2LocalMux
    port map (
            O => \N__57487\,
            I => \N__56955\
        );

    \I__13502\ : Glb2LocalMux
    port map (
            O => \N__57484\,
            I => \N__56955\
        );

    \I__13501\ : Glb2LocalMux
    port map (
            O => \N__57481\,
            I => \N__56955\
        );

    \I__13500\ : Glb2LocalMux
    port map (
            O => \N__57478\,
            I => \N__56955\
        );

    \I__13499\ : Glb2LocalMux
    port map (
            O => \N__57475\,
            I => \N__56955\
        );

    \I__13498\ : Glb2LocalMux
    port map (
            O => \N__57472\,
            I => \N__56955\
        );

    \I__13497\ : Glb2LocalMux
    port map (
            O => \N__57469\,
            I => \N__56955\
        );

    \I__13496\ : Glb2LocalMux
    port map (
            O => \N__57466\,
            I => \N__56955\
        );

    \I__13495\ : Glb2LocalMux
    port map (
            O => \N__57463\,
            I => \N__56955\
        );

    \I__13494\ : Glb2LocalMux
    port map (
            O => \N__57460\,
            I => \N__56955\
        );

    \I__13493\ : Glb2LocalMux
    port map (
            O => \N__57457\,
            I => \N__56955\
        );

    \I__13492\ : Glb2LocalMux
    port map (
            O => \N__57454\,
            I => \N__56955\
        );

    \I__13491\ : Glb2LocalMux
    port map (
            O => \N__57451\,
            I => \N__56955\
        );

    \I__13490\ : Glb2LocalMux
    port map (
            O => \N__57448\,
            I => \N__56955\
        );

    \I__13489\ : Glb2LocalMux
    port map (
            O => \N__57445\,
            I => \N__56955\
        );

    \I__13488\ : Glb2LocalMux
    port map (
            O => \N__57442\,
            I => \N__56955\
        );

    \I__13487\ : Glb2LocalMux
    port map (
            O => \N__57439\,
            I => \N__56955\
        );

    \I__13486\ : Glb2LocalMux
    port map (
            O => \N__57436\,
            I => \N__56955\
        );

    \I__13485\ : Glb2LocalMux
    port map (
            O => \N__57433\,
            I => \N__56955\
        );

    \I__13484\ : Glb2LocalMux
    port map (
            O => \N__57430\,
            I => \N__56955\
        );

    \I__13483\ : Glb2LocalMux
    port map (
            O => \N__57427\,
            I => \N__56955\
        );

    \I__13482\ : Glb2LocalMux
    port map (
            O => \N__57424\,
            I => \N__56955\
        );

    \I__13481\ : Glb2LocalMux
    port map (
            O => \N__57421\,
            I => \N__56955\
        );

    \I__13480\ : Glb2LocalMux
    port map (
            O => \N__57418\,
            I => \N__56955\
        );

    \I__13479\ : Glb2LocalMux
    port map (
            O => \N__57415\,
            I => \N__56955\
        );

    \I__13478\ : Glb2LocalMux
    port map (
            O => \N__57412\,
            I => \N__56955\
        );

    \I__13477\ : Glb2LocalMux
    port map (
            O => \N__57409\,
            I => \N__56955\
        );

    \I__13476\ : Glb2LocalMux
    port map (
            O => \N__57406\,
            I => \N__56955\
        );

    \I__13475\ : Glb2LocalMux
    port map (
            O => \N__57403\,
            I => \N__56955\
        );

    \I__13474\ : Glb2LocalMux
    port map (
            O => \N__57400\,
            I => \N__56955\
        );

    \I__13473\ : Glb2LocalMux
    port map (
            O => \N__57397\,
            I => \N__56955\
        );

    \I__13472\ : Glb2LocalMux
    port map (
            O => \N__57394\,
            I => \N__56955\
        );

    \I__13471\ : Glb2LocalMux
    port map (
            O => \N__57391\,
            I => \N__56955\
        );

    \I__13470\ : Glb2LocalMux
    port map (
            O => \N__57388\,
            I => \N__56955\
        );

    \I__13469\ : Glb2LocalMux
    port map (
            O => \N__57385\,
            I => \N__56955\
        );

    \I__13468\ : Glb2LocalMux
    port map (
            O => \N__57382\,
            I => \N__56955\
        );

    \I__13467\ : Glb2LocalMux
    port map (
            O => \N__57379\,
            I => \N__56955\
        );

    \I__13466\ : Glb2LocalMux
    port map (
            O => \N__57376\,
            I => \N__56955\
        );

    \I__13465\ : Glb2LocalMux
    port map (
            O => \N__57373\,
            I => \N__56955\
        );

    \I__13464\ : Glb2LocalMux
    port map (
            O => \N__57370\,
            I => \N__56955\
        );

    \I__13463\ : Glb2LocalMux
    port map (
            O => \N__57367\,
            I => \N__56955\
        );

    \I__13462\ : Glb2LocalMux
    port map (
            O => \N__57364\,
            I => \N__56955\
        );

    \I__13461\ : Glb2LocalMux
    port map (
            O => \N__57361\,
            I => \N__56955\
        );

    \I__13460\ : Glb2LocalMux
    port map (
            O => \N__57358\,
            I => \N__56955\
        );

    \I__13459\ : GlobalMux
    port map (
            O => \N__56955\,
            I => \N__56952\
        );

    \I__13458\ : gio2CtrlBuf
    port map (
            O => \N__56952\,
            I => reset_system_g
        );

    \I__13457\ : InMux
    port map (
            O => \N__56949\,
            I => \N__56946\
        );

    \I__13456\ : LocalMux
    port map (
            O => \N__56946\,
            I => \N__56943\
        );

    \I__13455\ : Odrv4
    port map (
            O => \N__56943\,
            I => \pid_front.O_4\
        );

    \I__13454\ : CascadeMux
    port map (
            O => \N__56940\,
            I => \N__56936\
        );

    \I__13453\ : CascadeMux
    port map (
            O => \N__56939\,
            I => \N__56932\
        );

    \I__13452\ : InMux
    port map (
            O => \N__56936\,
            I => \N__56929\
        );

    \I__13451\ : InMux
    port map (
            O => \N__56935\,
            I => \N__56926\
        );

    \I__13450\ : InMux
    port map (
            O => \N__56932\,
            I => \N__56923\
        );

    \I__13449\ : LocalMux
    port map (
            O => \N__56929\,
            I => \N__56920\
        );

    \I__13448\ : LocalMux
    port map (
            O => \N__56926\,
            I => \N__56915\
        );

    \I__13447\ : LocalMux
    port map (
            O => \N__56923\,
            I => \N__56915\
        );

    \I__13446\ : Span4Mux_v
    port map (
            O => \N__56920\,
            I => \N__56912\
        );

    \I__13445\ : Sp12to4
    port map (
            O => \N__56915\,
            I => \N__56909\
        );

    \I__13444\ : Sp12to4
    port map (
            O => \N__56912\,
            I => \N__56904\
        );

    \I__13443\ : Span12Mux_h
    port map (
            O => \N__56909\,
            I => \N__56904\
        );

    \I__13442\ : Odrv12
    port map (
            O => \N__56904\,
            I => \pid_front.error_d_regZ0Z_0\
        );

    \I__13441\ : InMux
    port map (
            O => \N__56901\,
            I => \N__56898\
        );

    \I__13440\ : LocalMux
    port map (
            O => \N__56898\,
            I => \pid_front.O_5\
        );

    \I__13439\ : InMux
    port map (
            O => \N__56895\,
            I => \N__56890\
        );

    \I__13438\ : InMux
    port map (
            O => \N__56894\,
            I => \N__56887\
        );

    \I__13437\ : CascadeMux
    port map (
            O => \N__56893\,
            I => \N__56884\
        );

    \I__13436\ : LocalMux
    port map (
            O => \N__56890\,
            I => \N__56881\
        );

    \I__13435\ : LocalMux
    port map (
            O => \N__56887\,
            I => \N__56878\
        );

    \I__13434\ : InMux
    port map (
            O => \N__56884\,
            I => \N__56875\
        );

    \I__13433\ : Span4Mux_v
    port map (
            O => \N__56881\,
            I => \N__56868\
        );

    \I__13432\ : Span4Mux_v
    port map (
            O => \N__56878\,
            I => \N__56868\
        );

    \I__13431\ : LocalMux
    port map (
            O => \N__56875\,
            I => \N__56868\
        );

    \I__13430\ : Sp12to4
    port map (
            O => \N__56868\,
            I => \N__56865\
        );

    \I__13429\ : Span12Mux_h
    port map (
            O => \N__56865\,
            I => \N__56862\
        );

    \I__13428\ : Odrv12
    port map (
            O => \N__56862\,
            I => \pid_front.error_d_regZ0Z_1\
        );

    \I__13427\ : InMux
    port map (
            O => \N__56859\,
            I => \N__56856\
        );

    \I__13426\ : LocalMux
    port map (
            O => \N__56856\,
            I => \N__56853\
        );

    \I__13425\ : Odrv4
    port map (
            O => \N__56853\,
            I => \pid_front.O_17\
        );

    \I__13424\ : InMux
    port map (
            O => \N__56850\,
            I => \N__56841\
        );

    \I__13423\ : InMux
    port map (
            O => \N__56849\,
            I => \N__56841\
        );

    \I__13422\ : InMux
    port map (
            O => \N__56848\,
            I => \N__56841\
        );

    \I__13421\ : LocalMux
    port map (
            O => \N__56841\,
            I => \N__56838\
        );

    \I__13420\ : Span12Mux_h
    port map (
            O => \N__56838\,
            I => \N__56835\
        );

    \I__13419\ : Odrv12
    port map (
            O => \N__56835\,
            I => \pid_front.error_d_regZ0Z_13\
        );

    \I__13418\ : InMux
    port map (
            O => \N__56832\,
            I => \N__56829\
        );

    \I__13417\ : LocalMux
    port map (
            O => \N__56829\,
            I => \N__56826\
        );

    \I__13416\ : Odrv4
    port map (
            O => \N__56826\,
            I => \pid_front.O_15\
        );

    \I__13415\ : InMux
    port map (
            O => \N__56823\,
            I => \N__56819\
        );

    \I__13414\ : InMux
    port map (
            O => \N__56822\,
            I => \N__56816\
        );

    \I__13413\ : LocalMux
    port map (
            O => \N__56819\,
            I => \N__56812\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__56816\,
            I => \N__56809\
        );

    \I__13411\ : InMux
    port map (
            O => \N__56815\,
            I => \N__56806\
        );

    \I__13410\ : Span4Mux_v
    port map (
            O => \N__56812\,
            I => \N__56803\
        );

    \I__13409\ : Span4Mux_v
    port map (
            O => \N__56809\,
            I => \N__56800\
        );

    \I__13408\ : LocalMux
    port map (
            O => \N__56806\,
            I => \N__56797\
        );

    \I__13407\ : Span4Mux_h
    port map (
            O => \N__56803\,
            I => \N__56794\
        );

    \I__13406\ : Sp12to4
    port map (
            O => \N__56800\,
            I => \N__56787\
        );

    \I__13405\ : Span12Mux_h
    port map (
            O => \N__56797\,
            I => \N__56787\
        );

    \I__13404\ : Sp12to4
    port map (
            O => \N__56794\,
            I => \N__56787\
        );

    \I__13403\ : Odrv12
    port map (
            O => \N__56787\,
            I => \pid_front.error_d_regZ0Z_11\
        );

    \I__13402\ : InMux
    port map (
            O => \N__56784\,
            I => \N__56781\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__56781\,
            I => \N__56778\
        );

    \I__13400\ : Odrv4
    port map (
            O => \N__56778\,
            I => \pid_front.O_13\
        );

    \I__13399\ : CascadeMux
    port map (
            O => \N__56775\,
            I => \N__56770\
        );

    \I__13398\ : InMux
    port map (
            O => \N__56774\,
            I => \N__56765\
        );

    \I__13397\ : InMux
    port map (
            O => \N__56773\,
            I => \N__56765\
        );

    \I__13396\ : InMux
    port map (
            O => \N__56770\,
            I => \N__56762\
        );

    \I__13395\ : LocalMux
    port map (
            O => \N__56765\,
            I => \N__56759\
        );

    \I__13394\ : LocalMux
    port map (
            O => \N__56762\,
            I => \N__56756\
        );

    \I__13393\ : Span4Mux_v
    port map (
            O => \N__56759\,
            I => \N__56753\
        );

    \I__13392\ : Span12Mux_h
    port map (
            O => \N__56756\,
            I => \N__56750\
        );

    \I__13391\ : Span4Mux_h
    port map (
            O => \N__56753\,
            I => \N__56747\
        );

    \I__13390\ : Span12Mux_h
    port map (
            O => \N__56750\,
            I => \N__56744\
        );

    \I__13389\ : Sp12to4
    port map (
            O => \N__56747\,
            I => \N__56741\
        );

    \I__13388\ : Odrv12
    port map (
            O => \N__56744\,
            I => \pid_front.error_d_regZ0Z_9\
        );

    \I__13387\ : Odrv12
    port map (
            O => \N__56741\,
            I => \pid_front.error_d_regZ0Z_9\
        );

    \I__13386\ : InMux
    port map (
            O => \N__56736\,
            I => \N__56733\
        );

    \I__13385\ : LocalMux
    port map (
            O => \N__56733\,
            I => \N__56730\
        );

    \I__13384\ : Odrv4
    port map (
            O => \N__56730\,
            I => \pid_front.O_20\
        );

    \I__13383\ : InMux
    port map (
            O => \N__56727\,
            I => \N__56724\
        );

    \I__13382\ : LocalMux
    port map (
            O => \N__56724\,
            I => \N__56720\
        );

    \I__13381\ : InMux
    port map (
            O => \N__56723\,
            I => \N__56717\
        );

    \I__13380\ : Span4Mux_h
    port map (
            O => \N__56720\,
            I => \N__56714\
        );

    \I__13379\ : LocalMux
    port map (
            O => \N__56717\,
            I => \N__56711\
        );

    \I__13378\ : Span4Mux_v
    port map (
            O => \N__56714\,
            I => \N__56705\
        );

    \I__13377\ : Span4Mux_h
    port map (
            O => \N__56711\,
            I => \N__56705\
        );

    \I__13376\ : InMux
    port map (
            O => \N__56710\,
            I => \N__56702\
        );

    \I__13375\ : Span4Mux_h
    port map (
            O => \N__56705\,
            I => \N__56699\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__56702\,
            I => \N__56696\
        );

    \I__13373\ : Span4Mux_h
    port map (
            O => \N__56699\,
            I => \N__56693\
        );

    \I__13372\ : Span12Mux_h
    port map (
            O => \N__56696\,
            I => \N__56690\
        );

    \I__13371\ : Span4Mux_h
    port map (
            O => \N__56693\,
            I => \N__56687\
        );

    \I__13370\ : Odrv12
    port map (
            O => \N__56690\,
            I => \pid_front.error_d_regZ0Z_16\
        );

    \I__13369\ : Odrv4
    port map (
            O => \N__56687\,
            I => \pid_front.error_d_regZ0Z_16\
        );

    \I__13368\ : InMux
    port map (
            O => \N__56682\,
            I => \N__56679\
        );

    \I__13367\ : LocalMux
    port map (
            O => \N__56679\,
            I => \N__56676\
        );

    \I__13366\ : Odrv4
    port map (
            O => \N__56676\,
            I => \pid_front.O_21\
        );

    \I__13365\ : InMux
    port map (
            O => \N__56673\,
            I => \N__56664\
        );

    \I__13364\ : InMux
    port map (
            O => \N__56672\,
            I => \N__56664\
        );

    \I__13363\ : InMux
    port map (
            O => \N__56671\,
            I => \N__56664\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__56664\,
            I => \N__56661\
        );

    \I__13361\ : Span4Mux_h
    port map (
            O => \N__56661\,
            I => \N__56658\
        );

    \I__13360\ : Span4Mux_h
    port map (
            O => \N__56658\,
            I => \N__56655\
        );

    \I__13359\ : Span4Mux_h
    port map (
            O => \N__56655\,
            I => \N__56652\
        );

    \I__13358\ : Odrv4
    port map (
            O => \N__56652\,
            I => \pid_front.error_d_regZ0Z_17\
        );

    \I__13357\ : InMux
    port map (
            O => \N__56649\,
            I => \N__56640\
        );

    \I__13356\ : InMux
    port map (
            O => \N__56648\,
            I => \N__56640\
        );

    \I__13355\ : InMux
    port map (
            O => \N__56647\,
            I => \N__56640\
        );

    \I__13354\ : LocalMux
    port map (
            O => \N__56640\,
            I => \N__56637\
        );

    \I__13353\ : Odrv12
    port map (
            O => \N__56637\,
            I => \pid_side.error_d_regZ0Z_7\
        );

    \I__13352\ : InMux
    port map (
            O => \N__56634\,
            I => \N__56631\
        );

    \I__13351\ : LocalMux
    port map (
            O => \N__56631\,
            I => \pid_side.O_1_20\
        );

    \I__13350\ : InMux
    port map (
            O => \N__56628\,
            I => \N__56619\
        );

    \I__13349\ : InMux
    port map (
            O => \N__56627\,
            I => \N__56619\
        );

    \I__13348\ : InMux
    port map (
            O => \N__56626\,
            I => \N__56619\
        );

    \I__13347\ : LocalMux
    port map (
            O => \N__56619\,
            I => \N__56616\
        );

    \I__13346\ : Span4Mux_v
    port map (
            O => \N__56616\,
            I => \N__56613\
        );

    \I__13345\ : Odrv4
    port map (
            O => \N__56613\,
            I => \pid_side.error_d_regZ0Z_16\
        );

    \I__13344\ : CEMux
    port map (
            O => \N__56610\,
            I => \N__56604\
        );

    \I__13343\ : CEMux
    port map (
            O => \N__56609\,
            I => \N__56600\
        );

    \I__13342\ : CEMux
    port map (
            O => \N__56608\,
            I => \N__56594\
        );

    \I__13341\ : CEMux
    port map (
            O => \N__56607\,
            I => \N__56589\
        );

    \I__13340\ : LocalMux
    port map (
            O => \N__56604\,
            I => \N__56586\
        );

    \I__13339\ : CEMux
    port map (
            O => \N__56603\,
            I => \N__56583\
        );

    \I__13338\ : LocalMux
    port map (
            O => \N__56600\,
            I => \N__56580\
        );

    \I__13337\ : CEMux
    port map (
            O => \N__56599\,
            I => \N__56577\
        );

    \I__13336\ : CEMux
    port map (
            O => \N__56598\,
            I => \N__56574\
        );

    \I__13335\ : CEMux
    port map (
            O => \N__56597\,
            I => \N__56571\
        );

    \I__13334\ : LocalMux
    port map (
            O => \N__56594\,
            I => \N__56568\
        );

    \I__13333\ : CEMux
    port map (
            O => \N__56593\,
            I => \N__56565\
        );

    \I__13332\ : CEMux
    port map (
            O => \N__56592\,
            I => \N__56561\
        );

    \I__13331\ : LocalMux
    port map (
            O => \N__56589\,
            I => \N__56558\
        );

    \I__13330\ : Span4Mux_v
    port map (
            O => \N__56586\,
            I => \N__56553\
        );

    \I__13329\ : LocalMux
    port map (
            O => \N__56583\,
            I => \N__56553\
        );

    \I__13328\ : Span4Mux_v
    port map (
            O => \N__56580\,
            I => \N__56544\
        );

    \I__13327\ : LocalMux
    port map (
            O => \N__56577\,
            I => \N__56544\
        );

    \I__13326\ : LocalMux
    port map (
            O => \N__56574\,
            I => \N__56544\
        );

    \I__13325\ : LocalMux
    port map (
            O => \N__56571\,
            I => \N__56544\
        );

    \I__13324\ : Span4Mux_v
    port map (
            O => \N__56568\,
            I => \N__56541\
        );

    \I__13323\ : LocalMux
    port map (
            O => \N__56565\,
            I => \N__56538\
        );

    \I__13322\ : CEMux
    port map (
            O => \N__56564\,
            I => \N__56535\
        );

    \I__13321\ : LocalMux
    port map (
            O => \N__56561\,
            I => \N__56532\
        );

    \I__13320\ : Span4Mux_v
    port map (
            O => \N__56558\,
            I => \N__56529\
        );

    \I__13319\ : Span4Mux_v
    port map (
            O => \N__56553\,
            I => \N__56522\
        );

    \I__13318\ : Span4Mux_v
    port map (
            O => \N__56544\,
            I => \N__56522\
        );

    \I__13317\ : Span4Mux_s1_h
    port map (
            O => \N__56541\,
            I => \N__56522\
        );

    \I__13316\ : Span4Mux_v
    port map (
            O => \N__56538\,
            I => \N__56515\
        );

    \I__13315\ : LocalMux
    port map (
            O => \N__56535\,
            I => \N__56515\
        );

    \I__13314\ : Span4Mux_v
    port map (
            O => \N__56532\,
            I => \N__56515\
        );

    \I__13313\ : Odrv4
    port map (
            O => \N__56529\,
            I => \pid_side.N_599_0\
        );

    \I__13312\ : Odrv4
    port map (
            O => \N__56522\,
            I => \pid_side.N_599_0\
        );

    \I__13311\ : Odrv4
    port map (
            O => \N__56515\,
            I => \pid_side.N_599_0\
        );

    \I__13310\ : InMux
    port map (
            O => \N__56508\,
            I => \N__56503\
        );

    \I__13309\ : InMux
    port map (
            O => \N__56507\,
            I => \N__56500\
        );

    \I__13308\ : InMux
    port map (
            O => \N__56506\,
            I => \N__56497\
        );

    \I__13307\ : LocalMux
    port map (
            O => \N__56503\,
            I => \N__56494\
        );

    \I__13306\ : LocalMux
    port map (
            O => \N__56500\,
            I => \N__56491\
        );

    \I__13305\ : LocalMux
    port map (
            O => \N__56497\,
            I => \N__56488\
        );

    \I__13304\ : Span4Mux_s3_h
    port map (
            O => \N__56494\,
            I => \N__56483\
        );

    \I__13303\ : Span4Mux_v
    port map (
            O => \N__56491\,
            I => \N__56480\
        );

    \I__13302\ : Span4Mux_v
    port map (
            O => \N__56488\,
            I => \N__56476\
        );

    \I__13301\ : InMux
    port map (
            O => \N__56487\,
            I => \N__56473\
        );

    \I__13300\ : InMux
    port map (
            O => \N__56486\,
            I => \N__56470\
        );

    \I__13299\ : Span4Mux_h
    port map (
            O => \N__56483\,
            I => \N__56467\
        );

    \I__13298\ : Span4Mux_h
    port map (
            O => \N__56480\,
            I => \N__56461\
        );

    \I__13297\ : InMux
    port map (
            O => \N__56479\,
            I => \N__56458\
        );

    \I__13296\ : Span4Mux_h
    port map (
            O => \N__56476\,
            I => \N__56455\
        );

    \I__13295\ : LocalMux
    port map (
            O => \N__56473\,
            I => \N__56451\
        );

    \I__13294\ : LocalMux
    port map (
            O => \N__56470\,
            I => \N__56448\
        );

    \I__13293\ : Span4Mux_h
    port map (
            O => \N__56467\,
            I => \N__56445\
        );

    \I__13292\ : InMux
    port map (
            O => \N__56466\,
            I => \N__56442\
        );

    \I__13291\ : InMux
    port map (
            O => \N__56465\,
            I => \N__56437\
        );

    \I__13290\ : InMux
    port map (
            O => \N__56464\,
            I => \N__56434\
        );

    \I__13289\ : Span4Mux_v
    port map (
            O => \N__56461\,
            I => \N__56428\
        );

    \I__13288\ : LocalMux
    port map (
            O => \N__56458\,
            I => \N__56428\
        );

    \I__13287\ : Span4Mux_v
    port map (
            O => \N__56455\,
            I => \N__56425\
        );

    \I__13286\ : InMux
    port map (
            O => \N__56454\,
            I => \N__56422\
        );

    \I__13285\ : Span4Mux_v
    port map (
            O => \N__56451\,
            I => \N__56417\
        );

    \I__13284\ : Span4Mux_s3_h
    port map (
            O => \N__56448\,
            I => \N__56417\
        );

    \I__13283\ : Span4Mux_h
    port map (
            O => \N__56445\,
            I => \N__56412\
        );

    \I__13282\ : LocalMux
    port map (
            O => \N__56442\,
            I => \N__56412\
        );

    \I__13281\ : CascadeMux
    port map (
            O => \N__56441\,
            I => \N__56409\
        );

    \I__13280\ : InMux
    port map (
            O => \N__56440\,
            I => \N__56406\
        );

    \I__13279\ : LocalMux
    port map (
            O => \N__56437\,
            I => \N__56403\
        );

    \I__13278\ : LocalMux
    port map (
            O => \N__56434\,
            I => \N__56400\
        );

    \I__13277\ : InMux
    port map (
            O => \N__56433\,
            I => \N__56397\
        );

    \I__13276\ : Span4Mux_h
    port map (
            O => \N__56428\,
            I => \N__56394\
        );

    \I__13275\ : Span4Mux_v
    port map (
            O => \N__56425\,
            I => \N__56389\
        );

    \I__13274\ : LocalMux
    port map (
            O => \N__56422\,
            I => \N__56389\
        );

    \I__13273\ : Span4Mux_h
    port map (
            O => \N__56417\,
            I => \N__56385\
        );

    \I__13272\ : Span4Mux_v
    port map (
            O => \N__56412\,
            I => \N__56381\
        );

    \I__13271\ : InMux
    port map (
            O => \N__56409\,
            I => \N__56378\
        );

    \I__13270\ : LocalMux
    port map (
            O => \N__56406\,
            I => \N__56375\
        );

    \I__13269\ : Span4Mux_v
    port map (
            O => \N__56403\,
            I => \N__56368\
        );

    \I__13268\ : Span4Mux_v
    port map (
            O => \N__56400\,
            I => \N__56368\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__56397\,
            I => \N__56368\
        );

    \I__13266\ : Span4Mux_h
    port map (
            O => \N__56394\,
            I => \N__56363\
        );

    \I__13265\ : Span4Mux_v
    port map (
            O => \N__56389\,
            I => \N__56363\
        );

    \I__13264\ : InMux
    port map (
            O => \N__56388\,
            I => \N__56360\
        );

    \I__13263\ : Sp12to4
    port map (
            O => \N__56385\,
            I => \N__56357\
        );

    \I__13262\ : InMux
    port map (
            O => \N__56384\,
            I => \N__56354\
        );

    \I__13261\ : Span4Mux_v
    port map (
            O => \N__56381\,
            I => \N__56345\
        );

    \I__13260\ : LocalMux
    port map (
            O => \N__56378\,
            I => \N__56345\
        );

    \I__13259\ : Span4Mux_v
    port map (
            O => \N__56375\,
            I => \N__56345\
        );

    \I__13258\ : Span4Mux_h
    port map (
            O => \N__56368\,
            I => \N__56345\
        );

    \I__13257\ : Odrv4
    port map (
            O => \N__56363\,
            I => uart_pc_data_0
        );

    \I__13256\ : LocalMux
    port map (
            O => \N__56360\,
            I => uart_pc_data_0
        );

    \I__13255\ : Odrv12
    port map (
            O => \N__56357\,
            I => uart_pc_data_0
        );

    \I__13254\ : LocalMux
    port map (
            O => \N__56354\,
            I => uart_pc_data_0
        );

    \I__13253\ : Odrv4
    port map (
            O => \N__56345\,
            I => uart_pc_data_0
        );

    \I__13252\ : InMux
    port map (
            O => \N__56334\,
            I => \N__56331\
        );

    \I__13251\ : LocalMux
    port map (
            O => \N__56331\,
            I => \N__56328\
        );

    \I__13250\ : Span4Mux_v
    port map (
            O => \N__56328\,
            I => \N__56325\
        );

    \I__13249\ : Span4Mux_v
    port map (
            O => \N__56325\,
            I => \N__56321\
        );

    \I__13248\ : InMux
    port map (
            O => \N__56324\,
            I => \N__56318\
        );

    \I__13247\ : Odrv4
    port map (
            O => \N__56321\,
            I => xy_kd_0
        );

    \I__13246\ : LocalMux
    port map (
            O => \N__56318\,
            I => xy_kd_0
        );

    \I__13245\ : InMux
    port map (
            O => \N__56313\,
            I => \N__56308\
        );

    \I__13244\ : InMux
    port map (
            O => \N__56312\,
            I => \N__56305\
        );

    \I__13243\ : InMux
    port map (
            O => \N__56311\,
            I => \N__56301\
        );

    \I__13242\ : LocalMux
    port map (
            O => \N__56308\,
            I => \N__56298\
        );

    \I__13241\ : LocalMux
    port map (
            O => \N__56305\,
            I => \N__56295\
        );

    \I__13240\ : InMux
    port map (
            O => \N__56304\,
            I => \N__56292\
        );

    \I__13239\ : LocalMux
    port map (
            O => \N__56301\,
            I => \N__56289\
        );

    \I__13238\ : Span4Mux_h
    port map (
            O => \N__56298\,
            I => \N__56286\
        );

    \I__13237\ : Span4Mux_h
    port map (
            O => \N__56295\,
            I => \N__56279\
        );

    \I__13236\ : LocalMux
    port map (
            O => \N__56292\,
            I => \N__56279\
        );

    \I__13235\ : Span4Mux_v
    port map (
            O => \N__56289\,
            I => \N__56275\
        );

    \I__13234\ : Span4Mux_h
    port map (
            O => \N__56286\,
            I => \N__56272\
        );

    \I__13233\ : InMux
    port map (
            O => \N__56285\,
            I => \N__56267\
        );

    \I__13232\ : InMux
    port map (
            O => \N__56284\,
            I => \N__56263\
        );

    \I__13231\ : Span4Mux_v
    port map (
            O => \N__56279\,
            I => \N__56260\
        );

    \I__13230\ : InMux
    port map (
            O => \N__56278\,
            I => \N__56257\
        );

    \I__13229\ : Span4Mux_v
    port map (
            O => \N__56275\,
            I => \N__56252\
        );

    \I__13228\ : Span4Mux_h
    port map (
            O => \N__56272\,
            I => \N__56252\
        );

    \I__13227\ : InMux
    port map (
            O => \N__56271\,
            I => \N__56249\
        );

    \I__13226\ : InMux
    port map (
            O => \N__56270\,
            I => \N__56246\
        );

    \I__13225\ : LocalMux
    port map (
            O => \N__56267\,
            I => \N__56243\
        );

    \I__13224\ : InMux
    port map (
            O => \N__56266\,
            I => \N__56239\
        );

    \I__13223\ : LocalMux
    port map (
            O => \N__56263\,
            I => \N__56236\
        );

    \I__13222\ : Span4Mux_v
    port map (
            O => \N__56260\,
            I => \N__56233\
        );

    \I__13221\ : LocalMux
    port map (
            O => \N__56257\,
            I => \N__56230\
        );

    \I__13220\ : Span4Mux_h
    port map (
            O => \N__56252\,
            I => \N__56225\
        );

    \I__13219\ : LocalMux
    port map (
            O => \N__56249\,
            I => \N__56225\
        );

    \I__13218\ : LocalMux
    port map (
            O => \N__56246\,
            I => \N__56221\
        );

    \I__13217\ : Span12Mux_v
    port map (
            O => \N__56243\,
            I => \N__56217\
        );

    \I__13216\ : InMux
    port map (
            O => \N__56242\,
            I => \N__56214\
        );

    \I__13215\ : LocalMux
    port map (
            O => \N__56239\,
            I => \N__56211\
        );

    \I__13214\ : Span4Mux_v
    port map (
            O => \N__56236\,
            I => \N__56208\
        );

    \I__13213\ : Span4Mux_v
    port map (
            O => \N__56233\,
            I => \N__56203\
        );

    \I__13212\ : Span4Mux_v
    port map (
            O => \N__56230\,
            I => \N__56203\
        );

    \I__13211\ : Span4Mux_v
    port map (
            O => \N__56225\,
            I => \N__56200\
        );

    \I__13210\ : InMux
    port map (
            O => \N__56224\,
            I => \N__56197\
        );

    \I__13209\ : Span4Mux_h
    port map (
            O => \N__56221\,
            I => \N__56194\
        );

    \I__13208\ : InMux
    port map (
            O => \N__56220\,
            I => \N__56191\
        );

    \I__13207\ : Span12Mux_h
    port map (
            O => \N__56217\,
            I => \N__56186\
        );

    \I__13206\ : LocalMux
    port map (
            O => \N__56214\,
            I => \N__56186\
        );

    \I__13205\ : Span4Mux_h
    port map (
            O => \N__56211\,
            I => \N__56183\
        );

    \I__13204\ : Span4Mux_h
    port map (
            O => \N__56208\,
            I => \N__56174\
        );

    \I__13203\ : Span4Mux_h
    port map (
            O => \N__56203\,
            I => \N__56174\
        );

    \I__13202\ : Span4Mux_v
    port map (
            O => \N__56200\,
            I => \N__56174\
        );

    \I__13201\ : LocalMux
    port map (
            O => \N__56197\,
            I => \N__56174\
        );

    \I__13200\ : Odrv4
    port map (
            O => \N__56194\,
            I => uart_pc_data_1
        );

    \I__13199\ : LocalMux
    port map (
            O => \N__56191\,
            I => uart_pc_data_1
        );

    \I__13198\ : Odrv12
    port map (
            O => \N__56186\,
            I => uart_pc_data_1
        );

    \I__13197\ : Odrv4
    port map (
            O => \N__56183\,
            I => uart_pc_data_1
        );

    \I__13196\ : Odrv4
    port map (
            O => \N__56174\,
            I => uart_pc_data_1
        );

    \I__13195\ : InMux
    port map (
            O => \N__56163\,
            I => \N__56160\
        );

    \I__13194\ : LocalMux
    port map (
            O => \N__56160\,
            I => \N__56157\
        );

    \I__13193\ : Span4Mux_v
    port map (
            O => \N__56157\,
            I => \N__56154\
        );

    \I__13192\ : Span4Mux_v
    port map (
            O => \N__56154\,
            I => \N__56150\
        );

    \I__13191\ : InMux
    port map (
            O => \N__56153\,
            I => \N__56147\
        );

    \I__13190\ : Odrv4
    port map (
            O => \N__56150\,
            I => xy_kd_1
        );

    \I__13189\ : LocalMux
    port map (
            O => \N__56147\,
            I => xy_kd_1
        );

    \I__13188\ : InMux
    port map (
            O => \N__56142\,
            I => \N__56136\
        );

    \I__13187\ : InMux
    port map (
            O => \N__56141\,
            I => \N__56133\
        );

    \I__13186\ : InMux
    port map (
            O => \N__56140\,
            I => \N__56129\
        );

    \I__13185\ : InMux
    port map (
            O => \N__56139\,
            I => \N__56126\
        );

    \I__13184\ : LocalMux
    port map (
            O => \N__56136\,
            I => \N__56121\
        );

    \I__13183\ : LocalMux
    port map (
            O => \N__56133\,
            I => \N__56118\
        );

    \I__13182\ : InMux
    port map (
            O => \N__56132\,
            I => \N__56115\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__56129\,
            I => \N__56112\
        );

    \I__13180\ : LocalMux
    port map (
            O => \N__56126\,
            I => \N__56107\
        );

    \I__13179\ : InMux
    port map (
            O => \N__56125\,
            I => \N__56102\
        );

    \I__13178\ : InMux
    port map (
            O => \N__56124\,
            I => \N__56099\
        );

    \I__13177\ : Span4Mux_v
    port map (
            O => \N__56121\,
            I => \N__56096\
        );

    \I__13176\ : Span4Mux_v
    port map (
            O => \N__56118\,
            I => \N__56093\
        );

    \I__13175\ : LocalMux
    port map (
            O => \N__56115\,
            I => \N__56090\
        );

    \I__13174\ : Span4Mux_v
    port map (
            O => \N__56112\,
            I => \N__56087\
        );

    \I__13173\ : InMux
    port map (
            O => \N__56111\,
            I => \N__56084\
        );

    \I__13172\ : InMux
    port map (
            O => \N__56110\,
            I => \N__56081\
        );

    \I__13171\ : Span4Mux_v
    port map (
            O => \N__56107\,
            I => \N__56078\
        );

    \I__13170\ : CascadeMux
    port map (
            O => \N__56106\,
            I => \N__56075\
        );

    \I__13169\ : InMux
    port map (
            O => \N__56105\,
            I => \N__56070\
        );

    \I__13168\ : LocalMux
    port map (
            O => \N__56102\,
            I => \N__56067\
        );

    \I__13167\ : LocalMux
    port map (
            O => \N__56099\,
            I => \N__56064\
        );

    \I__13166\ : Sp12to4
    port map (
            O => \N__56096\,
            I => \N__56061\
        );

    \I__13165\ : Sp12to4
    port map (
            O => \N__56093\,
            I => \N__56058\
        );

    \I__13164\ : Span4Mux_v
    port map (
            O => \N__56090\,
            I => \N__56053\
        );

    \I__13163\ : Span4Mux_h
    port map (
            O => \N__56087\,
            I => \N__56053\
        );

    \I__13162\ : LocalMux
    port map (
            O => \N__56084\,
            I => \N__56050\
        );

    \I__13161\ : LocalMux
    port map (
            O => \N__56081\,
            I => \N__56047\
        );

    \I__13160\ : Span4Mux_h
    port map (
            O => \N__56078\,
            I => \N__56043\
        );

    \I__13159\ : InMux
    port map (
            O => \N__56075\,
            I => \N__56040\
        );

    \I__13158\ : InMux
    port map (
            O => \N__56074\,
            I => \N__56037\
        );

    \I__13157\ : CascadeMux
    port map (
            O => \N__56073\,
            I => \N__56034\
        );

    \I__13156\ : LocalMux
    port map (
            O => \N__56070\,
            I => \N__56031\
        );

    \I__13155\ : Span4Mux_v
    port map (
            O => \N__56067\,
            I => \N__56028\
        );

    \I__13154\ : Span4Mux_v
    port map (
            O => \N__56064\,
            I => \N__56025\
        );

    \I__13153\ : Span12Mux_h
    port map (
            O => \N__56061\,
            I => \N__56020\
        );

    \I__13152\ : Span12Mux_s6_h
    port map (
            O => \N__56058\,
            I => \N__56020\
        );

    \I__13151\ : Span4Mux_v
    port map (
            O => \N__56053\,
            I => \N__56017\
        );

    \I__13150\ : Span4Mux_v
    port map (
            O => \N__56050\,
            I => \N__56013\
        );

    \I__13149\ : Span4Mux_v
    port map (
            O => \N__56047\,
            I => \N__56010\
        );

    \I__13148\ : InMux
    port map (
            O => \N__56046\,
            I => \N__56007\
        );

    \I__13147\ : Span4Mux_v
    port map (
            O => \N__56043\,
            I => \N__56002\
        );

    \I__13146\ : LocalMux
    port map (
            O => \N__56040\,
            I => \N__56002\
        );

    \I__13145\ : LocalMux
    port map (
            O => \N__56037\,
            I => \N__55998\
        );

    \I__13144\ : InMux
    port map (
            O => \N__56034\,
            I => \N__55995\
        );

    \I__13143\ : Span4Mux_v
    port map (
            O => \N__56031\,
            I => \N__55990\
        );

    \I__13142\ : Span4Mux_h
    port map (
            O => \N__56028\,
            I => \N__55990\
        );

    \I__13141\ : Sp12to4
    port map (
            O => \N__56025\,
            I => \N__55983\
        );

    \I__13140\ : Span12Mux_v
    port map (
            O => \N__56020\,
            I => \N__55983\
        );

    \I__13139\ : Sp12to4
    port map (
            O => \N__56017\,
            I => \N__55983\
        );

    \I__13138\ : InMux
    port map (
            O => \N__56016\,
            I => \N__55980\
        );

    \I__13137\ : Span4Mux_h
    port map (
            O => \N__56013\,
            I => \N__55971\
        );

    \I__13136\ : Span4Mux_v
    port map (
            O => \N__56010\,
            I => \N__55971\
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__56007\,
            I => \N__55971\
        );

    \I__13134\ : Span4Mux_v
    port map (
            O => \N__56002\,
            I => \N__55971\
        );

    \I__13133\ : InMux
    port map (
            O => \N__56001\,
            I => \N__55968\
        );

    \I__13132\ : Span4Mux_v
    port map (
            O => \N__55998\,
            I => \N__55965\
        );

    \I__13131\ : LocalMux
    port map (
            O => \N__55995\,
            I => uart_pc_data_2
        );

    \I__13130\ : Odrv4
    port map (
            O => \N__55990\,
            I => uart_pc_data_2
        );

    \I__13129\ : Odrv12
    port map (
            O => \N__55983\,
            I => uart_pc_data_2
        );

    \I__13128\ : LocalMux
    port map (
            O => \N__55980\,
            I => uart_pc_data_2
        );

    \I__13127\ : Odrv4
    port map (
            O => \N__55971\,
            I => uart_pc_data_2
        );

    \I__13126\ : LocalMux
    port map (
            O => \N__55968\,
            I => uart_pc_data_2
        );

    \I__13125\ : Odrv4
    port map (
            O => \N__55965\,
            I => uart_pc_data_2
        );

    \I__13124\ : InMux
    port map (
            O => \N__55950\,
            I => \N__55947\
        );

    \I__13123\ : LocalMux
    port map (
            O => \N__55947\,
            I => \N__55944\
        );

    \I__13122\ : Span4Mux_v
    port map (
            O => \N__55944\,
            I => \N__55940\
        );

    \I__13121\ : InMux
    port map (
            O => \N__55943\,
            I => \N__55937\
        );

    \I__13120\ : Odrv4
    port map (
            O => \N__55940\,
            I => xy_kd_2
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__55937\,
            I => xy_kd_2
        );

    \I__13118\ : InMux
    port map (
            O => \N__55932\,
            I => \N__55928\
        );

    \I__13117\ : InMux
    port map (
            O => \N__55931\,
            I => \N__55923\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__55928\,
            I => \N__55919\
        );

    \I__13115\ : InMux
    port map (
            O => \N__55927\,
            I => \N__55916\
        );

    \I__13114\ : InMux
    port map (
            O => \N__55926\,
            I => \N__55913\
        );

    \I__13113\ : LocalMux
    port map (
            O => \N__55923\,
            I => \N__55910\
        );

    \I__13112\ : InMux
    port map (
            O => \N__55922\,
            I => \N__55907\
        );

    \I__13111\ : Span4Mux_v
    port map (
            O => \N__55919\,
            I => \N__55904\
        );

    \I__13110\ : LocalMux
    port map (
            O => \N__55916\,
            I => \N__55900\
        );

    \I__13109\ : LocalMux
    port map (
            O => \N__55913\,
            I => \N__55895\
        );

    \I__13108\ : Span4Mux_s1_h
    port map (
            O => \N__55910\,
            I => \N__55892\
        );

    \I__13107\ : LocalMux
    port map (
            O => \N__55907\,
            I => \N__55889\
        );

    \I__13106\ : Span4Mux_v
    port map (
            O => \N__55904\,
            I => \N__55886\
        );

    \I__13105\ : InMux
    port map (
            O => \N__55903\,
            I => \N__55883\
        );

    \I__13104\ : Span4Mux_v
    port map (
            O => \N__55900\,
            I => \N__55880\
        );

    \I__13103\ : InMux
    port map (
            O => \N__55899\,
            I => \N__55877\
        );

    \I__13102\ : InMux
    port map (
            O => \N__55898\,
            I => \N__55872\
        );

    \I__13101\ : Span4Mux_v
    port map (
            O => \N__55895\,
            I => \N__55867\
        );

    \I__13100\ : Span4Mux_h
    port map (
            O => \N__55892\,
            I => \N__55867\
        );

    \I__13099\ : Span4Mux_h
    port map (
            O => \N__55889\,
            I => \N__55864\
        );

    \I__13098\ : Span4Mux_v
    port map (
            O => \N__55886\,
            I => \N__55859\
        );

    \I__13097\ : LocalMux
    port map (
            O => \N__55883\,
            I => \N__55859\
        );

    \I__13096\ : Span4Mux_v
    port map (
            O => \N__55880\,
            I => \N__55856\
        );

    \I__13095\ : LocalMux
    port map (
            O => \N__55877\,
            I => \N__55853\
        );

    \I__13094\ : InMux
    port map (
            O => \N__55876\,
            I => \N__55850\
        );

    \I__13093\ : InMux
    port map (
            O => \N__55875\,
            I => \N__55847\
        );

    \I__13092\ : LocalMux
    port map (
            O => \N__55872\,
            I => \N__55842\
        );

    \I__13091\ : Sp12to4
    port map (
            O => \N__55867\,
            I => \N__55839\
        );

    \I__13090\ : Sp12to4
    port map (
            O => \N__55864\,
            I => \N__55836\
        );

    \I__13089\ : Span4Mux_v
    port map (
            O => \N__55859\,
            I => \N__55832\
        );

    \I__13088\ : Span4Mux_v
    port map (
            O => \N__55856\,
            I => \N__55825\
        );

    \I__13087\ : Span4Mux_v
    port map (
            O => \N__55853\,
            I => \N__55825\
        );

    \I__13086\ : LocalMux
    port map (
            O => \N__55850\,
            I => \N__55825\
        );

    \I__13085\ : LocalMux
    port map (
            O => \N__55847\,
            I => \N__55822\
        );

    \I__13084\ : InMux
    port map (
            O => \N__55846\,
            I => \N__55819\
        );

    \I__13083\ : InMux
    port map (
            O => \N__55845\,
            I => \N__55814\
        );

    \I__13082\ : Span4Mux_v
    port map (
            O => \N__55842\,
            I => \N__55811\
        );

    \I__13081\ : Span12Mux_h
    port map (
            O => \N__55839\,
            I => \N__55806\
        );

    \I__13080\ : Span12Mux_v
    port map (
            O => \N__55836\,
            I => \N__55806\
        );

    \I__13079\ : InMux
    port map (
            O => \N__55835\,
            I => \N__55803\
        );

    \I__13078\ : Span4Mux_h
    port map (
            O => \N__55832\,
            I => \N__55794\
        );

    \I__13077\ : Span4Mux_h
    port map (
            O => \N__55825\,
            I => \N__55794\
        );

    \I__13076\ : Span4Mux_v
    port map (
            O => \N__55822\,
            I => \N__55794\
        );

    \I__13075\ : LocalMux
    port map (
            O => \N__55819\,
            I => \N__55794\
        );

    \I__13074\ : InMux
    port map (
            O => \N__55818\,
            I => \N__55789\
        );

    \I__13073\ : InMux
    port map (
            O => \N__55817\,
            I => \N__55789\
        );

    \I__13072\ : LocalMux
    port map (
            O => \N__55814\,
            I => \N__55786\
        );

    \I__13071\ : Odrv4
    port map (
            O => \N__55811\,
            I => uart_pc_data_5
        );

    \I__13070\ : Odrv12
    port map (
            O => \N__55806\,
            I => uart_pc_data_5
        );

    \I__13069\ : LocalMux
    port map (
            O => \N__55803\,
            I => uart_pc_data_5
        );

    \I__13068\ : Odrv4
    port map (
            O => \N__55794\,
            I => uart_pc_data_5
        );

    \I__13067\ : LocalMux
    port map (
            O => \N__55789\,
            I => uart_pc_data_5
        );

    \I__13066\ : Odrv4
    port map (
            O => \N__55786\,
            I => uart_pc_data_5
        );

    \I__13065\ : InMux
    port map (
            O => \N__55773\,
            I => \N__55770\
        );

    \I__13064\ : LocalMux
    port map (
            O => \N__55770\,
            I => \N__55767\
        );

    \I__13063\ : Span4Mux_v
    port map (
            O => \N__55767\,
            I => \N__55763\
        );

    \I__13062\ : InMux
    port map (
            O => \N__55766\,
            I => \N__55760\
        );

    \I__13061\ : Odrv4
    port map (
            O => \N__55763\,
            I => xy_kd_5
        );

    \I__13060\ : LocalMux
    port map (
            O => \N__55760\,
            I => xy_kd_5
        );

    \I__13059\ : InMux
    port map (
            O => \N__55755\,
            I => \N__55751\
        );

    \I__13058\ : InMux
    port map (
            O => \N__55754\,
            I => \N__55746\
        );

    \I__13057\ : LocalMux
    port map (
            O => \N__55751\,
            I => \N__55743\
        );

    \I__13056\ : InMux
    port map (
            O => \N__55750\,
            I => \N__55740\
        );

    \I__13055\ : InMux
    port map (
            O => \N__55749\,
            I => \N__55737\
        );

    \I__13054\ : LocalMux
    port map (
            O => \N__55746\,
            I => \N__55734\
        );

    \I__13053\ : Span4Mux_v
    port map (
            O => \N__55743\,
            I => \N__55727\
        );

    \I__13052\ : LocalMux
    port map (
            O => \N__55740\,
            I => \N__55724\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__55737\,
            I => \N__55720\
        );

    \I__13050\ : Span4Mux_v
    port map (
            O => \N__55734\,
            I => \N__55717\
        );

    \I__13049\ : InMux
    port map (
            O => \N__55733\,
            I => \N__55713\
        );

    \I__13048\ : InMux
    port map (
            O => \N__55732\,
            I => \N__55710\
        );

    \I__13047\ : InMux
    port map (
            O => \N__55731\,
            I => \N__55706\
        );

    \I__13046\ : InMux
    port map (
            O => \N__55730\,
            I => \N__55702\
        );

    \I__13045\ : Sp12to4
    port map (
            O => \N__55727\,
            I => \N__55699\
        );

    \I__13044\ : Span4Mux_v
    port map (
            O => \N__55724\,
            I => \N__55696\
        );

    \I__13043\ : InMux
    port map (
            O => \N__55723\,
            I => \N__55693\
        );

    \I__13042\ : Span4Mux_v
    port map (
            O => \N__55720\,
            I => \N__55688\
        );

    \I__13041\ : Span4Mux_h
    port map (
            O => \N__55717\,
            I => \N__55688\
        );

    \I__13040\ : InMux
    port map (
            O => \N__55716\,
            I => \N__55685\
        );

    \I__13039\ : LocalMux
    port map (
            O => \N__55713\,
            I => \N__55682\
        );

    \I__13038\ : LocalMux
    port map (
            O => \N__55710\,
            I => \N__55679\
        );

    \I__13037\ : InMux
    port map (
            O => \N__55709\,
            I => \N__55676\
        );

    \I__13036\ : LocalMux
    port map (
            O => \N__55706\,
            I => \N__55673\
        );

    \I__13035\ : InMux
    port map (
            O => \N__55705\,
            I => \N__55670\
        );

    \I__13034\ : LocalMux
    port map (
            O => \N__55702\,
            I => \N__55667\
        );

    \I__13033\ : Span12Mux_h
    port map (
            O => \N__55699\,
            I => \N__55659\
        );

    \I__13032\ : Sp12to4
    port map (
            O => \N__55696\,
            I => \N__55659\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__55693\,
            I => \N__55659\
        );

    \I__13030\ : Sp12to4
    port map (
            O => \N__55688\,
            I => \N__55656\
        );

    \I__13029\ : LocalMux
    port map (
            O => \N__55685\,
            I => \N__55653\
        );

    \I__13028\ : Span4Mux_v
    port map (
            O => \N__55682\,
            I => \N__55650\
        );

    \I__13027\ : Span4Mux_v
    port map (
            O => \N__55679\,
            I => \N__55647\
        );

    \I__13026\ : LocalMux
    port map (
            O => \N__55676\,
            I => \N__55644\
        );

    \I__13025\ : Span4Mux_h
    port map (
            O => \N__55673\,
            I => \N__55639\
        );

    \I__13024\ : LocalMux
    port map (
            O => \N__55670\,
            I => \N__55639\
        );

    \I__13023\ : Span4Mux_h
    port map (
            O => \N__55667\,
            I => \N__55636\
        );

    \I__13022\ : InMux
    port map (
            O => \N__55666\,
            I => \N__55633\
        );

    \I__13021\ : Span12Mux_v
    port map (
            O => \N__55659\,
            I => \N__55630\
        );

    \I__13020\ : Span12Mux_h
    port map (
            O => \N__55656\,
            I => \N__55625\
        );

    \I__13019\ : Span12Mux_s7_h
    port map (
            O => \N__55653\,
            I => \N__55625\
        );

    \I__13018\ : Span4Mux_h
    port map (
            O => \N__55650\,
            I => \N__55616\
        );

    \I__13017\ : Span4Mux_h
    port map (
            O => \N__55647\,
            I => \N__55616\
        );

    \I__13016\ : Span4Mux_v
    port map (
            O => \N__55644\,
            I => \N__55616\
        );

    \I__13015\ : Span4Mux_v
    port map (
            O => \N__55639\,
            I => \N__55616\
        );

    \I__13014\ : Odrv4
    port map (
            O => \N__55636\,
            I => uart_pc_data_6
        );

    \I__13013\ : LocalMux
    port map (
            O => \N__55633\,
            I => uart_pc_data_6
        );

    \I__13012\ : Odrv12
    port map (
            O => \N__55630\,
            I => uart_pc_data_6
        );

    \I__13011\ : Odrv12
    port map (
            O => \N__55625\,
            I => uart_pc_data_6
        );

    \I__13010\ : Odrv4
    port map (
            O => \N__55616\,
            I => uart_pc_data_6
        );

    \I__13009\ : InMux
    port map (
            O => \N__55605\,
            I => \N__55602\
        );

    \I__13008\ : LocalMux
    port map (
            O => \N__55602\,
            I => \N__55599\
        );

    \I__13007\ : Span4Mux_s0_h
    port map (
            O => \N__55599\,
            I => \N__55596\
        );

    \I__13006\ : Span4Mux_v
    port map (
            O => \N__55596\,
            I => \N__55592\
        );

    \I__13005\ : InMux
    port map (
            O => \N__55595\,
            I => \N__55589\
        );

    \I__13004\ : Odrv4
    port map (
            O => \N__55592\,
            I => xy_kd_6
        );

    \I__13003\ : LocalMux
    port map (
            O => \N__55589\,
            I => xy_kd_6
        );

    \I__13002\ : InMux
    port map (
            O => \N__55584\,
            I => \N__55578\
        );

    \I__13001\ : InMux
    port map (
            O => \N__55583\,
            I => \N__55575\
        );

    \I__13000\ : InMux
    port map (
            O => \N__55582\,
            I => \N__55571\
        );

    \I__12999\ : InMux
    port map (
            O => \N__55581\,
            I => \N__55568\
        );

    \I__12998\ : LocalMux
    port map (
            O => \N__55578\,
            I => \N__55562\
        );

    \I__12997\ : LocalMux
    port map (
            O => \N__55575\,
            I => \N__55559\
        );

    \I__12996\ : InMux
    port map (
            O => \N__55574\,
            I => \N__55556\
        );

    \I__12995\ : LocalMux
    port map (
            O => \N__55571\,
            I => \N__55553\
        );

    \I__12994\ : LocalMux
    port map (
            O => \N__55568\,
            I => \N__55550\
        );

    \I__12993\ : InMux
    port map (
            O => \N__55567\,
            I => \N__55545\
        );

    \I__12992\ : InMux
    port map (
            O => \N__55566\,
            I => \N__55542\
        );

    \I__12991\ : InMux
    port map (
            O => \N__55565\,
            I => \N__55538\
        );

    \I__12990\ : Span4Mux_v
    port map (
            O => \N__55562\,
            I => \N__55535\
        );

    \I__12989\ : Span4Mux_s3_h
    port map (
            O => \N__55559\,
            I => \N__55531\
        );

    \I__12988\ : LocalMux
    port map (
            O => \N__55556\,
            I => \N__55528\
        );

    \I__12987\ : Span4Mux_v
    port map (
            O => \N__55553\,
            I => \N__55525\
        );

    \I__12986\ : Span4Mux_v
    port map (
            O => \N__55550\,
            I => \N__55522\
        );

    \I__12985\ : InMux
    port map (
            O => \N__55549\,
            I => \N__55518\
        );

    \I__12984\ : InMux
    port map (
            O => \N__55548\,
            I => \N__55515\
        );

    \I__12983\ : LocalMux
    port map (
            O => \N__55545\,
            I => \N__55512\
        );

    \I__12982\ : LocalMux
    port map (
            O => \N__55542\,
            I => \N__55509\
        );

    \I__12981\ : InMux
    port map (
            O => \N__55541\,
            I => \N__55506\
        );

    \I__12980\ : LocalMux
    port map (
            O => \N__55538\,
            I => \N__55503\
        );

    \I__12979\ : Span4Mux_h
    port map (
            O => \N__55535\,
            I => \N__55500\
        );

    \I__12978\ : CascadeMux
    port map (
            O => \N__55534\,
            I => \N__55497\
        );

    \I__12977\ : Span4Mux_h
    port map (
            O => \N__55531\,
            I => \N__55494\
        );

    \I__12976\ : Span4Mux_v
    port map (
            O => \N__55528\,
            I => \N__55489\
        );

    \I__12975\ : Span4Mux_h
    port map (
            O => \N__55525\,
            I => \N__55489\
        );

    \I__12974\ : Span4Mux_h
    port map (
            O => \N__55522\,
            I => \N__55486\
        );

    \I__12973\ : InMux
    port map (
            O => \N__55521\,
            I => \N__55483\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__55518\,
            I => \N__55480\
        );

    \I__12971\ : LocalMux
    port map (
            O => \N__55515\,
            I => \N__55477\
        );

    \I__12970\ : Span4Mux_v
    port map (
            O => \N__55512\,
            I => \N__55474\
        );

    \I__12969\ : Span4Mux_v
    port map (
            O => \N__55509\,
            I => \N__55471\
        );

    \I__12968\ : LocalMux
    port map (
            O => \N__55506\,
            I => \N__55468\
        );

    \I__12967\ : Span4Mux_s3_h
    port map (
            O => \N__55503\,
            I => \N__55465\
        );

    \I__12966\ : Span4Mux_v
    port map (
            O => \N__55500\,
            I => \N__55462\
        );

    \I__12965\ : InMux
    port map (
            O => \N__55497\,
            I => \N__55459\
        );

    \I__12964\ : Sp12to4
    port map (
            O => \N__55494\,
            I => \N__55456\
        );

    \I__12963\ : Span4Mux_v
    port map (
            O => \N__55489\,
            I => \N__55453\
        );

    \I__12962\ : Span4Mux_v
    port map (
            O => \N__55486\,
            I => \N__55450\
        );

    \I__12961\ : LocalMux
    port map (
            O => \N__55483\,
            I => \N__55447\
        );

    \I__12960\ : Span4Mux_v
    port map (
            O => \N__55480\,
            I => \N__55436\
        );

    \I__12959\ : Span4Mux_v
    port map (
            O => \N__55477\,
            I => \N__55436\
        );

    \I__12958\ : Span4Mux_h
    port map (
            O => \N__55474\,
            I => \N__55436\
        );

    \I__12957\ : Span4Mux_h
    port map (
            O => \N__55471\,
            I => \N__55436\
        );

    \I__12956\ : Span4Mux_h
    port map (
            O => \N__55468\,
            I => \N__55431\
        );

    \I__12955\ : Span4Mux_h
    port map (
            O => \N__55465\,
            I => \N__55431\
        );

    \I__12954\ : Span4Mux_v
    port map (
            O => \N__55462\,
            I => \N__55428\
        );

    \I__12953\ : LocalMux
    port map (
            O => \N__55459\,
            I => \N__55421\
        );

    \I__12952\ : Span12Mux_v
    port map (
            O => \N__55456\,
            I => \N__55421\
        );

    \I__12951\ : Sp12to4
    port map (
            O => \N__55453\,
            I => \N__55421\
        );

    \I__12950\ : Span4Mux_v
    port map (
            O => \N__55450\,
            I => \N__55416\
        );

    \I__12949\ : Span4Mux_h
    port map (
            O => \N__55447\,
            I => \N__55416\
        );

    \I__12948\ : InMux
    port map (
            O => \N__55446\,
            I => \N__55413\
        );

    \I__12947\ : InMux
    port map (
            O => \N__55445\,
            I => \N__55410\
        );

    \I__12946\ : Odrv4
    port map (
            O => \N__55436\,
            I => uart_pc_data_7
        );

    \I__12945\ : Odrv4
    port map (
            O => \N__55431\,
            I => uart_pc_data_7
        );

    \I__12944\ : Odrv4
    port map (
            O => \N__55428\,
            I => uart_pc_data_7
        );

    \I__12943\ : Odrv12
    port map (
            O => \N__55421\,
            I => uart_pc_data_7
        );

    \I__12942\ : Odrv4
    port map (
            O => \N__55416\,
            I => uart_pc_data_7
        );

    \I__12941\ : LocalMux
    port map (
            O => \N__55413\,
            I => uart_pc_data_7
        );

    \I__12940\ : LocalMux
    port map (
            O => \N__55410\,
            I => uart_pc_data_7
        );

    \I__12939\ : InMux
    port map (
            O => \N__55395\,
            I => \N__55392\
        );

    \I__12938\ : LocalMux
    port map (
            O => \N__55392\,
            I => \N__55389\
        );

    \I__12937\ : Span4Mux_v
    port map (
            O => \N__55389\,
            I => \N__55385\
        );

    \I__12936\ : InMux
    port map (
            O => \N__55388\,
            I => \N__55382\
        );

    \I__12935\ : Odrv4
    port map (
            O => \N__55385\,
            I => xy_kd_7
        );

    \I__12934\ : LocalMux
    port map (
            O => \N__55382\,
            I => xy_kd_7
        );

    \I__12933\ : InMux
    port map (
            O => \N__55377\,
            I => \N__55374\
        );

    \I__12932\ : LocalMux
    port map (
            O => \N__55374\,
            I => \N__55369\
        );

    \I__12931\ : InMux
    port map (
            O => \N__55373\,
            I => \N__55366\
        );

    \I__12930\ : InMux
    port map (
            O => \N__55372\,
            I => \N__55363\
        );

    \I__12929\ : Span4Mux_v
    port map (
            O => \N__55369\,
            I => \N__55357\
        );

    \I__12928\ : LocalMux
    port map (
            O => \N__55366\,
            I => \N__55357\
        );

    \I__12927\ : LocalMux
    port map (
            O => \N__55363\,
            I => \N__55350\
        );

    \I__12926\ : InMux
    port map (
            O => \N__55362\,
            I => \N__55347\
        );

    \I__12925\ : Span4Mux_v
    port map (
            O => \N__55357\,
            I => \N__55344\
        );

    \I__12924\ : InMux
    port map (
            O => \N__55356\,
            I => \N__55339\
        );

    \I__12923\ : InMux
    port map (
            O => \N__55355\,
            I => \N__55336\
        );

    \I__12922\ : InMux
    port map (
            O => \N__55354\,
            I => \N__55333\
        );

    \I__12921\ : InMux
    port map (
            O => \N__55353\,
            I => \N__55329\
        );

    \I__12920\ : Span4Mux_v
    port map (
            O => \N__55350\,
            I => \N__55326\
        );

    \I__12919\ : LocalMux
    port map (
            O => \N__55347\,
            I => \N__55323\
        );

    \I__12918\ : Span4Mux_h
    port map (
            O => \N__55344\,
            I => \N__55320\
        );

    \I__12917\ : InMux
    port map (
            O => \N__55343\,
            I => \N__55317\
        );

    \I__12916\ : InMux
    port map (
            O => \N__55342\,
            I => \N__55314\
        );

    \I__12915\ : LocalMux
    port map (
            O => \N__55339\,
            I => \N__55311\
        );

    \I__12914\ : LocalMux
    port map (
            O => \N__55336\,
            I => \N__55308\
        );

    \I__12913\ : LocalMux
    port map (
            O => \N__55333\,
            I => \N__55305\
        );

    \I__12912\ : InMux
    port map (
            O => \N__55332\,
            I => \N__55302\
        );

    \I__12911\ : LocalMux
    port map (
            O => \N__55329\,
            I => \N__55299\
        );

    \I__12910\ : Span4Mux_v
    port map (
            O => \N__55326\,
            I => \N__55296\
        );

    \I__12909\ : Sp12to4
    port map (
            O => \N__55323\,
            I => \N__55293\
        );

    \I__12908\ : Span4Mux_v
    port map (
            O => \N__55320\,
            I => \N__55290\
        );

    \I__12907\ : LocalMux
    port map (
            O => \N__55317\,
            I => \N__55285\
        );

    \I__12906\ : LocalMux
    port map (
            O => \N__55314\,
            I => \N__55285\
        );

    \I__12905\ : Span12Mux_h
    port map (
            O => \N__55311\,
            I => \N__55281\
        );

    \I__12904\ : Span4Mux_v
    port map (
            O => \N__55308\,
            I => \N__55273\
        );

    \I__12903\ : Span4Mux_s3_h
    port map (
            O => \N__55305\,
            I => \N__55273\
        );

    \I__12902\ : LocalMux
    port map (
            O => \N__55302\,
            I => \N__55273\
        );

    \I__12901\ : Span4Mux_v
    port map (
            O => \N__55299\,
            I => \N__55270\
        );

    \I__12900\ : Sp12to4
    port map (
            O => \N__55296\,
            I => \N__55265\
        );

    \I__12899\ : Span12Mux_v
    port map (
            O => \N__55293\,
            I => \N__55265\
        );

    \I__12898\ : Span4Mux_v
    port map (
            O => \N__55290\,
            I => \N__55260\
        );

    \I__12897\ : Span4Mux_v
    port map (
            O => \N__55285\,
            I => \N__55260\
        );

    \I__12896\ : InMux
    port map (
            O => \N__55284\,
            I => \N__55257\
        );

    \I__12895\ : Span12Mux_v
    port map (
            O => \N__55281\,
            I => \N__55254\
        );

    \I__12894\ : InMux
    port map (
            O => \N__55280\,
            I => \N__55251\
        );

    \I__12893\ : Span4Mux_h
    port map (
            O => \N__55273\,
            I => \N__55248\
        );

    \I__12892\ : Sp12to4
    port map (
            O => \N__55270\,
            I => \N__55239\
        );

    \I__12891\ : Span12Mux_h
    port map (
            O => \N__55265\,
            I => \N__55239\
        );

    \I__12890\ : Sp12to4
    port map (
            O => \N__55260\,
            I => \N__55239\
        );

    \I__12889\ : LocalMux
    port map (
            O => \N__55257\,
            I => \N__55239\
        );

    \I__12888\ : Odrv12
    port map (
            O => \N__55254\,
            I => uart_pc_data_3
        );

    \I__12887\ : LocalMux
    port map (
            O => \N__55251\,
            I => uart_pc_data_3
        );

    \I__12886\ : Odrv4
    port map (
            O => \N__55248\,
            I => uart_pc_data_3
        );

    \I__12885\ : Odrv12
    port map (
            O => \N__55239\,
            I => uart_pc_data_3
        );

    \I__12884\ : InMux
    port map (
            O => \N__55230\,
            I => \N__55227\
        );

    \I__12883\ : LocalMux
    port map (
            O => \N__55227\,
            I => \N__55224\
        );

    \I__12882\ : Span4Mux_v
    port map (
            O => \N__55224\,
            I => \N__55220\
        );

    \I__12881\ : InMux
    port map (
            O => \N__55223\,
            I => \N__55217\
        );

    \I__12880\ : Odrv4
    port map (
            O => \N__55220\,
            I => xy_kd_3
        );

    \I__12879\ : LocalMux
    port map (
            O => \N__55217\,
            I => xy_kd_3
        );

    \I__12878\ : CEMux
    port map (
            O => \N__55212\,
            I => \N__55209\
        );

    \I__12877\ : LocalMux
    port map (
            O => \N__55209\,
            I => \N__55206\
        );

    \I__12876\ : Span4Mux_s3_h
    port map (
            O => \N__55206\,
            I => \N__55202\
        );

    \I__12875\ : CEMux
    port map (
            O => \N__55205\,
            I => \N__55199\
        );

    \I__12874\ : Span4Mux_h
    port map (
            O => \N__55202\,
            I => \N__55194\
        );

    \I__12873\ : LocalMux
    port map (
            O => \N__55199\,
            I => \N__55194\
        );

    \I__12872\ : Span4Mux_v
    port map (
            O => \N__55194\,
            I => \N__55191\
        );

    \I__12871\ : Span4Mux_h
    port map (
            O => \N__55191\,
            I => \N__55188\
        );

    \I__12870\ : Span4Mux_h
    port map (
            O => \N__55188\,
            I => \N__55185\
        );

    \I__12869\ : Span4Mux_h
    port map (
            O => \N__55185\,
            I => \N__55182\
        );

    \I__12868\ : Odrv4
    port map (
            O => \N__55182\,
            I => \Commands_frame_decoder.state_RNITUI31Z0Z_13\
        );

    \I__12867\ : InMux
    port map (
            O => \N__55179\,
            I => \N__55176\
        );

    \I__12866\ : LocalMux
    port map (
            O => \N__55176\,
            I => \N__55173\
        );

    \I__12865\ : Odrv4
    port map (
            O => \N__55173\,
            I => \pid_side.O_1_18\
        );

    \I__12864\ : InMux
    port map (
            O => \N__55170\,
            I => \N__55165\
        );

    \I__12863\ : InMux
    port map (
            O => \N__55169\,
            I => \N__55162\
        );

    \I__12862\ : InMux
    port map (
            O => \N__55168\,
            I => \N__55159\
        );

    \I__12861\ : LocalMux
    port map (
            O => \N__55165\,
            I => \N__55154\
        );

    \I__12860\ : LocalMux
    port map (
            O => \N__55162\,
            I => \N__55154\
        );

    \I__12859\ : LocalMux
    port map (
            O => \N__55159\,
            I => \N__55151\
        );

    \I__12858\ : Span4Mux_h
    port map (
            O => \N__55154\,
            I => \N__55148\
        );

    \I__12857\ : Span4Mux_h
    port map (
            O => \N__55151\,
            I => \N__55145\
        );

    \I__12856\ : Odrv4
    port map (
            O => \N__55148\,
            I => \pid_side.error_d_regZ0Z_14\
        );

    \I__12855\ : Odrv4
    port map (
            O => \N__55145\,
            I => \pid_side.error_d_regZ0Z_14\
        );

    \I__12854\ : InMux
    port map (
            O => \N__55140\,
            I => \N__55137\
        );

    \I__12853\ : LocalMux
    port map (
            O => \N__55137\,
            I => \pid_side.O_1_7\
        );

    \I__12852\ : InMux
    port map (
            O => \N__55134\,
            I => \N__55125\
        );

    \I__12851\ : InMux
    port map (
            O => \N__55133\,
            I => \N__55125\
        );

    \I__12850\ : InMux
    port map (
            O => \N__55132\,
            I => \N__55125\
        );

    \I__12849\ : LocalMux
    port map (
            O => \N__55125\,
            I => \N__55122\
        );

    \I__12848\ : Span4Mux_v
    port map (
            O => \N__55122\,
            I => \N__55119\
        );

    \I__12847\ : Odrv4
    port map (
            O => \N__55119\,
            I => \pid_side.error_d_regZ0Z_3\
        );

    \I__12846\ : InMux
    port map (
            O => \N__55116\,
            I => \N__55113\
        );

    \I__12845\ : LocalMux
    port map (
            O => \N__55113\,
            I => \N__55110\
        );

    \I__12844\ : Span4Mux_h
    port map (
            O => \N__55110\,
            I => \N__55107\
        );

    \I__12843\ : Odrv4
    port map (
            O => \N__55107\,
            I => \pid_side.O_1_17\
        );

    \I__12842\ : InMux
    port map (
            O => \N__55104\,
            I => \N__55095\
        );

    \I__12841\ : InMux
    port map (
            O => \N__55103\,
            I => \N__55095\
        );

    \I__12840\ : InMux
    port map (
            O => \N__55102\,
            I => \N__55095\
        );

    \I__12839\ : LocalMux
    port map (
            O => \N__55095\,
            I => \N__55092\
        );

    \I__12838\ : Span12Mux_v
    port map (
            O => \N__55092\,
            I => \N__55089\
        );

    \I__12837\ : Odrv12
    port map (
            O => \N__55089\,
            I => \pid_side.error_d_regZ0Z_13\
        );

    \I__12836\ : InMux
    port map (
            O => \N__55086\,
            I => \N__55083\
        );

    \I__12835\ : LocalMux
    port map (
            O => \N__55083\,
            I => \pid_side.O_1_14\
        );

    \I__12834\ : InMux
    port map (
            O => \N__55080\,
            I => \N__55075\
        );

    \I__12833\ : InMux
    port map (
            O => \N__55079\,
            I => \N__55070\
        );

    \I__12832\ : InMux
    port map (
            O => \N__55078\,
            I => \N__55070\
        );

    \I__12831\ : LocalMux
    port map (
            O => \N__55075\,
            I => \N__55067\
        );

    \I__12830\ : LocalMux
    port map (
            O => \N__55070\,
            I => \N__55064\
        );

    \I__12829\ : Span4Mux_v
    port map (
            O => \N__55067\,
            I => \N__55061\
        );

    \I__12828\ : Span4Mux_h
    port map (
            O => \N__55064\,
            I => \N__55058\
        );

    \I__12827\ : Odrv4
    port map (
            O => \N__55061\,
            I => \pid_side.error_d_regZ0Z_10\
        );

    \I__12826\ : Odrv4
    port map (
            O => \N__55058\,
            I => \pid_side.error_d_regZ0Z_10\
        );

    \I__12825\ : InMux
    port map (
            O => \N__55053\,
            I => \N__55050\
        );

    \I__12824\ : LocalMux
    port map (
            O => \N__55050\,
            I => \N__55047\
        );

    \I__12823\ : Odrv4
    port map (
            O => \N__55047\,
            I => \pid_side.O_1_23\
        );

    \I__12822\ : InMux
    port map (
            O => \N__55044\,
            I => \N__55035\
        );

    \I__12821\ : InMux
    port map (
            O => \N__55043\,
            I => \N__55035\
        );

    \I__12820\ : InMux
    port map (
            O => \N__55042\,
            I => \N__55035\
        );

    \I__12819\ : LocalMux
    port map (
            O => \N__55035\,
            I => \N__55032\
        );

    \I__12818\ : Odrv12
    port map (
            O => \N__55032\,
            I => \pid_side.error_d_regZ0Z_19\
        );

    \I__12817\ : InMux
    port map (
            O => \N__55029\,
            I => \N__55026\
        );

    \I__12816\ : LocalMux
    port map (
            O => \N__55026\,
            I => \N__55023\
        );

    \I__12815\ : Odrv4
    port map (
            O => \N__55023\,
            I => \pid_side.O_1_24\
        );

    \I__12814\ : InMux
    port map (
            O => \N__55020\,
            I => \N__55017\
        );

    \I__12813\ : LocalMux
    port map (
            O => \N__55017\,
            I => \pid_side.O_1_10\
        );

    \I__12812\ : InMux
    port map (
            O => \N__55014\,
            I => \N__55011\
        );

    \I__12811\ : LocalMux
    port map (
            O => \N__55011\,
            I => \N__55006\
        );

    \I__12810\ : InMux
    port map (
            O => \N__55010\,
            I => \N__55001\
        );

    \I__12809\ : InMux
    port map (
            O => \N__55009\,
            I => \N__55001\
        );

    \I__12808\ : Span4Mux_h
    port map (
            O => \N__55006\,
            I => \N__54996\
        );

    \I__12807\ : LocalMux
    port map (
            O => \N__55001\,
            I => \N__54996\
        );

    \I__12806\ : Odrv4
    port map (
            O => \N__54996\,
            I => \pid_side.error_d_regZ0Z_6\
        );

    \I__12805\ : InMux
    port map (
            O => \N__54993\,
            I => \N__54990\
        );

    \I__12804\ : LocalMux
    port map (
            O => \N__54990\,
            I => \N__54987\
        );

    \I__12803\ : Odrv4
    port map (
            O => \N__54987\,
            I => \pid_side.O_1_22\
        );

    \I__12802\ : InMux
    port map (
            O => \N__54984\,
            I => \N__54975\
        );

    \I__12801\ : InMux
    port map (
            O => \N__54983\,
            I => \N__54975\
        );

    \I__12800\ : InMux
    port map (
            O => \N__54982\,
            I => \N__54975\
        );

    \I__12799\ : LocalMux
    port map (
            O => \N__54975\,
            I => \N__54972\
        );

    \I__12798\ : Span4Mux_h
    port map (
            O => \N__54972\,
            I => \N__54969\
        );

    \I__12797\ : Odrv4
    port map (
            O => \N__54969\,
            I => \pid_side.error_d_regZ0Z_18\
        );

    \I__12796\ : InMux
    port map (
            O => \N__54966\,
            I => \N__54963\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__54963\,
            I => \pid_side.O_1_11\
        );

    \I__12794\ : InMux
    port map (
            O => \N__54960\,
            I => \N__54954\
        );

    \I__12793\ : InMux
    port map (
            O => \N__54959\,
            I => \N__54947\
        );

    \I__12792\ : InMux
    port map (
            O => \N__54958\,
            I => \N__54947\
        );

    \I__12791\ : InMux
    port map (
            O => \N__54957\,
            I => \N__54947\
        );

    \I__12790\ : LocalMux
    port map (
            O => \N__54954\,
            I => \pid_side.error_d_reg_prevZ0Z_7\
        );

    \I__12789\ : LocalMux
    port map (
            O => \N__54947\,
            I => \pid_side.error_d_reg_prevZ0Z_7\
        );

    \I__12788\ : InMux
    port map (
            O => \N__54942\,
            I => \N__54939\
        );

    \I__12787\ : LocalMux
    port map (
            O => \N__54939\,
            I => \N__54936\
        );

    \I__12786\ : Span4Mux_h
    port map (
            O => \N__54936\,
            I => \N__54933\
        );

    \I__12785\ : Odrv4
    port map (
            O => \N__54933\,
            I => \pid_side.error_p_reg_esr_RNIBNBR2Z0Z_7\
        );

    \I__12784\ : InMux
    port map (
            O => \N__54930\,
            I => \N__54924\
        );

    \I__12783\ : InMux
    port map (
            O => \N__54929\,
            I => \N__54917\
        );

    \I__12782\ : InMux
    port map (
            O => \N__54928\,
            I => \N__54917\
        );

    \I__12781\ : InMux
    port map (
            O => \N__54927\,
            I => \N__54917\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__54924\,
            I => \pid_side.error_p_regZ0Z_6\
        );

    \I__12779\ : LocalMux
    port map (
            O => \N__54917\,
            I => \pid_side.error_p_regZ0Z_6\
        );

    \I__12778\ : InMux
    port map (
            O => \N__54912\,
            I => \N__54906\
        );

    \I__12777\ : InMux
    port map (
            O => \N__54911\,
            I => \N__54899\
        );

    \I__12776\ : InMux
    port map (
            O => \N__54910\,
            I => \N__54899\
        );

    \I__12775\ : InMux
    port map (
            O => \N__54909\,
            I => \N__54899\
        );

    \I__12774\ : LocalMux
    port map (
            O => \N__54906\,
            I => \pid_side.error_d_reg_prevZ0Z_6\
        );

    \I__12773\ : LocalMux
    port map (
            O => \N__54899\,
            I => \pid_side.error_d_reg_prevZ0Z_6\
        );

    \I__12772\ : InMux
    port map (
            O => \N__54894\,
            I => \N__54891\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__54891\,
            I => \N__54888\
        );

    \I__12770\ : Span12Mux_h
    port map (
            O => \N__54888\,
            I => \N__54885\
        );

    \I__12769\ : Odrv12
    port map (
            O => \N__54885\,
            I => \pid_side.un1_pid_prereg_50_0\
        );

    \I__12768\ : InMux
    port map (
            O => \N__54882\,
            I => \N__54879\
        );

    \I__12767\ : LocalMux
    port map (
            O => \N__54879\,
            I => \N__54876\
        );

    \I__12766\ : Span4Mux_h
    port map (
            O => \N__54876\,
            I => \N__54873\
        );

    \I__12765\ : Odrv4
    port map (
            O => \N__54873\,
            I => \pid_side.O_1_15\
        );

    \I__12764\ : InMux
    port map (
            O => \N__54870\,
            I => \N__54865\
        );

    \I__12763\ : InMux
    port map (
            O => \N__54869\,
            I => \N__54860\
        );

    \I__12762\ : InMux
    port map (
            O => \N__54868\,
            I => \N__54860\
        );

    \I__12761\ : LocalMux
    port map (
            O => \N__54865\,
            I => \N__54857\
        );

    \I__12760\ : LocalMux
    port map (
            O => \N__54860\,
            I => \N__54854\
        );

    \I__12759\ : Span4Mux_h
    port map (
            O => \N__54857\,
            I => \N__54851\
        );

    \I__12758\ : Odrv4
    port map (
            O => \N__54854\,
            I => \pid_side.error_d_regZ0Z_11\
        );

    \I__12757\ : Odrv4
    port map (
            O => \N__54851\,
            I => \pid_side.error_d_regZ0Z_11\
        );

    \I__12756\ : InMux
    port map (
            O => \N__54846\,
            I => \N__54843\
        );

    \I__12755\ : LocalMux
    port map (
            O => \N__54843\,
            I => \N__54840\
        );

    \I__12754\ : Odrv4
    port map (
            O => \N__54840\,
            I => \pid_side.O_1_21\
        );

    \I__12753\ : InMux
    port map (
            O => \N__54837\,
            I => \N__54832\
        );

    \I__12752\ : InMux
    port map (
            O => \N__54836\,
            I => \N__54827\
        );

    \I__12751\ : InMux
    port map (
            O => \N__54835\,
            I => \N__54827\
        );

    \I__12750\ : LocalMux
    port map (
            O => \N__54832\,
            I => \pid_side.error_d_regZ0Z_17\
        );

    \I__12749\ : LocalMux
    port map (
            O => \N__54827\,
            I => \pid_side.error_d_regZ0Z_17\
        );

    \I__12748\ : InMux
    port map (
            O => \N__54822\,
            I => \N__54819\
        );

    \I__12747\ : LocalMux
    port map (
            O => \N__54819\,
            I => \N__54816\
        );

    \I__12746\ : Odrv4
    port map (
            O => \N__54816\,
            I => \pid_side.O_1_19\
        );

    \I__12745\ : InMux
    port map (
            O => \N__54813\,
            I => \N__54809\
        );

    \I__12744\ : InMux
    port map (
            O => \N__54812\,
            I => \N__54805\
        );

    \I__12743\ : LocalMux
    port map (
            O => \N__54809\,
            I => \N__54802\
        );

    \I__12742\ : InMux
    port map (
            O => \N__54808\,
            I => \N__54799\
        );

    \I__12741\ : LocalMux
    port map (
            O => \N__54805\,
            I => \N__54792\
        );

    \I__12740\ : Span4Mux_h
    port map (
            O => \N__54802\,
            I => \N__54792\
        );

    \I__12739\ : LocalMux
    port map (
            O => \N__54799\,
            I => \N__54792\
        );

    \I__12738\ : Span4Mux_h
    port map (
            O => \N__54792\,
            I => \N__54789\
        );

    \I__12737\ : Odrv4
    port map (
            O => \N__54789\,
            I => \pid_side.error_d_regZ0Z_15\
        );

    \I__12736\ : InMux
    port map (
            O => \N__54786\,
            I => \N__54783\
        );

    \I__12735\ : LocalMux
    port map (
            O => \N__54783\,
            I => \N__54780\
        );

    \I__12734\ : Odrv4
    port map (
            O => \N__54780\,
            I => \pid_side.O_1_12\
        );

    \I__12733\ : InMux
    port map (
            O => \N__54777\,
            I => \N__54768\
        );

    \I__12732\ : InMux
    port map (
            O => \N__54776\,
            I => \N__54768\
        );

    \I__12731\ : InMux
    port map (
            O => \N__54775\,
            I => \N__54768\
        );

    \I__12730\ : LocalMux
    port map (
            O => \N__54768\,
            I => \N__54765\
        );

    \I__12729\ : Odrv4
    port map (
            O => \N__54765\,
            I => \pid_side.error_d_regZ0Z_8\
        );

    \I__12728\ : InMux
    port map (
            O => \N__54762\,
            I => \N__54759\
        );

    \I__12727\ : LocalMux
    port map (
            O => \N__54759\,
            I => \N__54756\
        );

    \I__12726\ : Odrv4
    port map (
            O => \N__54756\,
            I => \pid_side.O_1_9\
        );

    \I__12725\ : InMux
    port map (
            O => \N__54753\,
            I => \N__54748\
        );

    \I__12724\ : InMux
    port map (
            O => \N__54752\,
            I => \N__54743\
        );

    \I__12723\ : InMux
    port map (
            O => \N__54751\,
            I => \N__54743\
        );

    \I__12722\ : LocalMux
    port map (
            O => \N__54748\,
            I => \N__54740\
        );

    \I__12721\ : LocalMux
    port map (
            O => \N__54743\,
            I => \N__54737\
        );

    \I__12720\ : Span4Mux_h
    port map (
            O => \N__54740\,
            I => \N__54734\
        );

    \I__12719\ : Span4Mux_h
    port map (
            O => \N__54737\,
            I => \N__54731\
        );

    \I__12718\ : Span4Mux_v
    port map (
            O => \N__54734\,
            I => \N__54728\
        );

    \I__12717\ : Span4Mux_v
    port map (
            O => \N__54731\,
            I => \N__54725\
        );

    \I__12716\ : Odrv4
    port map (
            O => \N__54728\,
            I => \pid_side.error_d_regZ0Z_5\
        );

    \I__12715\ : Odrv4
    port map (
            O => \N__54725\,
            I => \pid_side.error_d_regZ0Z_5\
        );

    \I__12714\ : InMux
    port map (
            O => \N__54720\,
            I => \N__54717\
        );

    \I__12713\ : LocalMux
    port map (
            O => \N__54717\,
            I => \N__54714\
        );

    \I__12712\ : Odrv4
    port map (
            O => \N__54714\,
            I => \pid_side.O_1_16\
        );

    \I__12711\ : InMux
    port map (
            O => \N__54711\,
            I => \N__54702\
        );

    \I__12710\ : InMux
    port map (
            O => \N__54710\,
            I => \N__54702\
        );

    \I__12709\ : InMux
    port map (
            O => \N__54709\,
            I => \N__54702\
        );

    \I__12708\ : LocalMux
    port map (
            O => \N__54702\,
            I => \N__54699\
        );

    \I__12707\ : Span4Mux_h
    port map (
            O => \N__54699\,
            I => \N__54696\
        );

    \I__12706\ : Odrv4
    port map (
            O => \N__54696\,
            I => \pid_side.error_d_regZ0Z_12\
        );

    \I__12705\ : InMux
    port map (
            O => \N__54693\,
            I => \N__54690\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__54690\,
            I => \pid_side.O_2_11\
        );

    \I__12703\ : InMux
    port map (
            O => \N__54687\,
            I => \N__54684\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__54684\,
            I => \pid_side.O_2_23\
        );

    \I__12701\ : InMux
    port map (
            O => \N__54681\,
            I => \N__54675\
        );

    \I__12700\ : InMux
    port map (
            O => \N__54680\,
            I => \N__54675\
        );

    \I__12699\ : LocalMux
    port map (
            O => \N__54675\,
            I => \N__54672\
        );

    \I__12698\ : Span4Mux_h
    port map (
            O => \N__54672\,
            I => \N__54669\
        );

    \I__12697\ : Span4Mux_v
    port map (
            O => \N__54669\,
            I => \N__54666\
        );

    \I__12696\ : Odrv4
    port map (
            O => \N__54666\,
            I => \pid_side.error_p_regZ0Z_19\
        );

    \I__12695\ : InMux
    port map (
            O => \N__54663\,
            I => \N__54660\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__54660\,
            I => \pid_side.O_2_16\
        );

    \I__12693\ : CascadeMux
    port map (
            O => \N__54657\,
            I => \N__54653\
        );

    \I__12692\ : CascadeMux
    port map (
            O => \N__54656\,
            I => \N__54650\
        );

    \I__12691\ : InMux
    port map (
            O => \N__54653\,
            I => \N__54642\
        );

    \I__12690\ : InMux
    port map (
            O => \N__54650\,
            I => \N__54642\
        );

    \I__12689\ : InMux
    port map (
            O => \N__54649\,
            I => \N__54642\
        );

    \I__12688\ : LocalMux
    port map (
            O => \N__54642\,
            I => \N__54639\
        );

    \I__12687\ : Span4Mux_h
    port map (
            O => \N__54639\,
            I => \N__54636\
        );

    \I__12686\ : Odrv4
    port map (
            O => \N__54636\,
            I => \pid_side.error_p_regZ0Z_12\
        );

    \I__12685\ : InMux
    port map (
            O => \N__54633\,
            I => \N__54630\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__54630\,
            I => \N__54626\
        );

    \I__12683\ : InMux
    port map (
            O => \N__54629\,
            I => \N__54623\
        );

    \I__12682\ : Span4Mux_v
    port map (
            O => \N__54626\,
            I => \N__54620\
        );

    \I__12681\ : LocalMux
    port map (
            O => \N__54623\,
            I => \pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6\
        );

    \I__12680\ : Odrv4
    port map (
            O => \N__54620\,
            I => \pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6\
        );

    \I__12679\ : CascadeMux
    port map (
            O => \N__54615\,
            I => \pid_side.un1_pid_prereg_60_0_cascade_\
        );

    \I__12678\ : CascadeMux
    port map (
            O => \N__54612\,
            I => \N__54609\
        );

    \I__12677\ : InMux
    port map (
            O => \N__54609\,
            I => \N__54606\
        );

    \I__12676\ : LocalMux
    port map (
            O => \N__54606\,
            I => \N__54603\
        );

    \I__12675\ : Span4Mux_h
    port map (
            O => \N__54603\,
            I => \N__54600\
        );

    \I__12674\ : Span4Mux_s1_h
    port map (
            O => \N__54600\,
            I => \N__54597\
        );

    \I__12673\ : Odrv4
    port map (
            O => \N__54597\,
            I => \pid_side.error_p_reg_esr_RNI1DBR2Z0Z_6\
        );

    \I__12672\ : CascadeMux
    port map (
            O => \N__54594\,
            I => \pid_side.N_1570_i_cascade_\
        );

    \I__12671\ : CascadeMux
    port map (
            O => \N__54591\,
            I => \N__54588\
        );

    \I__12670\ : InMux
    port map (
            O => \N__54588\,
            I => \N__54585\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__54585\,
            I => \N__54582\
        );

    \I__12668\ : Span4Mux_h
    port map (
            O => \N__54582\,
            I => \N__54579\
        );

    \I__12667\ : Odrv4
    port map (
            O => \N__54579\,
            I => \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7\
        );

    \I__12666\ : InMux
    port map (
            O => \N__54576\,
            I => \N__54573\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__54573\,
            I => \pid_side.un1_pid_prereg_70_0\
        );

    \I__12664\ : InMux
    port map (
            O => \N__54570\,
            I => \N__54564\
        );

    \I__12663\ : InMux
    port map (
            O => \N__54569\,
            I => \N__54557\
        );

    \I__12662\ : InMux
    port map (
            O => \N__54568\,
            I => \N__54557\
        );

    \I__12661\ : InMux
    port map (
            O => \N__54567\,
            I => \N__54557\
        );

    \I__12660\ : LocalMux
    port map (
            O => \N__54564\,
            I => \pid_side.error_p_regZ0Z_7\
        );

    \I__12659\ : LocalMux
    port map (
            O => \N__54557\,
            I => \pid_side.error_p_regZ0Z_7\
        );

    \I__12658\ : CascadeMux
    port map (
            O => \N__54552\,
            I => \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7_cascade_\
        );

    \I__12657\ : InMux
    port map (
            O => \N__54549\,
            I => \N__54546\
        );

    \I__12656\ : LocalMux
    port map (
            O => \N__54546\,
            I => \N__54543\
        );

    \I__12655\ : Span4Mux_v
    port map (
            O => \N__54543\,
            I => \N__54540\
        );

    \I__12654\ : Odrv4
    port map (
            O => \N__54540\,
            I => \pid_side.O_1_6\
        );

    \I__12653\ : InMux
    port map (
            O => \N__54537\,
            I => \N__54532\
        );

    \I__12652\ : InMux
    port map (
            O => \N__54536\,
            I => \N__54527\
        );

    \I__12651\ : InMux
    port map (
            O => \N__54535\,
            I => \N__54527\
        );

    \I__12650\ : LocalMux
    port map (
            O => \N__54532\,
            I => \pid_side.error_d_regZ0Z_2\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__54527\,
            I => \pid_side.error_d_regZ0Z_2\
        );

    \I__12648\ : InMux
    port map (
            O => \N__54522\,
            I => \N__54519\
        );

    \I__12647\ : LocalMux
    port map (
            O => \N__54519\,
            I => \N__54516\
        );

    \I__12646\ : Odrv4
    port map (
            O => \N__54516\,
            I => \pid_side.O_2_17\
        );

    \I__12645\ : InMux
    port map (
            O => \N__54513\,
            I => \N__54507\
        );

    \I__12644\ : InMux
    port map (
            O => \N__54512\,
            I => \N__54507\
        );

    \I__12643\ : LocalMux
    port map (
            O => \N__54507\,
            I => \N__54504\
        );

    \I__12642\ : Odrv4
    port map (
            O => \N__54504\,
            I => \pid_side.error_p_regZ0Z_13\
        );

    \I__12641\ : InMux
    port map (
            O => \N__54501\,
            I => \N__54498\
        );

    \I__12640\ : LocalMux
    port map (
            O => \N__54498\,
            I => \pid_side.O_2_12\
        );

    \I__12639\ : CascadeMux
    port map (
            O => \N__54495\,
            I => \N__54490\
        );

    \I__12638\ : InMux
    port map (
            O => \N__54494\,
            I => \N__54482\
        );

    \I__12637\ : InMux
    port map (
            O => \N__54493\,
            I => \N__54482\
        );

    \I__12636\ : InMux
    port map (
            O => \N__54490\,
            I => \N__54482\
        );

    \I__12635\ : InMux
    port map (
            O => \N__54489\,
            I => \N__54479\
        );

    \I__12634\ : LocalMux
    port map (
            O => \N__54482\,
            I => \N__54476\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__54479\,
            I => \pid_side.error_p_regZ0Z_8\
        );

    \I__12632\ : Odrv4
    port map (
            O => \N__54476\,
            I => \pid_side.error_p_regZ0Z_8\
        );

    \I__12631\ : InMux
    port map (
            O => \N__54471\,
            I => \N__54468\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__54468\,
            I => \N__54465\
        );

    \I__12629\ : Odrv4
    port map (
            O => \N__54465\,
            I => \pid_side.O_2_24\
        );

    \I__12628\ : InMux
    port map (
            O => \N__54462\,
            I => \N__54459\
        );

    \I__12627\ : LocalMux
    port map (
            O => \N__54459\,
            I => \N__54455\
        );

    \I__12626\ : InMux
    port map (
            O => \N__54458\,
            I => \N__54452\
        );

    \I__12625\ : Span4Mux_v
    port map (
            O => \N__54455\,
            I => \N__54447\
        );

    \I__12624\ : LocalMux
    port map (
            O => \N__54452\,
            I => \N__54447\
        );

    \I__12623\ : Sp12to4
    port map (
            O => \N__54447\,
            I => \N__54444\
        );

    \I__12622\ : Odrv12
    port map (
            O => \N__54444\,
            I => \pid_side.error_p_regZ0Z_20\
        );

    \I__12621\ : InMux
    port map (
            O => \N__54441\,
            I => \N__54438\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__54438\,
            I => \N__54435\
        );

    \I__12619\ : Odrv4
    port map (
            O => \N__54435\,
            I => \pid_side.O_2_18\
        );

    \I__12618\ : InMux
    port map (
            O => \N__54432\,
            I => \N__54428\
        );

    \I__12617\ : InMux
    port map (
            O => \N__54431\,
            I => \N__54425\
        );

    \I__12616\ : LocalMux
    port map (
            O => \N__54428\,
            I => \N__54422\
        );

    \I__12615\ : LocalMux
    port map (
            O => \N__54425\,
            I => \N__54419\
        );

    \I__12614\ : Span4Mux_h
    port map (
            O => \N__54422\,
            I => \N__54416\
        );

    \I__12613\ : Odrv12
    port map (
            O => \N__54419\,
            I => \pid_side.error_p_regZ0Z_14\
        );

    \I__12612\ : Odrv4
    port map (
            O => \N__54416\,
            I => \pid_side.error_p_regZ0Z_14\
        );

    \I__12611\ : InMux
    port map (
            O => \N__54411\,
            I => \N__54408\
        );

    \I__12610\ : LocalMux
    port map (
            O => \N__54408\,
            I => \pid_side.O_2_14\
        );

    \I__12609\ : InMux
    port map (
            O => \N__54405\,
            I => \N__54402\
        );

    \I__12608\ : LocalMux
    port map (
            O => \N__54402\,
            I => \N__54398\
        );

    \I__12607\ : InMux
    port map (
            O => \N__54401\,
            I => \N__54395\
        );

    \I__12606\ : Span4Mux_h
    port map (
            O => \N__54398\,
            I => \N__54392\
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__54395\,
            I => \N__54389\
        );

    \I__12604\ : Odrv4
    port map (
            O => \N__54392\,
            I => \pid_side.error_p_regZ0Z_10\
        );

    \I__12603\ : Odrv12
    port map (
            O => \N__54389\,
            I => \pid_side.error_p_regZ0Z_10\
        );

    \I__12602\ : InMux
    port map (
            O => \N__54384\,
            I => \N__54381\
        );

    \I__12601\ : LocalMux
    port map (
            O => \N__54381\,
            I => \pid_side.O_2_19\
        );

    \I__12600\ : InMux
    port map (
            O => \N__54378\,
            I => \N__54374\
        );

    \I__12599\ : InMux
    port map (
            O => \N__54377\,
            I => \N__54371\
        );

    \I__12598\ : LocalMux
    port map (
            O => \N__54374\,
            I => \N__54366\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__54371\,
            I => \N__54366\
        );

    \I__12596\ : Span4Mux_h
    port map (
            O => \N__54366\,
            I => \N__54363\
        );

    \I__12595\ : Odrv4
    port map (
            O => \N__54363\,
            I => \pid_side.error_p_regZ0Z_15\
        );

    \I__12594\ : InMux
    port map (
            O => \N__54360\,
            I => \N__54357\
        );

    \I__12593\ : LocalMux
    port map (
            O => \N__54357\,
            I => \pid_side.O_2_10\
        );

    \I__12592\ : InMux
    port map (
            O => \N__54354\,
            I => \N__54351\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__54351\,
            I => \pid_side.O_2_13\
        );

    \I__12590\ : InMux
    port map (
            O => \N__54348\,
            I => \N__54343\
        );

    \I__12589\ : InMux
    port map (
            O => \N__54347\,
            I => \N__54340\
        );

    \I__12588\ : InMux
    port map (
            O => \N__54346\,
            I => \N__54337\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__54343\,
            I => \N__54334\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__54340\,
            I => \pid_side.error_p_regZ0Z_9\
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__54337\,
            I => \pid_side.error_p_regZ0Z_9\
        );

    \I__12584\ : Odrv4
    port map (
            O => \N__54334\,
            I => \pid_side.error_p_regZ0Z_9\
        );

    \I__12583\ : InMux
    port map (
            O => \N__54327\,
            I => \N__54324\
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__54324\,
            I => \N__54321\
        );

    \I__12581\ : Span4Mux_h
    port map (
            O => \N__54321\,
            I => \N__54318\
        );

    \I__12580\ : Odrv4
    port map (
            O => \N__54318\,
            I => \pid_front.O_14\
        );

    \I__12579\ : InMux
    port map (
            O => \N__54315\,
            I => \N__54309\
        );

    \I__12578\ : InMux
    port map (
            O => \N__54314\,
            I => \N__54309\
        );

    \I__12577\ : LocalMux
    port map (
            O => \N__54309\,
            I => \N__54305\
        );

    \I__12576\ : InMux
    port map (
            O => \N__54308\,
            I => \N__54302\
        );

    \I__12575\ : Span4Mux_h
    port map (
            O => \N__54305\,
            I => \N__54297\
        );

    \I__12574\ : LocalMux
    port map (
            O => \N__54302\,
            I => \N__54297\
        );

    \I__12573\ : Sp12to4
    port map (
            O => \N__54297\,
            I => \N__54294\
        );

    \I__12572\ : Span12Mux_s7_v
    port map (
            O => \N__54294\,
            I => \N__54291\
        );

    \I__12571\ : Odrv12
    port map (
            O => \N__54291\,
            I => \pid_front.error_d_regZ0Z_10\
        );

    \I__12570\ : InMux
    port map (
            O => \N__54288\,
            I => \N__54285\
        );

    \I__12569\ : LocalMux
    port map (
            O => \N__54285\,
            I => \N__54282\
        );

    \I__12568\ : Odrv4
    port map (
            O => \N__54282\,
            I => \pid_side.O_2_8\
        );

    \I__12567\ : InMux
    port map (
            O => \N__54279\,
            I => \N__54273\
        );

    \I__12566\ : InMux
    port map (
            O => \N__54278\,
            I => \N__54273\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__54273\,
            I => \N__54270\
        );

    \I__12564\ : Odrv4
    port map (
            O => \N__54270\,
            I => \pid_side.error_p_regZ0Z_4\
        );

    \I__12563\ : InMux
    port map (
            O => \N__54267\,
            I => \N__54264\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__54264\,
            I => \pid_side.O_2_5\
        );

    \I__12561\ : CascadeMux
    port map (
            O => \N__54261\,
            I => \N__54258\
        );

    \I__12560\ : InMux
    port map (
            O => \N__54258\,
            I => \N__54252\
        );

    \I__12559\ : InMux
    port map (
            O => \N__54257\,
            I => \N__54252\
        );

    \I__12558\ : LocalMux
    port map (
            O => \N__54252\,
            I => \N__54249\
        );

    \I__12557\ : Odrv4
    port map (
            O => \N__54249\,
            I => \pid_side.error_p_regZ0Z_1\
        );

    \I__12556\ : InMux
    port map (
            O => \N__54246\,
            I => \N__54243\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__54243\,
            I => \pid_side.O_2_7\
        );

    \I__12554\ : InMux
    port map (
            O => \N__54240\,
            I => \N__54234\
        );

    \I__12553\ : InMux
    port map (
            O => \N__54239\,
            I => \N__54234\
        );

    \I__12552\ : LocalMux
    port map (
            O => \N__54234\,
            I => \pid_side.error_p_regZ0Z_3\
        );

    \I__12551\ : InMux
    port map (
            O => \N__54231\,
            I => \N__54228\
        );

    \I__12550\ : LocalMux
    port map (
            O => \N__54228\,
            I => \N__54225\
        );

    \I__12549\ : Span4Mux_h
    port map (
            O => \N__54225\,
            I => \N__54222\
        );

    \I__12548\ : Odrv4
    port map (
            O => \N__54222\,
            I => \pid_side.O_2_22\
        );

    \I__12547\ : InMux
    port map (
            O => \N__54219\,
            I => \N__54213\
        );

    \I__12546\ : InMux
    port map (
            O => \N__54218\,
            I => \N__54213\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__54213\,
            I => \N__54210\
        );

    \I__12544\ : Span4Mux_v
    port map (
            O => \N__54210\,
            I => \N__54207\
        );

    \I__12543\ : Odrv4
    port map (
            O => \N__54207\,
            I => \pid_side.error_p_regZ0Z_18\
        );

    \I__12542\ : InMux
    port map (
            O => \N__54204\,
            I => \N__54201\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__54201\,
            I => \pid_side.O_2_6\
        );

    \I__12540\ : InMux
    port map (
            O => \N__54198\,
            I => \N__54192\
        );

    \I__12539\ : InMux
    port map (
            O => \N__54197\,
            I => \N__54192\
        );

    \I__12538\ : LocalMux
    port map (
            O => \N__54192\,
            I => \pid_side.error_p_regZ0Z_2\
        );

    \I__12537\ : InMux
    port map (
            O => \N__54189\,
            I => \N__54186\
        );

    \I__12536\ : LocalMux
    port map (
            O => \N__54186\,
            I => \N__54183\
        );

    \I__12535\ : Odrv4
    port map (
            O => \N__54183\,
            I => \pid_side.O_2_20\
        );

    \I__12534\ : InMux
    port map (
            O => \N__54180\,
            I => \N__54174\
        );

    \I__12533\ : InMux
    port map (
            O => \N__54179\,
            I => \N__54174\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__54174\,
            I => \N__54171\
        );

    \I__12531\ : Span4Mux_v
    port map (
            O => \N__54171\,
            I => \N__54168\
        );

    \I__12530\ : Span4Mux_h
    port map (
            O => \N__54168\,
            I => \N__54165\
        );

    \I__12529\ : Odrv4
    port map (
            O => \N__54165\,
            I => \pid_side.error_p_regZ0Z_16\
        );

    \I__12528\ : InMux
    port map (
            O => \N__54162\,
            I => \N__54159\
        );

    \I__12527\ : LocalMux
    port map (
            O => \N__54159\,
            I => \N__54156\
        );

    \I__12526\ : Odrv4
    port map (
            O => \N__54156\,
            I => \pid_side.O_2_21\
        );

    \I__12525\ : InMux
    port map (
            O => \N__54153\,
            I => \N__54147\
        );

    \I__12524\ : InMux
    port map (
            O => \N__54152\,
            I => \N__54147\
        );

    \I__12523\ : LocalMux
    port map (
            O => \N__54147\,
            I => \N__54144\
        );

    \I__12522\ : Odrv4
    port map (
            O => \N__54144\,
            I => \pid_side.error_p_regZ0Z_17\
        );

    \I__12521\ : InMux
    port map (
            O => \N__54141\,
            I => \N__54136\
        );

    \I__12520\ : InMux
    port map (
            O => \N__54140\,
            I => \N__54133\
        );

    \I__12519\ : InMux
    port map (
            O => \N__54139\,
            I => \N__54130\
        );

    \I__12518\ : LocalMux
    port map (
            O => \N__54136\,
            I => \pid_side.error_d_reg_prevZ0Z_9\
        );

    \I__12517\ : LocalMux
    port map (
            O => \N__54133\,
            I => \pid_side.error_d_reg_prevZ0Z_9\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__54130\,
            I => \pid_side.error_d_reg_prevZ0Z_9\
        );

    \I__12515\ : CascadeMux
    port map (
            O => \N__54123\,
            I => \N__54118\
        );

    \I__12514\ : InMux
    port map (
            O => \N__54122\,
            I => \N__54113\
        );

    \I__12513\ : InMux
    port map (
            O => \N__54121\,
            I => \N__54113\
        );

    \I__12512\ : InMux
    port map (
            O => \N__54118\,
            I => \N__54110\
        );

    \I__12511\ : LocalMux
    port map (
            O => \N__54113\,
            I => \N__54107\
        );

    \I__12510\ : LocalMux
    port map (
            O => \N__54110\,
            I => \pid_side.un1_pid_prereg_41\
        );

    \I__12509\ : Odrv4
    port map (
            O => \N__54107\,
            I => \pid_side.un1_pid_prereg_41\
        );

    \I__12508\ : InMux
    port map (
            O => \N__54102\,
            I => \N__54099\
        );

    \I__12507\ : LocalMux
    port map (
            O => \N__54099\,
            I => \N__54096\
        );

    \I__12506\ : Span4Mux_v
    port map (
            O => \N__54096\,
            I => \N__54091\
        );

    \I__12505\ : InMux
    port map (
            O => \N__54095\,
            I => \N__54086\
        );

    \I__12504\ : InMux
    port map (
            O => \N__54094\,
            I => \N__54086\
        );

    \I__12503\ : Odrv4
    port map (
            O => \N__54091\,
            I => \pid_side.un1_pid_prereg_42\
        );

    \I__12502\ : LocalMux
    port map (
            O => \N__54086\,
            I => \pid_side.un1_pid_prereg_42\
        );

    \I__12501\ : CascadeMux
    port map (
            O => \N__54081\,
            I => \N__54078\
        );

    \I__12500\ : InMux
    port map (
            O => \N__54078\,
            I => \N__54072\
        );

    \I__12499\ : InMux
    port map (
            O => \N__54077\,
            I => \N__54072\
        );

    \I__12498\ : LocalMux
    port map (
            O => \N__54072\,
            I => \pid_side.error_d_reg_prevZ0Z_17\
        );

    \I__12497\ : InMux
    port map (
            O => \N__54069\,
            I => \N__54066\
        );

    \I__12496\ : LocalMux
    port map (
            O => \N__54066\,
            I => \N__54063\
        );

    \I__12495\ : Span4Mux_h
    port map (
            O => \N__54063\,
            I => \N__54060\
        );

    \I__12494\ : Odrv4
    port map (
            O => \N__54060\,
            I => \pid_side.O_1_13\
        );

    \I__12493\ : InMux
    port map (
            O => \N__54057\,
            I => \N__54054\
        );

    \I__12492\ : LocalMux
    port map (
            O => \N__54054\,
            I => \N__54049\
        );

    \I__12491\ : InMux
    port map (
            O => \N__54053\,
            I => \N__54044\
        );

    \I__12490\ : InMux
    port map (
            O => \N__54052\,
            I => \N__54044\
        );

    \I__12489\ : Sp12to4
    port map (
            O => \N__54049\,
            I => \N__54039\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__54044\,
            I => \N__54039\
        );

    \I__12487\ : Odrv12
    port map (
            O => \N__54039\,
            I => \pid_side.error_d_regZ0Z_9\
        );

    \I__12486\ : CascadeMux
    port map (
            O => \N__54036\,
            I => \N__54031\
        );

    \I__12485\ : CascadeMux
    port map (
            O => \N__54035\,
            I => \N__54025\
        );

    \I__12484\ : InMux
    port map (
            O => \N__54034\,
            I => \N__54022\
        );

    \I__12483\ : InMux
    port map (
            O => \N__54031\,
            I => \N__54015\
        );

    \I__12482\ : InMux
    port map (
            O => \N__54030\,
            I => \N__54015\
        );

    \I__12481\ : InMux
    port map (
            O => \N__54029\,
            I => \N__54015\
        );

    \I__12480\ : InMux
    port map (
            O => \N__54028\,
            I => \N__54010\
        );

    \I__12479\ : InMux
    port map (
            O => \N__54025\,
            I => \N__54010\
        );

    \I__12478\ : LocalMux
    port map (
            O => \N__54022\,
            I => \N__54007\
        );

    \I__12477\ : LocalMux
    port map (
            O => \N__54015\,
            I => \N__54002\
        );

    \I__12476\ : LocalMux
    port map (
            O => \N__54010\,
            I => \N__54002\
        );

    \I__12475\ : Span4Mux_h
    port map (
            O => \N__54007\,
            I => \N__53999\
        );

    \I__12474\ : Span4Mux_h
    port map (
            O => \N__54002\,
            I => \N__53996\
        );

    \I__12473\ : Odrv4
    port map (
            O => \N__53999\,
            I => \pid_side.un1_pid_prereg_93\
        );

    \I__12472\ : Odrv4
    port map (
            O => \N__53996\,
            I => \pid_side.un1_pid_prereg_93\
        );

    \I__12471\ : CascadeMux
    port map (
            O => \N__53991\,
            I => \N__53987\
        );

    \I__12470\ : InMux
    port map (
            O => \N__53990\,
            I => \N__53984\
        );

    \I__12469\ : InMux
    port map (
            O => \N__53987\,
            I => \N__53975\
        );

    \I__12468\ : LocalMux
    port map (
            O => \N__53984\,
            I => \N__53971\
        );

    \I__12467\ : InMux
    port map (
            O => \N__53983\,
            I => \N__53962\
        );

    \I__12466\ : InMux
    port map (
            O => \N__53982\,
            I => \N__53962\
        );

    \I__12465\ : InMux
    port map (
            O => \N__53981\,
            I => \N__53962\
        );

    \I__12464\ : InMux
    port map (
            O => \N__53980\,
            I => \N__53962\
        );

    \I__12463\ : InMux
    port map (
            O => \N__53979\,
            I => \N__53957\
        );

    \I__12462\ : InMux
    port map (
            O => \N__53978\,
            I => \N__53957\
        );

    \I__12461\ : LocalMux
    port map (
            O => \N__53975\,
            I => \N__53954\
        );

    \I__12460\ : InMux
    port map (
            O => \N__53974\,
            I => \N__53951\
        );

    \I__12459\ : Span4Mux_h
    port map (
            O => \N__53971\,
            I => \N__53948\
        );

    \I__12458\ : LocalMux
    port map (
            O => \N__53962\,
            I => \N__53939\
        );

    \I__12457\ : LocalMux
    port map (
            O => \N__53957\,
            I => \N__53939\
        );

    \I__12456\ : Span4Mux_v
    port map (
            O => \N__53954\,
            I => \N__53939\
        );

    \I__12455\ : LocalMux
    port map (
            O => \N__53951\,
            I => \N__53939\
        );

    \I__12454\ : Span4Mux_v
    port map (
            O => \N__53948\,
            I => \N__53936\
        );

    \I__12453\ : Span4Mux_v
    port map (
            O => \N__53939\,
            I => \N__53933\
        );

    \I__12452\ : Odrv4
    port map (
            O => \N__53936\,
            I => \pid_side.un1_pid_prereg_92\
        );

    \I__12451\ : Odrv4
    port map (
            O => \N__53933\,
            I => \pid_side.un1_pid_prereg_92\
        );

    \I__12450\ : InMux
    port map (
            O => \N__53928\,
            I => \N__53925\
        );

    \I__12449\ : LocalMux
    port map (
            O => \N__53925\,
            I => \N__53922\
        );

    \I__12448\ : Span4Mux_h
    port map (
            O => \N__53922\,
            I => \N__53919\
        );

    \I__12447\ : Odrv4
    port map (
            O => \N__53919\,
            I => \pid_front.O_12\
        );

    \I__12446\ : CascadeMux
    port map (
            O => \N__53916\,
            I => \N__53912\
        );

    \I__12445\ : InMux
    port map (
            O => \N__53915\,
            I => \N__53908\
        );

    \I__12444\ : InMux
    port map (
            O => \N__53912\,
            I => \N__53905\
        );

    \I__12443\ : InMux
    port map (
            O => \N__53911\,
            I => \N__53902\
        );

    \I__12442\ : LocalMux
    port map (
            O => \N__53908\,
            I => \N__53899\
        );

    \I__12441\ : LocalMux
    port map (
            O => \N__53905\,
            I => \N__53894\
        );

    \I__12440\ : LocalMux
    port map (
            O => \N__53902\,
            I => \N__53894\
        );

    \I__12439\ : Span4Mux_v
    port map (
            O => \N__53899\,
            I => \N__53891\
        );

    \I__12438\ : Span4Mux_h
    port map (
            O => \N__53894\,
            I => \N__53888\
        );

    \I__12437\ : Span4Mux_h
    port map (
            O => \N__53891\,
            I => \N__53885\
        );

    \I__12436\ : Span4Mux_h
    port map (
            O => \N__53888\,
            I => \N__53882\
        );

    \I__12435\ : Sp12to4
    port map (
            O => \N__53885\,
            I => \N__53879\
        );

    \I__12434\ : Span4Mux_h
    port map (
            O => \N__53882\,
            I => \N__53876\
        );

    \I__12433\ : Span12Mux_h
    port map (
            O => \N__53879\,
            I => \N__53873\
        );

    \I__12432\ : Span4Mux_h
    port map (
            O => \N__53876\,
            I => \N__53870\
        );

    \I__12431\ : Odrv12
    port map (
            O => \N__53873\,
            I => \pid_front.error_d_regZ0Z_8\
        );

    \I__12430\ : Odrv4
    port map (
            O => \N__53870\,
            I => \pid_front.error_d_regZ0Z_8\
        );

    \I__12429\ : InMux
    port map (
            O => \N__53865\,
            I => \N__53862\
        );

    \I__12428\ : LocalMux
    port map (
            O => \N__53862\,
            I => \N__53859\
        );

    \I__12427\ : Span4Mux_h
    port map (
            O => \N__53859\,
            I => \N__53856\
        );

    \I__12426\ : Odrv4
    port map (
            O => \N__53856\,
            I => \pid_front.O_16\
        );

    \I__12425\ : InMux
    port map (
            O => \N__53853\,
            I => \N__53850\
        );

    \I__12424\ : LocalMux
    port map (
            O => \N__53850\,
            I => \N__53845\
        );

    \I__12423\ : InMux
    port map (
            O => \N__53849\,
            I => \N__53840\
        );

    \I__12422\ : InMux
    port map (
            O => \N__53848\,
            I => \N__53840\
        );

    \I__12421\ : Span4Mux_h
    port map (
            O => \N__53845\,
            I => \N__53835\
        );

    \I__12420\ : LocalMux
    port map (
            O => \N__53840\,
            I => \N__53835\
        );

    \I__12419\ : Sp12to4
    port map (
            O => \N__53835\,
            I => \N__53832\
        );

    \I__12418\ : Span12Mux_s7_v
    port map (
            O => \N__53832\,
            I => \N__53829\
        );

    \I__12417\ : Span12Mux_h
    port map (
            O => \N__53829\,
            I => \N__53826\
        );

    \I__12416\ : Odrv12
    port map (
            O => \N__53826\,
            I => \pid_front.error_d_regZ0Z_12\
        );

    \I__12415\ : CascadeMux
    port map (
            O => \N__53823\,
            I => \N__53820\
        );

    \I__12414\ : InMux
    port map (
            O => \N__53820\,
            I => \N__53816\
        );

    \I__12413\ : InMux
    port map (
            O => \N__53819\,
            I => \N__53811\
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__53816\,
            I => \N__53808\
        );

    \I__12411\ : InMux
    port map (
            O => \N__53815\,
            I => \N__53803\
        );

    \I__12410\ : InMux
    port map (
            O => \N__53814\,
            I => \N__53803\
        );

    \I__12409\ : LocalMux
    port map (
            O => \N__53811\,
            I => \pid_side.error_p_regZ0Z_5\
        );

    \I__12408\ : Odrv4
    port map (
            O => \N__53808\,
            I => \pid_side.error_p_regZ0Z_5\
        );

    \I__12407\ : LocalMux
    port map (
            O => \N__53803\,
            I => \pid_side.error_p_regZ0Z_5\
        );

    \I__12406\ : InMux
    port map (
            O => \N__53796\,
            I => \N__53792\
        );

    \I__12405\ : CascadeMux
    port map (
            O => \N__53795\,
            I => \N__53789\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__53792\,
            I => \N__53785\
        );

    \I__12403\ : InMux
    port map (
            O => \N__53789\,
            I => \N__53779\
        );

    \I__12402\ : InMux
    port map (
            O => \N__53788\,
            I => \N__53779\
        );

    \I__12401\ : Span4Mux_v
    port map (
            O => \N__53785\,
            I => \N__53776\
        );

    \I__12400\ : InMux
    port map (
            O => \N__53784\,
            I => \N__53773\
        );

    \I__12399\ : LocalMux
    port map (
            O => \N__53779\,
            I => \N__53770\
        );

    \I__12398\ : Odrv4
    port map (
            O => \N__53776\,
            I => \pid_side.error_d_reg_prevZ0Z_5\
        );

    \I__12397\ : LocalMux
    port map (
            O => \N__53773\,
            I => \pid_side.error_d_reg_prevZ0Z_5\
        );

    \I__12396\ : Odrv4
    port map (
            O => \N__53770\,
            I => \pid_side.error_d_reg_prevZ0Z_5\
        );

    \I__12395\ : CascadeMux
    port map (
            O => \N__53763\,
            I => \pid_side.N_1566_i_cascade_\
        );

    \I__12394\ : CascadeMux
    port map (
            O => \N__53760\,
            I => \pid_side.N_1578_i_cascade_\
        );

    \I__12393\ : CascadeMux
    port map (
            O => \N__53757\,
            I => \N__53753\
        );

    \I__12392\ : CascadeMux
    port map (
            O => \N__53756\,
            I => \N__53750\
        );

    \I__12391\ : InMux
    port map (
            O => \N__53753\,
            I => \N__53747\
        );

    \I__12390\ : InMux
    port map (
            O => \N__53750\,
            I => \N__53744\
        );

    \I__12389\ : LocalMux
    port map (
            O => \N__53747\,
            I => \N__53741\
        );

    \I__12388\ : LocalMux
    port map (
            O => \N__53744\,
            I => \N__53738\
        );

    \I__12387\ : Span4Mux_h
    port map (
            O => \N__53741\,
            I => \N__53735\
        );

    \I__12386\ : Odrv4
    port map (
            O => \N__53738\,
            I => \pid_side.error_d_reg_esr_RNID3MD1Z0Z_9\
        );

    \I__12385\ : Odrv4
    port map (
            O => \N__53735\,
            I => \pid_side.error_d_reg_esr_RNID3MD1Z0Z_9\
        );

    \I__12384\ : CascadeMux
    port map (
            O => \N__53730\,
            I => \pid_side.N_1574_i_cascade_\
        );

    \I__12383\ : CascadeMux
    port map (
            O => \N__53727\,
            I => \N__53724\
        );

    \I__12382\ : InMux
    port map (
            O => \N__53724\,
            I => \N__53721\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__53721\,
            I => \N__53718\
        );

    \I__12380\ : Span4Mux_v
    port map (
            O => \N__53718\,
            I => \N__53715\
        );

    \I__12379\ : Odrv4
    port map (
            O => \N__53715\,
            I => \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8\
        );

    \I__12378\ : InMux
    port map (
            O => \N__53712\,
            I => \N__53709\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__53709\,
            I => \pid_side.un1_pid_prereg_80_0\
        );

    \I__12376\ : CascadeMux
    port map (
            O => \N__53706\,
            I => \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8_cascade_\
        );

    \I__12375\ : InMux
    port map (
            O => \N__53703\,
            I => \N__53700\
        );

    \I__12374\ : LocalMux
    port map (
            O => \N__53700\,
            I => \N__53697\
        );

    \I__12373\ : Span4Mux_h
    port map (
            O => \N__53697\,
            I => \N__53694\
        );

    \I__12372\ : Odrv4
    port map (
            O => \N__53694\,
            I => \pid_side.error_p_reg_esr_RNIL1CR2Z0Z_8\
        );

    \I__12371\ : InMux
    port map (
            O => \N__53691\,
            I => \N__53685\
        );

    \I__12370\ : InMux
    port map (
            O => \N__53690\,
            I => \N__53678\
        );

    \I__12369\ : InMux
    port map (
            O => \N__53689\,
            I => \N__53678\
        );

    \I__12368\ : InMux
    port map (
            O => \N__53688\,
            I => \N__53678\
        );

    \I__12367\ : LocalMux
    port map (
            O => \N__53685\,
            I => \pid_side.error_d_reg_prevZ0Z_8\
        );

    \I__12366\ : LocalMux
    port map (
            O => \N__53678\,
            I => \pid_side.error_d_reg_prevZ0Z_8\
        );

    \I__12365\ : CascadeMux
    port map (
            O => \N__53673\,
            I => \N__53669\
        );

    \I__12364\ : InMux
    port map (
            O => \N__53672\,
            I => \N__53666\
        );

    \I__12363\ : InMux
    port map (
            O => \N__53669\,
            I => \N__53663\
        );

    \I__12362\ : LocalMux
    port map (
            O => \N__53666\,
            I => \pid_side.un1_pid_prereg_2\
        );

    \I__12361\ : LocalMux
    port map (
            O => \N__53663\,
            I => \pid_side.un1_pid_prereg_2\
        );

    \I__12360\ : CascadeMux
    port map (
            O => \N__53658\,
            I => \pid_side.un1_pid_prereg_2_cascade_\
        );

    \I__12359\ : InMux
    port map (
            O => \N__53655\,
            I => \N__53652\
        );

    \I__12358\ : LocalMux
    port map (
            O => \N__53652\,
            I => \N__53649\
        );

    \I__12357\ : Odrv4
    port map (
            O => \N__53649\,
            I => \pid_side.error_p_reg_esr_RNIRPSK1Z0Z_2\
        );

    \I__12356\ : InMux
    port map (
            O => \N__53646\,
            I => \N__53639\
        );

    \I__12355\ : InMux
    port map (
            O => \N__53645\,
            I => \N__53639\
        );

    \I__12354\ : InMux
    port map (
            O => \N__53644\,
            I => \N__53636\
        );

    \I__12353\ : LocalMux
    port map (
            O => \N__53639\,
            I => \N__53633\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__53636\,
            I => \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2\
        );

    \I__12351\ : Odrv4
    port map (
            O => \N__53633\,
            I => \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2\
        );

    \I__12350\ : CascadeMux
    port map (
            O => \N__53628\,
            I => \N__53625\
        );

    \I__12349\ : InMux
    port map (
            O => \N__53625\,
            I => \N__53620\
        );

    \I__12348\ : InMux
    port map (
            O => \N__53624\,
            I => \N__53615\
        );

    \I__12347\ : InMux
    port map (
            O => \N__53623\,
            I => \N__53615\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__53620\,
            I => \pid_side.un1_pid_prereg_0\
        );

    \I__12345\ : LocalMux
    port map (
            O => \N__53615\,
            I => \pid_side.un1_pid_prereg_0\
        );

    \I__12344\ : InMux
    port map (
            O => \N__53610\,
            I => \N__53604\
        );

    \I__12343\ : InMux
    port map (
            O => \N__53609\,
            I => \N__53604\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__53604\,
            I => \pid_side.error_d_reg_prevZ0Z_3\
        );

    \I__12341\ : InMux
    port map (
            O => \N__53601\,
            I => \N__53596\
        );

    \I__12340\ : InMux
    port map (
            O => \N__53600\,
            I => \N__53591\
        );

    \I__12339\ : InMux
    port map (
            O => \N__53599\,
            I => \N__53591\
        );

    \I__12338\ : LocalMux
    port map (
            O => \N__53596\,
            I => \pid_side.un1_pid_prereg_3\
        );

    \I__12337\ : LocalMux
    port map (
            O => \N__53591\,
            I => \pid_side.un1_pid_prereg_3\
        );

    \I__12336\ : CascadeMux
    port map (
            O => \N__53586\,
            I => \N__53583\
        );

    \I__12335\ : InMux
    port map (
            O => \N__53583\,
            I => \N__53577\
        );

    \I__12334\ : InMux
    port map (
            O => \N__53582\,
            I => \N__53577\
        );

    \I__12333\ : LocalMux
    port map (
            O => \N__53577\,
            I => \pid_side.error_d_reg_prevZ0Z_2\
        );

    \I__12332\ : InMux
    port map (
            O => \N__53574\,
            I => \N__53570\
        );

    \I__12331\ : InMux
    port map (
            O => \N__53573\,
            I => \N__53567\
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__53570\,
            I => \N__53564\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__53567\,
            I => \N__53561\
        );

    \I__12328\ : Odrv4
    port map (
            O => \N__53564\,
            I => \pid_side.error_d_reg_prevZ0Z_14\
        );

    \I__12327\ : Odrv4
    port map (
            O => \N__53561\,
            I => \pid_side.error_d_reg_prevZ0Z_14\
        );

    \I__12326\ : CascadeMux
    port map (
            O => \N__53556\,
            I => \pid_side.un1_pid_prereg_47_cascade_\
        );

    \I__12325\ : CascadeMux
    port map (
            O => \N__53553\,
            I => \N__53550\
        );

    \I__12324\ : InMux
    port map (
            O => \N__53550\,
            I => \N__53547\
        );

    \I__12323\ : LocalMux
    port map (
            O => \N__53547\,
            I => \N__53544\
        );

    \I__12322\ : Span4Mux_h
    port map (
            O => \N__53544\,
            I => \N__53541\
        );

    \I__12321\ : Odrv4
    port map (
            O => \N__53541\,
            I => \pid_side.error_d_reg_prev_esr_RNIVB6H1Z0Z_17\
        );

    \I__12320\ : InMux
    port map (
            O => \N__53538\,
            I => \N__53534\
        );

    \I__12319\ : InMux
    port map (
            O => \N__53537\,
            I => \N__53531\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__53534\,
            I => \N__53528\
        );

    \I__12317\ : LocalMux
    port map (
            O => \N__53531\,
            I => \N__53523\
        );

    \I__12316\ : Span4Mux_h
    port map (
            O => \N__53528\,
            I => \N__53523\
        );

    \I__12315\ : Odrv4
    port map (
            O => \N__53523\,
            I => \pid_side.error_d_reg_prevZ0Z_10\
        );

    \I__12314\ : InMux
    port map (
            O => \N__53520\,
            I => \N__53517\
        );

    \I__12313\ : LocalMux
    port map (
            O => \N__53517\,
            I => \N__53514\
        );

    \I__12312\ : Odrv4
    port map (
            O => \N__53514\,
            I => \pid_side.O_1_4\
        );

    \I__12311\ : CascadeMux
    port map (
            O => \N__53511\,
            I => \N__53506\
        );

    \I__12310\ : CascadeMux
    port map (
            O => \N__53510\,
            I => \N__53503\
        );

    \I__12309\ : InMux
    port map (
            O => \N__53509\,
            I => \N__53500\
        );

    \I__12308\ : InMux
    port map (
            O => \N__53506\,
            I => \N__53497\
        );

    \I__12307\ : InMux
    port map (
            O => \N__53503\,
            I => \N__53494\
        );

    \I__12306\ : LocalMux
    port map (
            O => \N__53500\,
            I => \N__53491\
        );

    \I__12305\ : LocalMux
    port map (
            O => \N__53497\,
            I => \N__53486\
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__53494\,
            I => \N__53486\
        );

    \I__12303\ : Span4Mux_h
    port map (
            O => \N__53491\,
            I => \N__53483\
        );

    \I__12302\ : Span4Mux_h
    port map (
            O => \N__53486\,
            I => \N__53480\
        );

    \I__12301\ : Span4Mux_v
    port map (
            O => \N__53483\,
            I => \N__53475\
        );

    \I__12300\ : Span4Mux_v
    port map (
            O => \N__53480\,
            I => \N__53475\
        );

    \I__12299\ : Odrv4
    port map (
            O => \N__53475\,
            I => \pid_side.error_d_regZ0Z_0\
        );

    \I__12298\ : InMux
    port map (
            O => \N__53472\,
            I => \N__53469\
        );

    \I__12297\ : LocalMux
    port map (
            O => \N__53469\,
            I => \N__53466\
        );

    \I__12296\ : Span4Mux_v
    port map (
            O => \N__53466\,
            I => \N__53463\
        );

    \I__12295\ : Odrv4
    port map (
            O => \N__53463\,
            I => \pid_side.O_1_8\
        );

    \I__12294\ : InMux
    port map (
            O => \N__53460\,
            I => \N__53451\
        );

    \I__12293\ : InMux
    port map (
            O => \N__53459\,
            I => \N__53451\
        );

    \I__12292\ : InMux
    port map (
            O => \N__53458\,
            I => \N__53451\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__53451\,
            I => \N__53448\
        );

    \I__12290\ : Odrv12
    port map (
            O => \N__53448\,
            I => \pid_side.error_d_regZ0Z_4\
        );

    \I__12289\ : InMux
    port map (
            O => \N__53445\,
            I => \N__53442\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__53442\,
            I => \N__53439\
        );

    \I__12287\ : Odrv4
    port map (
            O => \N__53439\,
            I => \pid_side.O_1_5\
        );

    \I__12286\ : InMux
    port map (
            O => \N__53436\,
            I => \N__53432\
        );

    \I__12285\ : CascadeMux
    port map (
            O => \N__53435\,
            I => \N__53428\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__53432\,
            I => \N__53425\
        );

    \I__12283\ : InMux
    port map (
            O => \N__53431\,
            I => \N__53420\
        );

    \I__12282\ : InMux
    port map (
            O => \N__53428\,
            I => \N__53420\
        );

    \I__12281\ : Span4Mux_h
    port map (
            O => \N__53425\,
            I => \N__53415\
        );

    \I__12280\ : LocalMux
    port map (
            O => \N__53420\,
            I => \N__53415\
        );

    \I__12279\ : Span4Mux_v
    port map (
            O => \N__53415\,
            I => \N__53412\
        );

    \I__12278\ : Odrv4
    port map (
            O => \N__53412\,
            I => \pid_side.error_d_regZ0Z_1\
        );

    \I__12277\ : InMux
    port map (
            O => \N__53409\,
            I => \N__53406\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__53406\,
            I => \N__53402\
        );

    \I__12275\ : CascadeMux
    port map (
            O => \N__53405\,
            I => \N__53398\
        );

    \I__12274\ : Span4Mux_v
    port map (
            O => \N__53402\,
            I => \N__53393\
        );

    \I__12273\ : InMux
    port map (
            O => \N__53401\,
            I => \N__53390\
        );

    \I__12272\ : InMux
    port map (
            O => \N__53398\,
            I => \N__53387\
        );

    \I__12271\ : InMux
    port map (
            O => \N__53397\,
            I => \N__53383\
        );

    \I__12270\ : InMux
    port map (
            O => \N__53396\,
            I => \N__53380\
        );

    \I__12269\ : Span4Mux_h
    port map (
            O => \N__53393\,
            I => \N__53376\
        );

    \I__12268\ : LocalMux
    port map (
            O => \N__53390\,
            I => \N__53371\
        );

    \I__12267\ : LocalMux
    port map (
            O => \N__53387\,
            I => \N__53371\
        );

    \I__12266\ : InMux
    port map (
            O => \N__53386\,
            I => \N__53367\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__53383\,
            I => \N__53364\
        );

    \I__12264\ : LocalMux
    port map (
            O => \N__53380\,
            I => \N__53361\
        );

    \I__12263\ : InMux
    port map (
            O => \N__53379\,
            I => \N__53357\
        );

    \I__12262\ : Span4Mux_v
    port map (
            O => \N__53376\,
            I => \N__53354\
        );

    \I__12261\ : Span4Mux_v
    port map (
            O => \N__53371\,
            I => \N__53351\
        );

    \I__12260\ : InMux
    port map (
            O => \N__53370\,
            I => \N__53346\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__53367\,
            I => \N__53343\
        );

    \I__12258\ : Span4Mux_v
    port map (
            O => \N__53364\,
            I => \N__53340\
        );

    \I__12257\ : Span4Mux_h
    port map (
            O => \N__53361\,
            I => \N__53337\
        );

    \I__12256\ : InMux
    port map (
            O => \N__53360\,
            I => \N__53334\
        );

    \I__12255\ : LocalMux
    port map (
            O => \N__53357\,
            I => \N__53331\
        );

    \I__12254\ : Span4Mux_h
    port map (
            O => \N__53354\,
            I => \N__53326\
        );

    \I__12253\ : Span4Mux_h
    port map (
            O => \N__53351\,
            I => \N__53326\
        );

    \I__12252\ : InMux
    port map (
            O => \N__53350\,
            I => \N__53321\
        );

    \I__12251\ : InMux
    port map (
            O => \N__53349\,
            I => \N__53318\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__53346\,
            I => \N__53315\
        );

    \I__12249\ : Span4Mux_v
    port map (
            O => \N__53343\,
            I => \N__53312\
        );

    \I__12248\ : Span4Mux_v
    port map (
            O => \N__53340\,
            I => \N__53309\
        );

    \I__12247\ : Sp12to4
    port map (
            O => \N__53337\,
            I => \N__53306\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__53334\,
            I => \N__53303\
        );

    \I__12245\ : Span4Mux_v
    port map (
            O => \N__53331\,
            I => \N__53300\
        );

    \I__12244\ : Span4Mux_v
    port map (
            O => \N__53326\,
            I => \N__53297\
        );

    \I__12243\ : InMux
    port map (
            O => \N__53325\,
            I => \N__53294\
        );

    \I__12242\ : InMux
    port map (
            O => \N__53324\,
            I => \N__53291\
        );

    \I__12241\ : LocalMux
    port map (
            O => \N__53321\,
            I => \N__53288\
        );

    \I__12240\ : LocalMux
    port map (
            O => \N__53318\,
            I => \N__53283\
        );

    \I__12239\ : Span4Mux_h
    port map (
            O => \N__53315\,
            I => \N__53283\
        );

    \I__12238\ : Span4Mux_h
    port map (
            O => \N__53312\,
            I => \N__53280\
        );

    \I__12237\ : Sp12to4
    port map (
            O => \N__53309\,
            I => \N__53275\
        );

    \I__12236\ : Span12Mux_v
    port map (
            O => \N__53306\,
            I => \N__53275\
        );

    \I__12235\ : Span4Mux_h
    port map (
            O => \N__53303\,
            I => \N__53266\
        );

    \I__12234\ : Span4Mux_h
    port map (
            O => \N__53300\,
            I => \N__53266\
        );

    \I__12233\ : Span4Mux_v
    port map (
            O => \N__53297\,
            I => \N__53266\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__53294\,
            I => \N__53266\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__53291\,
            I => uart_pc_data_4
        );

    \I__12230\ : Odrv12
    port map (
            O => \N__53288\,
            I => uart_pc_data_4
        );

    \I__12229\ : Odrv4
    port map (
            O => \N__53283\,
            I => uart_pc_data_4
        );

    \I__12228\ : Odrv4
    port map (
            O => \N__53280\,
            I => uart_pc_data_4
        );

    \I__12227\ : Odrv12
    port map (
            O => \N__53275\,
            I => uart_pc_data_4
        );

    \I__12226\ : Odrv4
    port map (
            O => \N__53266\,
            I => uart_pc_data_4
        );

    \I__12225\ : InMux
    port map (
            O => \N__53253\,
            I => \N__53250\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__53250\,
            I => \N__53246\
        );

    \I__12223\ : InMux
    port map (
            O => \N__53249\,
            I => \N__53243\
        );

    \I__12222\ : Span4Mux_s2_h
    port map (
            O => \N__53246\,
            I => \N__53240\
        );

    \I__12221\ : LocalMux
    port map (
            O => \N__53243\,
            I => \N__53237\
        );

    \I__12220\ : Span4Mux_v
    port map (
            O => \N__53240\,
            I => \N__53232\
        );

    \I__12219\ : Span4Mux_s2_h
    port map (
            O => \N__53237\,
            I => \N__53232\
        );

    \I__12218\ : Odrv4
    port map (
            O => \N__53232\,
            I => xy_kd_4
        );

    \I__12217\ : InMux
    port map (
            O => \N__53229\,
            I => \N__53225\
        );

    \I__12216\ : InMux
    port map (
            O => \N__53228\,
            I => \N__53221\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__53225\,
            I => \N__53218\
        );

    \I__12214\ : InMux
    port map (
            O => \N__53224\,
            I => \N__53215\
        );

    \I__12213\ : LocalMux
    port map (
            O => \N__53221\,
            I => \N__53212\
        );

    \I__12212\ : Span4Mux_h
    port map (
            O => \N__53218\,
            I => \N__53206\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__53215\,
            I => \N__53206\
        );

    \I__12210\ : Span4Mux_h
    port map (
            O => \N__53212\,
            I => \N__53201\
        );

    \I__12209\ : InMux
    port map (
            O => \N__53211\,
            I => \N__53198\
        );

    \I__12208\ : Span4Mux_v
    port map (
            O => \N__53206\,
            I => \N__53195\
        );

    \I__12207\ : InMux
    port map (
            O => \N__53205\,
            I => \N__53192\
        );

    \I__12206\ : InMux
    port map (
            O => \N__53204\,
            I => \N__53189\
        );

    \I__12205\ : Span4Mux_v
    port map (
            O => \N__53201\,
            I => \N__53186\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__53198\,
            I => \N__53181\
        );

    \I__12203\ : Span4Mux_v
    port map (
            O => \N__53195\,
            I => \N__53178\
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__53192\,
            I => \N__53173\
        );

    \I__12201\ : LocalMux
    port map (
            O => \N__53189\,
            I => \N__53173\
        );

    \I__12200\ : Span4Mux_v
    port map (
            O => \N__53186\,
            I => \N__53170\
        );

    \I__12199\ : InMux
    port map (
            O => \N__53185\,
            I => \N__53167\
        );

    \I__12198\ : InMux
    port map (
            O => \N__53184\,
            I => \N__53164\
        );

    \I__12197\ : Span12Mux_v
    port map (
            O => \N__53181\,
            I => \N__53161\
        );

    \I__12196\ : Sp12to4
    port map (
            O => \N__53178\,
            I => \N__53156\
        );

    \I__12195\ : Span12Mux_v
    port map (
            O => \N__53173\,
            I => \N__53156\
        );

    \I__12194\ : Span4Mux_v
    port map (
            O => \N__53170\,
            I => \N__53149\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__53167\,
            I => \N__53149\
        );

    \I__12192\ : LocalMux
    port map (
            O => \N__53164\,
            I => \N__53149\
        );

    \I__12191\ : Odrv12
    port map (
            O => \N__53161\,
            I => uart_drone_data_6
        );

    \I__12190\ : Odrv12
    port map (
            O => \N__53156\,
            I => uart_drone_data_6
        );

    \I__12189\ : Odrv4
    port map (
            O => \N__53149\,
            I => uart_drone_data_6
        );

    \I__12188\ : InMux
    port map (
            O => \N__53142\,
            I => \N__53136\
        );

    \I__12187\ : InMux
    port map (
            O => \N__53141\,
            I => \N__53136\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__53136\,
            I => \drone_H_disp_side_14\
        );

    \I__12185\ : CEMux
    port map (
            O => \N__53133\,
            I => \N__53130\
        );

    \I__12184\ : LocalMux
    port map (
            O => \N__53130\,
            I => \N__53126\
        );

    \I__12183\ : CEMux
    port map (
            O => \N__53129\,
            I => \N__53123\
        );

    \I__12182\ : Span4Mux_v
    port map (
            O => \N__53126\,
            I => \N__53118\
        );

    \I__12181\ : LocalMux
    port map (
            O => \N__53123\,
            I => \N__53118\
        );

    \I__12180\ : Span4Mux_h
    port map (
            O => \N__53118\,
            I => \N__53114\
        );

    \I__12179\ : CEMux
    port map (
            O => \N__53117\,
            I => \N__53111\
        );

    \I__12178\ : Span4Mux_h
    port map (
            O => \N__53114\,
            I => \N__53108\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__53111\,
            I => \N__53105\
        );

    \I__12176\ : Span4Mux_h
    port map (
            O => \N__53108\,
            I => \N__53102\
        );

    \I__12175\ : Span4Mux_v
    port map (
            O => \N__53105\,
            I => \N__53099\
        );

    \I__12174\ : Odrv4
    port map (
            O => \N__53102\,
            I => \dron_frame_decoder_1.N_497_0\
        );

    \I__12173\ : Odrv4
    port map (
            O => \N__53099\,
            I => \dron_frame_decoder_1.N_497_0\
        );

    \I__12172\ : InMux
    port map (
            O => \N__53094\,
            I => \N__53091\
        );

    \I__12171\ : LocalMux
    port map (
            O => \N__53091\,
            I => \N__53088\
        );

    \I__12170\ : Span4Mux_v
    port map (
            O => \N__53088\,
            I => \N__53085\
        );

    \I__12169\ : Odrv4
    port map (
            O => \N__53085\,
            I => \pid_front.O_9\
        );

    \I__12168\ : InMux
    port map (
            O => \N__53082\,
            I => \N__53073\
        );

    \I__12167\ : InMux
    port map (
            O => \N__53081\,
            I => \N__53073\
        );

    \I__12166\ : InMux
    port map (
            O => \N__53080\,
            I => \N__53073\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__53073\,
            I => \N__53070\
        );

    \I__12164\ : Span4Mux_h
    port map (
            O => \N__53070\,
            I => \N__53067\
        );

    \I__12163\ : Span4Mux_h
    port map (
            O => \N__53067\,
            I => \N__53064\
        );

    \I__12162\ : Span4Mux_h
    port map (
            O => \N__53064\,
            I => \N__53061\
        );

    \I__12161\ : Odrv4
    port map (
            O => \N__53061\,
            I => \pid_front.error_d_regZ0Z_5\
        );

    \I__12160\ : InMux
    port map (
            O => \N__53058\,
            I => \N__53055\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__53055\,
            I => \N__53051\
        );

    \I__12158\ : InMux
    port map (
            O => \N__53054\,
            I => \N__53048\
        );

    \I__12157\ : Odrv12
    port map (
            O => \N__53051\,
            I => \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__53048\,
            I => \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1\
        );

    \I__12155\ : CascadeMux
    port map (
            O => \N__53043\,
            I => \N__53040\
        );

    \I__12154\ : InMux
    port map (
            O => \N__53040\,
            I => \N__53037\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__53037\,
            I => \N__53034\
        );

    \I__12152\ : Odrv12
    port map (
            O => \N__53034\,
            I => \pid_side.error_p_reg_esr_RNI5PH23Z0Z_1\
        );

    \I__12151\ : InMux
    port map (
            O => \N__53031\,
            I => \N__53028\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__53028\,
            I => \N__53025\
        );

    \I__12149\ : Odrv4
    port map (
            O => \N__53025\,
            I => \pid_side.O_2_4\
        );

    \I__12148\ : InMux
    port map (
            O => \N__53022\,
            I => \N__53013\
        );

    \I__12147\ : InMux
    port map (
            O => \N__53021\,
            I => \N__53013\
        );

    \I__12146\ : InMux
    port map (
            O => \N__53020\,
            I => \N__53013\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__53013\,
            I => \pid_side.error_p_regZ0Z_0\
        );

    \I__12144\ : InMux
    port map (
            O => \N__53010\,
            I => \N__53007\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__53007\,
            I => \N__53004\
        );

    \I__12142\ : Span4Mux_h
    port map (
            O => \N__53004\,
            I => \N__53001\
        );

    \I__12141\ : Odrv4
    port map (
            O => \N__53001\,
            I => \pid_side.state_RNINK4UZ0Z_0\
        );

    \I__12140\ : InMux
    port map (
            O => \N__52998\,
            I => \N__52992\
        );

    \I__12139\ : InMux
    port map (
            O => \N__52997\,
            I => \N__52992\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__52992\,
            I => \pid_side.error_p_reg_esr_RNIE47JZ0Z_9\
        );

    \I__12137\ : InMux
    port map (
            O => \N__52989\,
            I => \N__52986\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__52986\,
            I => \N__52982\
        );

    \I__12135\ : InMux
    port map (
            O => \N__52985\,
            I => \N__52979\
        );

    \I__12134\ : Odrv4
    port map (
            O => \N__52982\,
            I => \pid_side.error_d_reg_prevZ0Z_15\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__52979\,
            I => \pid_side.error_d_reg_prevZ0Z_15\
        );

    \I__12132\ : InMux
    port map (
            O => \N__52974\,
            I => \N__52971\
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__52971\,
            I => \N__52966\
        );

    \I__12130\ : InMux
    port map (
            O => \N__52970\,
            I => \N__52961\
        );

    \I__12129\ : InMux
    port map (
            O => \N__52969\,
            I => \N__52961\
        );

    \I__12128\ : Odrv4
    port map (
            O => \N__52966\,
            I => \pid_side.un1_pid_prereg_24\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__52961\,
            I => \pid_side.un1_pid_prereg_24\
        );

    \I__12126\ : InMux
    port map (
            O => \N__52956\,
            I => \N__52947\
        );

    \I__12125\ : InMux
    port map (
            O => \N__52955\,
            I => \N__52947\
        );

    \I__12124\ : InMux
    port map (
            O => \N__52954\,
            I => \N__52947\
        );

    \I__12123\ : LocalMux
    port map (
            O => \N__52947\,
            I => \N__52944\
        );

    \I__12122\ : Span4Mux_v
    port map (
            O => \N__52944\,
            I => \N__52941\
        );

    \I__12121\ : Odrv4
    port map (
            O => \N__52941\,
            I => \pid_side.un1_pid_prereg_48\
        );

    \I__12120\ : InMux
    port map (
            O => \N__52938\,
            I => \N__52935\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__52935\,
            I => \N__52931\
        );

    \I__12118\ : InMux
    port map (
            O => \N__52934\,
            I => \N__52928\
        );

    \I__12117\ : Odrv12
    port map (
            O => \N__52931\,
            I => \pid_side.un1_pid_prereg_36\
        );

    \I__12116\ : LocalMux
    port map (
            O => \N__52928\,
            I => \pid_side.un1_pid_prereg_36\
        );

    \I__12115\ : CascadeMux
    port map (
            O => \N__52923\,
            I => \N__52920\
        );

    \I__12114\ : InMux
    port map (
            O => \N__52920\,
            I => \N__52917\
        );

    \I__12113\ : LocalMux
    port map (
            O => \N__52917\,
            I => \N__52914\
        );

    \I__12112\ : Span4Mux_h
    port map (
            O => \N__52914\,
            I => \N__52911\
        );

    \I__12111\ : Odrv4
    port map (
            O => \N__52911\,
            I => \pid_side.error_d_reg_prev_esr_RNIOHC23Z0Z_16\
        );

    \I__12110\ : CascadeMux
    port map (
            O => \N__52908\,
            I => \N__52905\
        );

    \I__12109\ : InMux
    port map (
            O => \N__52905\,
            I => \N__52899\
        );

    \I__12108\ : InMux
    port map (
            O => \N__52904\,
            I => \N__52899\
        );

    \I__12107\ : LocalMux
    port map (
            O => \N__52899\,
            I => \pid_side.error_d_reg_prevZ0Z_18\
        );

    \I__12106\ : InMux
    port map (
            O => \N__52896\,
            I => \N__52893\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__52893\,
            I => \N__52890\
        );

    \I__12104\ : Span4Mux_v
    port map (
            O => \N__52890\,
            I => \N__52886\
        );

    \I__12103\ : InMux
    port map (
            O => \N__52889\,
            I => \N__52883\
        );

    \I__12102\ : Odrv4
    port map (
            O => \N__52886\,
            I => \pid_side.un1_pid_prereg_47\
        );

    \I__12101\ : LocalMux
    port map (
            O => \N__52883\,
            I => \pid_side.un1_pid_prereg_47\
        );

    \I__12100\ : InMux
    port map (
            O => \N__52878\,
            I => \N__52874\
        );

    \I__12099\ : InMux
    port map (
            O => \N__52877\,
            I => \N__52871\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__52874\,
            I => \N__52868\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__52871\,
            I => \N__52865\
        );

    \I__12096\ : Odrv4
    port map (
            O => \N__52868\,
            I => \pid_side.error_d_reg_esr_RNI76TK1Z0Z_5\
        );

    \I__12095\ : Odrv4
    port map (
            O => \N__52865\,
            I => \pid_side.error_d_reg_esr_RNI76TK1Z0Z_5\
        );

    \I__12094\ : CascadeMux
    port map (
            O => \N__52860\,
            I => \pid_side.un1_pid_prereg_40_0_cascade_\
        );

    \I__12093\ : CascadeMux
    port map (
            O => \N__52857\,
            I => \N__52854\
        );

    \I__12092\ : InMux
    port map (
            O => \N__52854\,
            I => \N__52851\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__52851\,
            I => \N__52848\
        );

    \I__12090\ : Odrv4
    port map (
            O => \N__52848\,
            I => \pid_side.error_d_reg_esr_RNI86Q93Z0Z_5\
        );

    \I__12089\ : InMux
    port map (
            O => \N__52845\,
            I => \N__52839\
        );

    \I__12088\ : InMux
    port map (
            O => \N__52844\,
            I => \N__52839\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__52839\,
            I => \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4\
        );

    \I__12086\ : CascadeMux
    port map (
            O => \N__52836\,
            I => \pid_side.un1_pid_prereg_17_cascade_\
        );

    \I__12085\ : InMux
    port map (
            O => \N__52833\,
            I => \N__52830\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__52830\,
            I => \N__52827\
        );

    \I__12083\ : Odrv4
    port map (
            O => \N__52827\,
            I => \pid_side.error_p_reg_esr_RNI10TK1Z0Z_3\
        );

    \I__12082\ : CascadeMux
    port map (
            O => \N__52824\,
            I => \N__52821\
        );

    \I__12081\ : InMux
    port map (
            O => \N__52821\,
            I => \N__52815\
        );

    \I__12080\ : InMux
    port map (
            O => \N__52820\,
            I => \N__52815\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__52815\,
            I => \pid_side.error_d_reg_prevZ0Z_4\
        );

    \I__12078\ : InMux
    port map (
            O => \N__52812\,
            I => \N__52806\
        );

    \I__12077\ : InMux
    port map (
            O => \N__52811\,
            I => \N__52806\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__52806\,
            I => \pid_side.un1_pid_prereg_17\
        );

    \I__12075\ : CascadeMux
    port map (
            O => \N__52803\,
            I => \N__52800\
        );

    \I__12074\ : InMux
    port map (
            O => \N__52800\,
            I => \N__52797\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__52797\,
            I => \N__52794\
        );

    \I__12072\ : Odrv4
    port map (
            O => \N__52794\,
            I => \pid_side.error_p_reg_esr_RNISPP93Z0Z_2\
        );

    \I__12071\ : InMux
    port map (
            O => \N__52791\,
            I => \N__52788\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__52788\,
            I => \N__52785\
        );

    \I__12069\ : Span4Mux_v
    port map (
            O => \N__52785\,
            I => \N__52782\
        );

    \I__12068\ : Odrv4
    port map (
            O => \N__52782\,
            I => \pid_side.O_2_9\
        );

    \I__12067\ : CascadeMux
    port map (
            O => \N__52779\,
            I => \N__52776\
        );

    \I__12066\ : InMux
    port map (
            O => \N__52776\,
            I => \N__52773\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__52773\,
            I => \drone_H_disp_side_i_13\
        );

    \I__12064\ : InMux
    port map (
            O => \N__52770\,
            I => \N__52766\
        );

    \I__12063\ : InMux
    port map (
            O => \N__52769\,
            I => \N__52763\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__52766\,
            I => \N__52760\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__52763\,
            I => \N__52757\
        );

    \I__12060\ : Span12Mux_s4_h
    port map (
            O => \N__52760\,
            I => \N__52754\
        );

    \I__12059\ : Span4Mux_s3_h
    port map (
            O => \N__52757\,
            I => \N__52751\
        );

    \I__12058\ : Odrv12
    port map (
            O => \N__52754\,
            I => \pid_side.error_14\
        );

    \I__12057\ : Odrv4
    port map (
            O => \N__52751\,
            I => \pid_side.error_14\
        );

    \I__12056\ : InMux
    port map (
            O => \N__52746\,
            I => \pid_side.error_cry_9\
        );

    \I__12055\ : InMux
    port map (
            O => \N__52743\,
            I => \pid_side.error_cry_10\
        );

    \I__12054\ : InMux
    port map (
            O => \N__52740\,
            I => \N__52737\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__52737\,
            I => \N__52733\
        );

    \I__12052\ : InMux
    port map (
            O => \N__52736\,
            I => \N__52730\
        );

    \I__12051\ : Span4Mux_s3_h
    port map (
            O => \N__52733\,
            I => \N__52727\
        );

    \I__12050\ : LocalMux
    port map (
            O => \N__52730\,
            I => \N__52724\
        );

    \I__12049\ : Span4Mux_v
    port map (
            O => \N__52727\,
            I => \N__52721\
        );

    \I__12048\ : Span4Mux_s3_h
    port map (
            O => \N__52724\,
            I => \N__52718\
        );

    \I__12047\ : Odrv4
    port map (
            O => \N__52721\,
            I => \pid_side.error_15\
        );

    \I__12046\ : Odrv4
    port map (
            O => \N__52718\,
            I => \pid_side.error_15\
        );

    \I__12045\ : InMux
    port map (
            O => \N__52713\,
            I => \N__52710\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__52710\,
            I => \N__52705\
        );

    \I__12043\ : InMux
    port map (
            O => \N__52709\,
            I => \N__52702\
        );

    \I__12042\ : InMux
    port map (
            O => \N__52708\,
            I => \N__52699\
        );

    \I__12041\ : Span4Mux_h
    port map (
            O => \N__52705\,
            I => \N__52694\
        );

    \I__12040\ : LocalMux
    port map (
            O => \N__52702\,
            I => \N__52694\
        );

    \I__12039\ : LocalMux
    port map (
            O => \N__52699\,
            I => \N__52690\
        );

    \I__12038\ : Span4Mux_v
    port map (
            O => \N__52694\,
            I => \N__52687\
        );

    \I__12037\ : InMux
    port map (
            O => \N__52693\,
            I => \N__52684\
        );

    \I__12036\ : Span4Mux_v
    port map (
            O => \N__52690\,
            I => \N__52680\
        );

    \I__12035\ : Span4Mux_h
    port map (
            O => \N__52687\,
            I => \N__52676\
        );

    \I__12034\ : LocalMux
    port map (
            O => \N__52684\,
            I => \N__52673\
        );

    \I__12033\ : InMux
    port map (
            O => \N__52683\,
            I => \N__52670\
        );

    \I__12032\ : Span4Mux_h
    port map (
            O => \N__52680\,
            I => \N__52667\
        );

    \I__12031\ : InMux
    port map (
            O => \N__52679\,
            I => \N__52664\
        );

    \I__12030\ : Span4Mux_h
    port map (
            O => \N__52676\,
            I => \N__52656\
        );

    \I__12029\ : Span4Mux_v
    port map (
            O => \N__52673\,
            I => \N__52656\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__52670\,
            I => \N__52656\
        );

    \I__12027\ : Span4Mux_v
    port map (
            O => \N__52667\,
            I => \N__52653\
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__52664\,
            I => \N__52650\
        );

    \I__12025\ : CascadeMux
    port map (
            O => \N__52663\,
            I => \N__52646\
        );

    \I__12024\ : Span4Mux_v
    port map (
            O => \N__52656\,
            I => \N__52643\
        );

    \I__12023\ : Span4Mux_v
    port map (
            O => \N__52653\,
            I => \N__52638\
        );

    \I__12022\ : Span4Mux_h
    port map (
            O => \N__52650\,
            I => \N__52638\
        );

    \I__12021\ : InMux
    port map (
            O => \N__52649\,
            I => \N__52635\
        );

    \I__12020\ : InMux
    port map (
            O => \N__52646\,
            I => \N__52632\
        );

    \I__12019\ : Span4Mux_v
    port map (
            O => \N__52643\,
            I => \N__52629\
        );

    \I__12018\ : Span4Mux_v
    port map (
            O => \N__52638\,
            I => \N__52626\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__52635\,
            I => \N__52621\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__52632\,
            I => \N__52621\
        );

    \I__12015\ : Odrv4
    port map (
            O => \N__52629\,
            I => uart_drone_data_3
        );

    \I__12014\ : Odrv4
    port map (
            O => \N__52626\,
            I => uart_drone_data_3
        );

    \I__12013\ : Odrv4
    port map (
            O => \N__52621\,
            I => uart_drone_data_3
        );

    \I__12012\ : InMux
    port map (
            O => \N__52614\,
            I => \N__52608\
        );

    \I__12011\ : InMux
    port map (
            O => \N__52613\,
            I => \N__52608\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__52608\,
            I => \drone_H_disp_side_11\
        );

    \I__12009\ : InMux
    port map (
            O => \N__52605\,
            I => \N__52602\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__52602\,
            I => \N__52599\
        );

    \I__12007\ : Span4Mux_v
    port map (
            O => \N__52599\,
            I => \N__52594\
        );

    \I__12006\ : InMux
    port map (
            O => \N__52598\,
            I => \N__52591\
        );

    \I__12005\ : InMux
    port map (
            O => \N__52597\,
            I => \N__52587\
        );

    \I__12004\ : Span4Mux_h
    port map (
            O => \N__52594\,
            I => \N__52583\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__52591\,
            I => \N__52580\
        );

    \I__12002\ : InMux
    port map (
            O => \N__52590\,
            I => \N__52577\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__52587\,
            I => \N__52573\
        );

    \I__12000\ : InMux
    port map (
            O => \N__52586\,
            I => \N__52570\
        );

    \I__11999\ : Span4Mux_h
    port map (
            O => \N__52583\,
            I => \N__52565\
        );

    \I__11998\ : Span4Mux_v
    port map (
            O => \N__52580\,
            I => \N__52565\
        );

    \I__11997\ : LocalMux
    port map (
            O => \N__52577\,
            I => \N__52562\
        );

    \I__11996\ : InMux
    port map (
            O => \N__52576\,
            I => \N__52559\
        );

    \I__11995\ : Span4Mux_h
    port map (
            O => \N__52573\,
            I => \N__52556\
        );

    \I__11994\ : LocalMux
    port map (
            O => \N__52570\,
            I => \N__52553\
        );

    \I__11993\ : Span4Mux_h
    port map (
            O => \N__52565\,
            I => \N__52546\
        );

    \I__11992\ : Span4Mux_v
    port map (
            O => \N__52562\,
            I => \N__52546\
        );

    \I__11991\ : LocalMux
    port map (
            O => \N__52559\,
            I => \N__52546\
        );

    \I__11990\ : Span4Mux_v
    port map (
            O => \N__52556\,
            I => \N__52543\
        );

    \I__11989\ : Sp12to4
    port map (
            O => \N__52553\,
            I => \N__52538\
        );

    \I__11988\ : Span4Mux_v
    port map (
            O => \N__52546\,
            I => \N__52535\
        );

    \I__11987\ : Span4Mux_v
    port map (
            O => \N__52543\,
            I => \N__52532\
        );

    \I__11986\ : InMux
    port map (
            O => \N__52542\,
            I => \N__52529\
        );

    \I__11985\ : InMux
    port map (
            O => \N__52541\,
            I => \N__52526\
        );

    \I__11984\ : Span12Mux_v
    port map (
            O => \N__52538\,
            I => \N__52523\
        );

    \I__11983\ : Span4Mux_v
    port map (
            O => \N__52535\,
            I => \N__52520\
        );

    \I__11982\ : Span4Mux_v
    port map (
            O => \N__52532\,
            I => \N__52513\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__52529\,
            I => \N__52513\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__52526\,
            I => \N__52513\
        );

    \I__11979\ : Odrv12
    port map (
            O => \N__52523\,
            I => uart_drone_data_4
        );

    \I__11978\ : Odrv4
    port map (
            O => \N__52520\,
            I => uart_drone_data_4
        );

    \I__11977\ : Odrv4
    port map (
            O => \N__52513\,
            I => uart_drone_data_4
        );

    \I__11976\ : CascadeMux
    port map (
            O => \N__52506\,
            I => \N__52503\
        );

    \I__11975\ : InMux
    port map (
            O => \N__52503\,
            I => \N__52498\
        );

    \I__11974\ : InMux
    port map (
            O => \N__52502\,
            I => \N__52493\
        );

    \I__11973\ : InMux
    port map (
            O => \N__52501\,
            I => \N__52493\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__52498\,
            I => \drone_H_disp_side_12\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__52493\,
            I => \drone_H_disp_side_12\
        );

    \I__11970\ : InMux
    port map (
            O => \N__52488\,
            I => \N__52485\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__52485\,
            I => \N__52481\
        );

    \I__11968\ : InMux
    port map (
            O => \N__52484\,
            I => \N__52478\
        );

    \I__11967\ : Span4Mux_v
    port map (
            O => \N__52481\,
            I => \N__52472\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__52478\,
            I => \N__52472\
        );

    \I__11965\ : InMux
    port map (
            O => \N__52477\,
            I => \N__52469\
        );

    \I__11964\ : Span4Mux_h
    port map (
            O => \N__52472\,
            I => \N__52464\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__52469\,
            I => \N__52461\
        );

    \I__11962\ : InMux
    port map (
            O => \N__52468\,
            I => \N__52458\
        );

    \I__11961\ : InMux
    port map (
            O => \N__52467\,
            I => \N__52454\
        );

    \I__11960\ : Span4Mux_h
    port map (
            O => \N__52464\,
            I => \N__52449\
        );

    \I__11959\ : Span4Mux_v
    port map (
            O => \N__52461\,
            I => \N__52449\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__52458\,
            I => \N__52446\
        );

    \I__11957\ : InMux
    port map (
            O => \N__52457\,
            I => \N__52443\
        );

    \I__11956\ : LocalMux
    port map (
            O => \N__52454\,
            I => \N__52440\
        );

    \I__11955\ : Span4Mux_h
    port map (
            O => \N__52449\,
            I => \N__52433\
        );

    \I__11954\ : Span4Mux_v
    port map (
            O => \N__52446\,
            I => \N__52433\
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__52443\,
            I => \N__52433\
        );

    \I__11952\ : Sp12to4
    port map (
            O => \N__52440\,
            I => \N__52430\
        );

    \I__11951\ : Span4Mux_v
    port map (
            O => \N__52433\,
            I => \N__52427\
        );

    \I__11950\ : Span12Mux_v
    port map (
            O => \N__52430\,
            I => \N__52423\
        );

    \I__11949\ : Span4Mux_v
    port map (
            O => \N__52427\,
            I => \N__52420\
        );

    \I__11948\ : InMux
    port map (
            O => \N__52426\,
            I => \N__52417\
        );

    \I__11947\ : Odrv12
    port map (
            O => \N__52423\,
            I => uart_drone_data_5
        );

    \I__11946\ : Odrv4
    port map (
            O => \N__52420\,
            I => uart_drone_data_5
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__52417\,
            I => uart_drone_data_5
        );

    \I__11944\ : CascadeMux
    port map (
            O => \N__52410\,
            I => \N__52407\
        );

    \I__11943\ : InMux
    port map (
            O => \N__52407\,
            I => \N__52403\
        );

    \I__11942\ : InMux
    port map (
            O => \N__52406\,
            I => \N__52400\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__52403\,
            I => \drone_H_disp_side_13\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__52400\,
            I => \drone_H_disp_side_13\
        );

    \I__11939\ : InMux
    port map (
            O => \N__52395\,
            I => \N__52392\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__52392\,
            I => \N__52388\
        );

    \I__11937\ : InMux
    port map (
            O => \N__52391\,
            I => \N__52385\
        );

    \I__11936\ : Span4Mux_v
    port map (
            O => \N__52388\,
            I => \N__52379\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__52385\,
            I => \N__52379\
        );

    \I__11934\ : InMux
    port map (
            O => \N__52384\,
            I => \N__52375\
        );

    \I__11933\ : Span4Mux_v
    port map (
            O => \N__52379\,
            I => \N__52371\
        );

    \I__11932\ : InMux
    port map (
            O => \N__52378\,
            I => \N__52368\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__52375\,
            I => \N__52365\
        );

    \I__11930\ : InMux
    port map (
            O => \N__52374\,
            I => \N__52362\
        );

    \I__11929\ : Span4Mux_h
    port map (
            O => \N__52371\,
            I => \N__52356\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__52368\,
            I => \N__52356\
        );

    \I__11927\ : Span4Mux_h
    port map (
            O => \N__52365\,
            I => \N__52351\
        );

    \I__11926\ : LocalMux
    port map (
            O => \N__52362\,
            I => \N__52351\
        );

    \I__11925\ : InMux
    port map (
            O => \N__52361\,
            I => \N__52348\
        );

    \I__11924\ : Span4Mux_v
    port map (
            O => \N__52356\,
            I => \N__52344\
        );

    \I__11923\ : Sp12to4
    port map (
            O => \N__52351\,
            I => \N__52341\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__52348\,
            I => \N__52338\
        );

    \I__11921\ : CascadeMux
    port map (
            O => \N__52347\,
            I => \N__52335\
        );

    \I__11920\ : Span4Mux_v
    port map (
            O => \N__52344\,
            I => \N__52332\
        );

    \I__11919\ : Span12Mux_v
    port map (
            O => \N__52341\,
            I => \N__52327\
        );

    \I__11918\ : Span12Mux_v
    port map (
            O => \N__52338\,
            I => \N__52327\
        );

    \I__11917\ : InMux
    port map (
            O => \N__52335\,
            I => \N__52324\
        );

    \I__11916\ : Odrv4
    port map (
            O => \N__52332\,
            I => uart_drone_data_7
        );

    \I__11915\ : Odrv12
    port map (
            O => \N__52327\,
            I => uart_drone_data_7
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__52324\,
            I => uart_drone_data_7
        );

    \I__11913\ : InMux
    port map (
            O => \N__52317\,
            I => \N__52314\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__52314\,
            I => \drone_H_disp_side_15\
        );

    \I__11911\ : InMux
    port map (
            O => \N__52311\,
            I => \N__52308\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__52308\,
            I => \N__52304\
        );

    \I__11909\ : InMux
    port map (
            O => \N__52307\,
            I => \N__52301\
        );

    \I__11908\ : Span4Mux_v
    port map (
            O => \N__52304\,
            I => \N__52295\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__52301\,
            I => \N__52295\
        );

    \I__11906\ : InMux
    port map (
            O => \N__52300\,
            I => \N__52292\
        );

    \I__11905\ : Span4Mux_v
    port map (
            O => \N__52295\,
            I => \N__52288\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__52292\,
            I => \N__52285\
        );

    \I__11903\ : InMux
    port map (
            O => \N__52291\,
            I => \N__52282\
        );

    \I__11902\ : Span4Mux_h
    port map (
            O => \N__52288\,
            I => \N__52279\
        );

    \I__11901\ : Span4Mux_v
    port map (
            O => \N__52285\,
            I => \N__52274\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__52282\,
            I => \N__52274\
        );

    \I__11899\ : Span4Mux_h
    port map (
            O => \N__52279\,
            I => \N__52268\
        );

    \I__11898\ : Span4Mux_v
    port map (
            O => \N__52274\,
            I => \N__52268\
        );

    \I__11897\ : InMux
    port map (
            O => \N__52273\,
            I => \N__52265\
        );

    \I__11896\ : Span4Mux_h
    port map (
            O => \N__52268\,
            I => \N__52260\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__52265\,
            I => \N__52260\
        );

    \I__11894\ : Span4Mux_v
    port map (
            O => \N__52260\,
            I => \N__52256\
        );

    \I__11893\ : InMux
    port map (
            O => \N__52259\,
            I => \N__52253\
        );

    \I__11892\ : Sp12to4
    port map (
            O => \N__52256\,
            I => \N__52248\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__52253\,
            I => \N__52248\
        );

    \I__11890\ : Span12Mux_s10_h
    port map (
            O => \N__52248\,
            I => \N__52244\
        );

    \I__11889\ : InMux
    port map (
            O => \N__52247\,
            I => \N__52241\
        );

    \I__11888\ : Odrv12
    port map (
            O => \N__52244\,
            I => uart_drone_data_0
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__52241\,
            I => uart_drone_data_0
        );

    \I__11886\ : InMux
    port map (
            O => \N__52236\,
            I => \N__52233\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__52233\,
            I => \dron_frame_decoder_1.drone_H_disp_side_8\
        );

    \I__11884\ : InMux
    port map (
            O => \N__52230\,
            I => \N__52227\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__52227\,
            I => \N__52224\
        );

    \I__11882\ : Span4Mux_h
    port map (
            O => \N__52224\,
            I => \N__52221\
        );

    \I__11881\ : Odrv4
    port map (
            O => \N__52221\,
            I => \pid_front.O_10\
        );

    \I__11880\ : InMux
    port map (
            O => \N__52218\,
            I => \N__52213\
        );

    \I__11879\ : InMux
    port map (
            O => \N__52217\,
            I => \N__52208\
        );

    \I__11878\ : InMux
    port map (
            O => \N__52216\,
            I => \N__52208\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__52213\,
            I => \N__52203\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__52208\,
            I => \N__52203\
        );

    \I__11875\ : Span4Mux_h
    port map (
            O => \N__52203\,
            I => \N__52200\
        );

    \I__11874\ : Span4Mux_h
    port map (
            O => \N__52200\,
            I => \N__52197\
        );

    \I__11873\ : Span4Mux_h
    port map (
            O => \N__52197\,
            I => \N__52194\
        );

    \I__11872\ : Odrv4
    port map (
            O => \N__52194\,
            I => \pid_front.error_d_regZ0Z_6\
        );

    \I__11871\ : InMux
    port map (
            O => \N__52191\,
            I => \N__52188\
        );

    \I__11870\ : LocalMux
    port map (
            O => \N__52188\,
            I => \drone_H_disp_side_i_6\
        );

    \I__11869\ : CascadeMux
    port map (
            O => \N__52185\,
            I => \N__52182\
        );

    \I__11868\ : InMux
    port map (
            O => \N__52182\,
            I => \N__52179\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__52179\,
            I => \N__52176\
        );

    \I__11866\ : Odrv4
    port map (
            O => \N__52176\,
            I => side_command_2
        );

    \I__11865\ : InMux
    port map (
            O => \N__52173\,
            I => \N__52170\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__52170\,
            I => \N__52167\
        );

    \I__11863\ : Span4Mux_s3_h
    port map (
            O => \N__52167\,
            I => \N__52163\
        );

    \I__11862\ : InMux
    port map (
            O => \N__52166\,
            I => \N__52160\
        );

    \I__11861\ : Span4Mux_v
    port map (
            O => \N__52163\,
            I => \N__52157\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__52160\,
            I => \N__52154\
        );

    \I__11859\ : Odrv4
    port map (
            O => \N__52157\,
            I => \pid_side.error_6\
        );

    \I__11858\ : Odrv12
    port map (
            O => \N__52154\,
            I => \pid_side.error_6\
        );

    \I__11857\ : InMux
    port map (
            O => \N__52149\,
            I => \pid_side.error_cry_1_0\
        );

    \I__11856\ : InMux
    port map (
            O => \N__52146\,
            I => \N__52143\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__52143\,
            I => \drone_H_disp_side_i_7\
        );

    \I__11854\ : CascadeMux
    port map (
            O => \N__52140\,
            I => \N__52137\
        );

    \I__11853\ : InMux
    port map (
            O => \N__52137\,
            I => \N__52134\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__52134\,
            I => side_command_3
        );

    \I__11851\ : InMux
    port map (
            O => \N__52131\,
            I => \N__52128\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__52128\,
            I => \N__52124\
        );

    \I__11849\ : InMux
    port map (
            O => \N__52127\,
            I => \N__52121\
        );

    \I__11848\ : Span12Mux_s4_h
    port map (
            O => \N__52124\,
            I => \N__52118\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__52121\,
            I => \N__52115\
        );

    \I__11846\ : Odrv12
    port map (
            O => \N__52118\,
            I => \pid_side.error_7\
        );

    \I__11845\ : Odrv12
    port map (
            O => \N__52115\,
            I => \pid_side.error_7\
        );

    \I__11844\ : InMux
    port map (
            O => \N__52110\,
            I => \pid_side.error_cry_2_0\
        );

    \I__11843\ : InMux
    port map (
            O => \N__52107\,
            I => \N__52104\
        );

    \I__11842\ : LocalMux
    port map (
            O => \N__52104\,
            I => \drone_H_disp_side_i_8\
        );

    \I__11841\ : CascadeMux
    port map (
            O => \N__52101\,
            I => \N__52098\
        );

    \I__11840\ : InMux
    port map (
            O => \N__52098\,
            I => \N__52095\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__52095\,
            I => \N__52092\
        );

    \I__11838\ : Span4Mux_h
    port map (
            O => \N__52092\,
            I => \N__52089\
        );

    \I__11837\ : Odrv4
    port map (
            O => \N__52089\,
            I => side_command_4
        );

    \I__11836\ : InMux
    port map (
            O => \N__52086\,
            I => \N__52083\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__52083\,
            I => \N__52079\
        );

    \I__11834\ : InMux
    port map (
            O => \N__52082\,
            I => \N__52076\
        );

    \I__11833\ : Span4Mux_v
    port map (
            O => \N__52079\,
            I => \N__52071\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__52076\,
            I => \N__52071\
        );

    \I__11831\ : Span4Mux_v
    port map (
            O => \N__52071\,
            I => \N__52068\
        );

    \I__11830\ : Odrv4
    port map (
            O => \N__52068\,
            I => \pid_side.error_8\
        );

    \I__11829\ : InMux
    port map (
            O => \N__52065\,
            I => \bfn_21_18_0_\
        );

    \I__11828\ : InMux
    port map (
            O => \N__52062\,
            I => \N__52059\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__52059\,
            I => \N__52056\
        );

    \I__11826\ : Span4Mux_v
    port map (
            O => \N__52056\,
            I => \N__52053\
        );

    \I__11825\ : Span4Mux_h
    port map (
            O => \N__52053\,
            I => \N__52050\
        );

    \I__11824\ : Span4Mux_h
    port map (
            O => \N__52050\,
            I => \N__52047\
        );

    \I__11823\ : Odrv4
    port map (
            O => \N__52047\,
            I => \drone_H_disp_side_i_9\
        );

    \I__11822\ : CascadeMux
    port map (
            O => \N__52044\,
            I => \N__52041\
        );

    \I__11821\ : InMux
    port map (
            O => \N__52041\,
            I => \N__52038\
        );

    \I__11820\ : LocalMux
    port map (
            O => \N__52038\,
            I => \N__52035\
        );

    \I__11819\ : Odrv4
    port map (
            O => \N__52035\,
            I => side_command_5
        );

    \I__11818\ : InMux
    port map (
            O => \N__52032\,
            I => \N__52029\
        );

    \I__11817\ : LocalMux
    port map (
            O => \N__52029\,
            I => \N__52025\
        );

    \I__11816\ : InMux
    port map (
            O => \N__52028\,
            I => \N__52022\
        );

    \I__11815\ : Span4Mux_v
    port map (
            O => \N__52025\,
            I => \N__52017\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__52022\,
            I => \N__52017\
        );

    \I__11813\ : Span4Mux_v
    port map (
            O => \N__52017\,
            I => \N__52014\
        );

    \I__11812\ : Odrv4
    port map (
            O => \N__52014\,
            I => \pid_side.error_9\
        );

    \I__11811\ : InMux
    port map (
            O => \N__52011\,
            I => \pid_side.error_cry_4\
        );

    \I__11810\ : InMux
    port map (
            O => \N__52008\,
            I => \N__52005\
        );

    \I__11809\ : LocalMux
    port map (
            O => \N__52005\,
            I => \N__52002\
        );

    \I__11808\ : Span12Mux_s6_h
    port map (
            O => \N__52002\,
            I => \N__51999\
        );

    \I__11807\ : Odrv12
    port map (
            O => \N__51999\,
            I => \drone_H_disp_side_i_10\
        );

    \I__11806\ : CascadeMux
    port map (
            O => \N__51996\,
            I => \N__51993\
        );

    \I__11805\ : InMux
    port map (
            O => \N__51993\,
            I => \N__51990\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__51990\,
            I => \N__51987\
        );

    \I__11803\ : Span4Mux_h
    port map (
            O => \N__51987\,
            I => \N__51984\
        );

    \I__11802\ : Odrv4
    port map (
            O => \N__51984\,
            I => side_command_6
        );

    \I__11801\ : InMux
    port map (
            O => \N__51981\,
            I => \N__51978\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__51978\,
            I => \N__51974\
        );

    \I__11799\ : InMux
    port map (
            O => \N__51977\,
            I => \N__51971\
        );

    \I__11798\ : Span4Mux_v
    port map (
            O => \N__51974\,
            I => \N__51968\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__51971\,
            I => \N__51965\
        );

    \I__11796\ : Span4Mux_h
    port map (
            O => \N__51968\,
            I => \N__51962\
        );

    \I__11795\ : Span4Mux_s3_h
    port map (
            O => \N__51965\,
            I => \N__51959\
        );

    \I__11794\ : Odrv4
    port map (
            O => \N__51962\,
            I => \pid_side.error_10\
        );

    \I__11793\ : Odrv4
    port map (
            O => \N__51959\,
            I => \pid_side.error_10\
        );

    \I__11792\ : InMux
    port map (
            O => \N__51954\,
            I => \pid_side.error_cry_5\
        );

    \I__11791\ : InMux
    port map (
            O => \N__51951\,
            I => \N__51948\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__51948\,
            I => \pid_side.error_axbZ0Z_7\
        );

    \I__11789\ : InMux
    port map (
            O => \N__51945\,
            I => \N__51942\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__51942\,
            I => \N__51938\
        );

    \I__11787\ : InMux
    port map (
            O => \N__51941\,
            I => \N__51935\
        );

    \I__11786\ : Span4Mux_v
    port map (
            O => \N__51938\,
            I => \N__51932\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__51935\,
            I => \N__51929\
        );

    \I__11784\ : Span4Mux_h
    port map (
            O => \N__51932\,
            I => \N__51926\
        );

    \I__11783\ : Span4Mux_s3_h
    port map (
            O => \N__51929\,
            I => \N__51923\
        );

    \I__11782\ : Odrv4
    port map (
            O => \N__51926\,
            I => \pid_side.error_11\
        );

    \I__11781\ : Odrv4
    port map (
            O => \N__51923\,
            I => \pid_side.error_11\
        );

    \I__11780\ : InMux
    port map (
            O => \N__51918\,
            I => \pid_side.error_cry_6\
        );

    \I__11779\ : InMux
    port map (
            O => \N__51915\,
            I => \N__51912\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__51912\,
            I => \pid_side.error_axb_8_l_ofxZ0\
        );

    \I__11777\ : InMux
    port map (
            O => \N__51909\,
            I => \N__51906\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__51906\,
            I => \N__51902\
        );

    \I__11775\ : InMux
    port map (
            O => \N__51905\,
            I => \N__51899\
        );

    \I__11774\ : Span4Mux_s3_h
    port map (
            O => \N__51902\,
            I => \N__51896\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__51899\,
            I => \N__51893\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__51896\,
            I => \N__51890\
        );

    \I__11771\ : Span4Mux_s3_h
    port map (
            O => \N__51893\,
            I => \N__51887\
        );

    \I__11770\ : Odrv4
    port map (
            O => \N__51890\,
            I => \pid_side.error_12\
        );

    \I__11769\ : Odrv4
    port map (
            O => \N__51887\,
            I => \pid_side.error_12\
        );

    \I__11768\ : InMux
    port map (
            O => \N__51882\,
            I => \pid_side.error_cry_7\
        );

    \I__11767\ : InMux
    port map (
            O => \N__51879\,
            I => \N__51876\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__51876\,
            I => \drone_H_disp_side_i_12\
        );

    \I__11765\ : InMux
    port map (
            O => \N__51873\,
            I => \N__51870\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__51870\,
            I => \N__51866\
        );

    \I__11763\ : InMux
    port map (
            O => \N__51869\,
            I => \N__51863\
        );

    \I__11762\ : Span4Mux_s3_h
    port map (
            O => \N__51866\,
            I => \N__51860\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__51863\,
            I => \N__51857\
        );

    \I__11760\ : Span4Mux_v
    port map (
            O => \N__51860\,
            I => \N__51854\
        );

    \I__11759\ : Span4Mux_s3_h
    port map (
            O => \N__51857\,
            I => \N__51851\
        );

    \I__11758\ : Odrv4
    port map (
            O => \N__51854\,
            I => \pid_side.error_13\
        );

    \I__11757\ : Odrv4
    port map (
            O => \N__51851\,
            I => \pid_side.error_13\
        );

    \I__11756\ : InMux
    port map (
            O => \N__51846\,
            I => \pid_side.error_cry_8\
        );

    \I__11755\ : InMux
    port map (
            O => \N__51843\,
            I => \N__51837\
        );

    \I__11754\ : InMux
    port map (
            O => \N__51842\,
            I => \N__51837\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__51837\,
            I => \pid_side.error_d_reg_prevZ0Z_19\
        );

    \I__11752\ : CascadeMux
    port map (
            O => \N__51834\,
            I => \N__51830\
        );

    \I__11751\ : InMux
    port map (
            O => \N__51833\,
            I => \N__51827\
        );

    \I__11750\ : InMux
    port map (
            O => \N__51830\,
            I => \N__51823\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__51827\,
            I => \N__51820\
        );

    \I__11748\ : InMux
    port map (
            O => \N__51826\,
            I => \N__51817\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__51823\,
            I => \pid_side.un1_pid_prereg_57\
        );

    \I__11746\ : Odrv4
    port map (
            O => \N__51820\,
            I => \pid_side.un1_pid_prereg_57\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__51817\,
            I => \pid_side.un1_pid_prereg_57\
        );

    \I__11744\ : CEMux
    port map (
            O => \N__51810\,
            I => \N__51806\
        );

    \I__11743\ : CEMux
    port map (
            O => \N__51809\,
            I => \N__51803\
        );

    \I__11742\ : LocalMux
    port map (
            O => \N__51806\,
            I => \N__51800\
        );

    \I__11741\ : LocalMux
    port map (
            O => \N__51803\,
            I => \N__51797\
        );

    \I__11740\ : Span4Mux_h
    port map (
            O => \N__51800\,
            I => \N__51794\
        );

    \I__11739\ : Span4Mux_h
    port map (
            O => \N__51797\,
            I => \N__51789\
        );

    \I__11738\ : Span4Mux_h
    port map (
            O => \N__51794\,
            I => \N__51789\
        );

    \I__11737\ : Odrv4
    port map (
            O => \N__51789\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__11736\ : InMux
    port map (
            O => \N__51786\,
            I => \N__51783\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__51783\,
            I => \N__51780\
        );

    \I__11734\ : Span4Mux_v
    port map (
            O => \N__51780\,
            I => \N__51776\
        );

    \I__11733\ : InMux
    port map (
            O => \N__51779\,
            I => \N__51773\
        );

    \I__11732\ : Span4Mux_h
    port map (
            O => \N__51776\,
            I => \N__51769\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__51773\,
            I => \N__51766\
        );

    \I__11730\ : InMux
    port map (
            O => \N__51772\,
            I => \N__51763\
        );

    \I__11729\ : Odrv4
    port map (
            O => \N__51769\,
            I => \drone_H_disp_side_0\
        );

    \I__11728\ : Odrv12
    port map (
            O => \N__51766\,
            I => \drone_H_disp_side_0\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__51763\,
            I => \drone_H_disp_side_0\
        );

    \I__11726\ : InMux
    port map (
            O => \N__51756\,
            I => \N__51753\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__51753\,
            I => \pid_side.error_axb_0\
        );

    \I__11724\ : InMux
    port map (
            O => \N__51750\,
            I => \N__51747\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__51747\,
            I => \pid_side.error_axbZ0Z_1\
        );

    \I__11722\ : InMux
    port map (
            O => \N__51744\,
            I => \N__51741\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__51741\,
            I => \N__51737\
        );

    \I__11720\ : InMux
    port map (
            O => \N__51740\,
            I => \N__51734\
        );

    \I__11719\ : Span4Mux_v
    port map (
            O => \N__51737\,
            I => \N__51731\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__51734\,
            I => \N__51728\
        );

    \I__11717\ : Span4Mux_h
    port map (
            O => \N__51731\,
            I => \N__51725\
        );

    \I__11716\ : Span4Mux_s1_h
    port map (
            O => \N__51728\,
            I => \N__51722\
        );

    \I__11715\ : Odrv4
    port map (
            O => \N__51725\,
            I => \pid_side.error_1\
        );

    \I__11714\ : Odrv4
    port map (
            O => \N__51722\,
            I => \pid_side.error_1\
        );

    \I__11713\ : InMux
    port map (
            O => \N__51717\,
            I => \pid_side.error_cry_0\
        );

    \I__11712\ : InMux
    port map (
            O => \N__51714\,
            I => \N__51711\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__51711\,
            I => \pid_side.error_axbZ0Z_2\
        );

    \I__11710\ : InMux
    port map (
            O => \N__51708\,
            I => \N__51705\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__51705\,
            I => \N__51701\
        );

    \I__11708\ : InMux
    port map (
            O => \N__51704\,
            I => \N__51698\
        );

    \I__11707\ : Span4Mux_v
    port map (
            O => \N__51701\,
            I => \N__51695\
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__51698\,
            I => \N__51692\
        );

    \I__11705\ : Span4Mux_h
    port map (
            O => \N__51695\,
            I => \N__51689\
        );

    \I__11704\ : Span4Mux_s1_h
    port map (
            O => \N__51692\,
            I => \N__51686\
        );

    \I__11703\ : Odrv4
    port map (
            O => \N__51689\,
            I => \pid_side.error_2\
        );

    \I__11702\ : Odrv4
    port map (
            O => \N__51686\,
            I => \pid_side.error_2\
        );

    \I__11701\ : InMux
    port map (
            O => \N__51681\,
            I => \pid_side.error_cry_1\
        );

    \I__11700\ : InMux
    port map (
            O => \N__51678\,
            I => \N__51675\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__51675\,
            I => \pid_side.error_axbZ0Z_3\
        );

    \I__11698\ : InMux
    port map (
            O => \N__51672\,
            I => \N__51669\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__51669\,
            I => \N__51666\
        );

    \I__11696\ : Span4Mux_v
    port map (
            O => \N__51666\,
            I => \N__51662\
        );

    \I__11695\ : InMux
    port map (
            O => \N__51665\,
            I => \N__51659\
        );

    \I__11694\ : Span4Mux_v
    port map (
            O => \N__51662\,
            I => \N__51654\
        );

    \I__11693\ : LocalMux
    port map (
            O => \N__51659\,
            I => \N__51654\
        );

    \I__11692\ : Span4Mux_s0_h
    port map (
            O => \N__51654\,
            I => \N__51651\
        );

    \I__11691\ : Odrv4
    port map (
            O => \N__51651\,
            I => \pid_side.error_3\
        );

    \I__11690\ : InMux
    port map (
            O => \N__51648\,
            I => \pid_side.error_cry_2\
        );

    \I__11689\ : InMux
    port map (
            O => \N__51645\,
            I => \N__51642\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__51642\,
            I => \drone_H_disp_side_i_4\
        );

    \I__11687\ : CascadeMux
    port map (
            O => \N__51639\,
            I => \N__51636\
        );

    \I__11686\ : InMux
    port map (
            O => \N__51636\,
            I => \N__51633\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__51633\,
            I => \N__51630\
        );

    \I__11684\ : Odrv4
    port map (
            O => \N__51630\,
            I => side_command_0
        );

    \I__11683\ : InMux
    port map (
            O => \N__51627\,
            I => \N__51624\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__51624\,
            I => \N__51621\
        );

    \I__11681\ : Span4Mux_s3_h
    port map (
            O => \N__51621\,
            I => \N__51617\
        );

    \I__11680\ : InMux
    port map (
            O => \N__51620\,
            I => \N__51614\
        );

    \I__11679\ : Span4Mux_v
    port map (
            O => \N__51617\,
            I => \N__51611\
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__51614\,
            I => \N__51608\
        );

    \I__11677\ : Odrv4
    port map (
            O => \N__51611\,
            I => \pid_side.error_4\
        );

    \I__11676\ : Odrv12
    port map (
            O => \N__51608\,
            I => \pid_side.error_4\
        );

    \I__11675\ : InMux
    port map (
            O => \N__51603\,
            I => \pid_side.error_cry_3\
        );

    \I__11674\ : InMux
    port map (
            O => \N__51600\,
            I => \N__51597\
        );

    \I__11673\ : LocalMux
    port map (
            O => \N__51597\,
            I => \N__51594\
        );

    \I__11672\ : Odrv4
    port map (
            O => \N__51594\,
            I => \drone_H_disp_side_i_5\
        );

    \I__11671\ : CascadeMux
    port map (
            O => \N__51591\,
            I => \N__51588\
        );

    \I__11670\ : InMux
    port map (
            O => \N__51588\,
            I => \N__51585\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__51585\,
            I => side_command_1
        );

    \I__11668\ : InMux
    port map (
            O => \N__51582\,
            I => \N__51579\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__51579\,
            I => \N__51576\
        );

    \I__11666\ : Span4Mux_s3_h
    port map (
            O => \N__51576\,
            I => \N__51572\
        );

    \I__11665\ : InMux
    port map (
            O => \N__51575\,
            I => \N__51569\
        );

    \I__11664\ : Span4Mux_v
    port map (
            O => \N__51572\,
            I => \N__51566\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__51569\,
            I => \N__51563\
        );

    \I__11662\ : Odrv4
    port map (
            O => \N__51566\,
            I => \pid_side.error_5\
        );

    \I__11661\ : Odrv12
    port map (
            O => \N__51563\,
            I => \pid_side.error_5\
        );

    \I__11660\ : InMux
    port map (
            O => \N__51558\,
            I => \pid_side.error_cry_0_0\
        );

    \I__11659\ : InMux
    port map (
            O => \N__51555\,
            I => \N__51552\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__51552\,
            I => \pid_side.un1_pid_prereg_107_0\
        );

    \I__11657\ : InMux
    port map (
            O => \N__51549\,
            I => \N__51545\
        );

    \I__11656\ : InMux
    port map (
            O => \N__51548\,
            I => \N__51542\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__51545\,
            I => \pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__51542\,
            I => \pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11\
        );

    \I__11653\ : InMux
    port map (
            O => \N__51537\,
            I => \N__51528\
        );

    \I__11652\ : InMux
    port map (
            O => \N__51536\,
            I => \N__51528\
        );

    \I__11651\ : InMux
    port map (
            O => \N__51535\,
            I => \N__51528\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__51528\,
            I => \pid_side.error_d_reg_prevZ0Z_12\
        );

    \I__11649\ : InMux
    port map (
            O => \N__51525\,
            I => \N__51520\
        );

    \I__11648\ : InMux
    port map (
            O => \N__51524\,
            I => \N__51515\
        );

    \I__11647\ : InMux
    port map (
            O => \N__51523\,
            I => \N__51515\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__51520\,
            I => \N__51510\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__51515\,
            I => \N__51510\
        );

    \I__11644\ : Odrv12
    port map (
            O => \N__51510\,
            I => \pid_side.error_d_reg_prev_esr_RNI2VN9Z0Z_12\
        );

    \I__11643\ : InMux
    port map (
            O => \N__51507\,
            I => \N__51503\
        );

    \I__11642\ : InMux
    port map (
            O => \N__51506\,
            I => \N__51500\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__51503\,
            I => \pid_side.error_d_reg_prevZ0Z_11\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__51500\,
            I => \pid_side.error_d_reg_prevZ0Z_11\
        );

    \I__11639\ : InMux
    port map (
            O => \N__51495\,
            I => \N__51492\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__51492\,
            I => \N__51489\
        );

    \I__11637\ : Span4Mux_h
    port map (
            O => \N__51489\,
            I => \N__51486\
        );

    \I__11636\ : Odrv4
    port map (
            O => \N__51486\,
            I => \pid_side.O_2_15\
        );

    \I__11635\ : InMux
    port map (
            O => \N__51483\,
            I => \N__51479\
        );

    \I__11634\ : InMux
    port map (
            O => \N__51482\,
            I => \N__51476\
        );

    \I__11633\ : LocalMux
    port map (
            O => \N__51479\,
            I => \N__51473\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__51476\,
            I => \pid_side.error_p_regZ0Z_11\
        );

    \I__11631\ : Odrv4
    port map (
            O => \N__51473\,
            I => \pid_side.error_p_regZ0Z_11\
        );

    \I__11630\ : InMux
    port map (
            O => \N__51468\,
            I => \N__51465\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__51465\,
            I => \N__51462\
        );

    \I__11628\ : Span12Mux_s9_h
    port map (
            O => \N__51462\,
            I => \N__51459\
        );

    \I__11627\ : Odrv12
    port map (
            O => \N__51459\,
            I => \ppm_encoder_1.N_291\
        );

    \I__11626\ : InMux
    port map (
            O => \N__51456\,
            I => \N__51453\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__51453\,
            I => \N__51445\
        );

    \I__11624\ : InMux
    port map (
            O => \N__51452\,
            I => \N__51442\
        );

    \I__11623\ : InMux
    port map (
            O => \N__51451\,
            I => \N__51437\
        );

    \I__11622\ : InMux
    port map (
            O => \N__51450\,
            I => \N__51437\
        );

    \I__11621\ : CascadeMux
    port map (
            O => \N__51449\,
            I => \N__51433\
        );

    \I__11620\ : CascadeMux
    port map (
            O => \N__51448\,
            I => \N__51428\
        );

    \I__11619\ : Span4Mux_v
    port map (
            O => \N__51445\,
            I => \N__51419\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__51442\,
            I => \N__51419\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__51437\,
            I => \N__51419\
        );

    \I__11616\ : InMux
    port map (
            O => \N__51436\,
            I => \N__51416\
        );

    \I__11615\ : InMux
    port map (
            O => \N__51433\,
            I => \N__51412\
        );

    \I__11614\ : CascadeMux
    port map (
            O => \N__51432\,
            I => \N__51406\
        );

    \I__11613\ : InMux
    port map (
            O => \N__51431\,
            I => \N__51401\
        );

    \I__11612\ : InMux
    port map (
            O => \N__51428\,
            I => \N__51397\
        );

    \I__11611\ : InMux
    port map (
            O => \N__51427\,
            I => \N__51394\
        );

    \I__11610\ : InMux
    port map (
            O => \N__51426\,
            I => \N__51391\
        );

    \I__11609\ : Span4Mux_v
    port map (
            O => \N__51419\,
            I => \N__51386\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__51416\,
            I => \N__51386\
        );

    \I__11607\ : InMux
    port map (
            O => \N__51415\,
            I => \N__51383\
        );

    \I__11606\ : LocalMux
    port map (
            O => \N__51412\,
            I => \N__51378\
        );

    \I__11605\ : InMux
    port map (
            O => \N__51411\,
            I => \N__51375\
        );

    \I__11604\ : InMux
    port map (
            O => \N__51410\,
            I => \N__51372\
        );

    \I__11603\ : InMux
    port map (
            O => \N__51409\,
            I => \N__51369\
        );

    \I__11602\ : InMux
    port map (
            O => \N__51406\,
            I => \N__51366\
        );

    \I__11601\ : InMux
    port map (
            O => \N__51405\,
            I => \N__51362\
        );

    \I__11600\ : InMux
    port map (
            O => \N__51404\,
            I => \N__51359\
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__51401\,
            I => \N__51356\
        );

    \I__11598\ : CascadeMux
    port map (
            O => \N__51400\,
            I => \N__51353\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__51397\,
            I => \N__51350\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__51394\,
            I => \N__51347\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__51391\,
            I => \N__51342\
        );

    \I__11594\ : Span4Mux_v
    port map (
            O => \N__51386\,
            I => \N__51342\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__51383\,
            I => \N__51339\
        );

    \I__11592\ : InMux
    port map (
            O => \N__51382\,
            I => \N__51334\
        );

    \I__11591\ : InMux
    port map (
            O => \N__51381\,
            I => \N__51334\
        );

    \I__11590\ : Span4Mux_v
    port map (
            O => \N__51378\,
            I => \N__51329\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__51375\,
            I => \N__51329\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__51372\,
            I => \N__51324\
        );

    \I__11587\ : LocalMux
    port map (
            O => \N__51369\,
            I => \N__51324\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__51366\,
            I => \N__51321\
        );

    \I__11585\ : InMux
    port map (
            O => \N__51365\,
            I => \N__51318\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__51362\,
            I => \N__51315\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__51359\,
            I => \N__51310\
        );

    \I__11582\ : Span4Mux_h
    port map (
            O => \N__51356\,
            I => \N__51310\
        );

    \I__11581\ : InMux
    port map (
            O => \N__51353\,
            I => \N__51307\
        );

    \I__11580\ : Span4Mux_h
    port map (
            O => \N__51350\,
            I => \N__51298\
        );

    \I__11579\ : Span4Mux_v
    port map (
            O => \N__51347\,
            I => \N__51298\
        );

    \I__11578\ : Span4Mux_h
    port map (
            O => \N__51342\,
            I => \N__51298\
        );

    \I__11577\ : Span4Mux_h
    port map (
            O => \N__51339\,
            I => \N__51298\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__51334\,
            I => \N__51291\
        );

    \I__11575\ : Span4Mux_v
    port map (
            O => \N__51329\,
            I => \N__51291\
        );

    \I__11574\ : Span4Mux_v
    port map (
            O => \N__51324\,
            I => \N__51291\
        );

    \I__11573\ : Span4Mux_v
    port map (
            O => \N__51321\,
            I => \N__51282\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__51318\,
            I => \N__51282\
        );

    \I__11571\ : Span4Mux_h
    port map (
            O => \N__51315\,
            I => \N__51282\
        );

    \I__11570\ : Span4Mux_v
    port map (
            O => \N__51310\,
            I => \N__51282\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__51307\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__11568\ : Odrv4
    port map (
            O => \N__51298\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__11567\ : Odrv4
    port map (
            O => \N__51291\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__11566\ : Odrv4
    port map (
            O => \N__51282\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__11565\ : InMux
    port map (
            O => \N__51273\,
            I => \N__51270\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__51270\,
            I => \N__51266\
        );

    \I__11563\ : InMux
    port map (
            O => \N__51269\,
            I => \N__51262\
        );

    \I__11562\ : Span4Mux_v
    port map (
            O => \N__51266\,
            I => \N__51259\
        );

    \I__11561\ : InMux
    port map (
            O => \N__51265\,
            I => \N__51256\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__51262\,
            I => \N__51249\
        );

    \I__11559\ : Sp12to4
    port map (
            O => \N__51259\,
            I => \N__51249\
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__51256\,
            I => \N__51249\
        );

    \I__11557\ : Odrv12
    port map (
            O => \N__51249\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__11556\ : InMux
    port map (
            O => \N__51246\,
            I => \N__51243\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__51243\,
            I => \N__51240\
        );

    \I__11554\ : Span4Mux_h
    port map (
            O => \N__51240\,
            I => \N__51237\
        );

    \I__11553\ : Span4Mux_h
    port map (
            O => \N__51237\,
            I => \N__51234\
        );

    \I__11552\ : Span4Mux_v
    port map (
            O => \N__51234\,
            I => \N__51231\
        );

    \I__11551\ : Odrv4
    port map (
            O => \N__51231\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\
        );

    \I__11550\ : CascadeMux
    port map (
            O => \N__51228\,
            I => \N__51223\
        );

    \I__11549\ : InMux
    port map (
            O => \N__51227\,
            I => \N__51220\
        );

    \I__11548\ : InMux
    port map (
            O => \N__51226\,
            I => \N__51215\
        );

    \I__11547\ : InMux
    port map (
            O => \N__51223\,
            I => \N__51215\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__51220\,
            I => \N__51210\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__51215\,
            I => \N__51210\
        );

    \I__11544\ : Span4Mux_v
    port map (
            O => \N__51210\,
            I => \N__51207\
        );

    \I__11543\ : Odrv4
    port map (
            O => \N__51207\,
            I => \pid_side.un1_pid_prereg_56\
        );

    \I__11542\ : CascadeMux
    port map (
            O => \N__51204\,
            I => \N__51201\
        );

    \I__11541\ : InMux
    port map (
            O => \N__51201\,
            I => \N__51198\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__51198\,
            I => \pid_side.error_d_reg_prev_esr_RNIO9BH1Z0Z_20\
        );

    \I__11539\ : InMux
    port map (
            O => \N__51195\,
            I => \N__51192\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__51192\,
            I => \N__51189\
        );

    \I__11537\ : Odrv4
    port map (
            O => \N__51189\,
            I => \pid_side.error_d_reg_prev_esr_RNILJFJ2Z0Z_12\
        );

    \I__11536\ : CascadeMux
    port map (
            O => \N__51186\,
            I => \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10_cascade_\
        );

    \I__11535\ : CascadeMux
    port map (
            O => \N__51183\,
            I => \N__51180\
        );

    \I__11534\ : InMux
    port map (
            O => \N__51180\,
            I => \N__51176\
        );

    \I__11533\ : InMux
    port map (
            O => \N__51179\,
            I => \N__51173\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__51176\,
            I => \N__51170\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__51173\,
            I => \pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10\
        );

    \I__11530\ : Odrv4
    port map (
            O => \N__51170\,
            I => \pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10\
        );

    \I__11529\ : CascadeMux
    port map (
            O => \N__51165\,
            I => \N__51162\
        );

    \I__11528\ : InMux
    port map (
            O => \N__51162\,
            I => \N__51159\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__51159\,
            I => \N__51155\
        );

    \I__11526\ : InMux
    port map (
            O => \N__51158\,
            I => \N__51152\
        );

    \I__11525\ : Odrv4
    port map (
            O => \N__51155\,
            I => \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11\
        );

    \I__11524\ : LocalMux
    port map (
            O => \N__51152\,
            I => \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11\
        );

    \I__11523\ : CascadeMux
    port map (
            O => \N__51147\,
            I => \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11_cascade_\
        );

    \I__11522\ : InMux
    port map (
            O => \N__51144\,
            I => \N__51138\
        );

    \I__11521\ : InMux
    port map (
            O => \N__51143\,
            I => \N__51138\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__51138\,
            I => \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10\
        );

    \I__11519\ : CascadeMux
    port map (
            O => \N__51135\,
            I => \N__51132\
        );

    \I__11518\ : InMux
    port map (
            O => \N__51132\,
            I => \N__51129\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__51129\,
            I => \N__51126\
        );

    \I__11516\ : Odrv4
    port map (
            O => \N__51126\,
            I => \pid_side.error_d_reg_prev_esr_RNIQCA21Z0Z_10\
        );

    \I__11515\ : InMux
    port map (
            O => \N__51123\,
            I => \N__51119\
        );

    \I__11514\ : CascadeMux
    port map (
            O => \N__51122\,
            I => \N__51116\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__51119\,
            I => \N__51113\
        );

    \I__11512\ : InMux
    port map (
            O => \N__51116\,
            I => \N__51110\
        );

    \I__11511\ : Odrv12
    port map (
            O => \N__51113\,
            I => \pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__51110\,
            I => \pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12\
        );

    \I__11509\ : CascadeMux
    port map (
            O => \N__51105\,
            I => \pid_side.N_1590_i_cascade_\
        );

    \I__11508\ : InMux
    port map (
            O => \N__51102\,
            I => \N__51099\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__51099\,
            I => \N__51096\
        );

    \I__11506\ : Odrv4
    port map (
            O => \N__51096\,
            I => \pid_side.error_d_reg_esr_RNIVTFJ2Z0Z_12\
        );

    \I__11505\ : InMux
    port map (
            O => \N__51093\,
            I => \N__51090\
        );

    \I__11504\ : LocalMux
    port map (
            O => \N__51090\,
            I => \N__51087\
        );

    \I__11503\ : Odrv4
    port map (
            O => \N__51087\,
            I => \pid_side.error_d_reg_prev_esr_RNI4NA21Z0Z_12\
        );

    \I__11502\ : InMux
    port map (
            O => \N__51084\,
            I => \N__51081\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__51081\,
            I => \pid_side.error_d_reg_prev_esr_RNIDP5H1Z0Z_14\
        );

    \I__11500\ : InMux
    port map (
            O => \N__51078\,
            I => \N__51075\
        );

    \I__11499\ : LocalMux
    port map (
            O => \N__51075\,
            I => \pid_side.error_d_reg_esr_RNIKMFP2Z0Z_10\
        );

    \I__11498\ : InMux
    port map (
            O => \N__51072\,
            I => \N__51069\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__51069\,
            I => \pid_side.N_1582_i\
        );

    \I__11496\ : CascadeMux
    port map (
            O => \N__51066\,
            I => \pid_side.N_1582_i_cascade_\
        );

    \I__11495\ : InMux
    port map (
            O => \N__51063\,
            I => \N__51060\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__51060\,
            I => \pid_side.error_d_reg_esr_RNI104E2Z0Z_10\
        );

    \I__11493\ : InMux
    port map (
            O => \N__51057\,
            I => \N__51054\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__51054\,
            I => \N__51051\
        );

    \I__11491\ : Odrv4
    port map (
            O => \N__51051\,
            I => \pid_side.error_d_reg_prev_esr_RNIKCB23Z0Z_13\
        );

    \I__11490\ : InMux
    port map (
            O => \N__51048\,
            I => \N__51043\
        );

    \I__11489\ : InMux
    port map (
            O => \N__51047\,
            I => \N__51038\
        );

    \I__11488\ : InMux
    port map (
            O => \N__51046\,
            I => \N__51038\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__51043\,
            I => \pid_side.un1_pid_prereg_23\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__51038\,
            I => \pid_side.un1_pid_prereg_23\
        );

    \I__11485\ : CascadeMux
    port map (
            O => \N__51033\,
            I => \N__51030\
        );

    \I__11484\ : InMux
    port map (
            O => \N__51030\,
            I => \N__51027\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__51027\,
            I => \N__51023\
        );

    \I__11482\ : InMux
    port map (
            O => \N__51026\,
            I => \N__51020\
        );

    \I__11481\ : Odrv12
    port map (
            O => \N__51023\,
            I => \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__51020\,
            I => \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13\
        );

    \I__11479\ : CascadeMux
    port map (
            O => \N__51015\,
            I => \N__51012\
        );

    \I__11478\ : InMux
    port map (
            O => \N__51012\,
            I => \N__51006\
        );

    \I__11477\ : InMux
    port map (
            O => \N__51011\,
            I => \N__51006\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__51006\,
            I => \pid_side.un1_pid_prereg_18\
        );

    \I__11475\ : CascadeMux
    port map (
            O => \N__51003\,
            I => \N__51000\
        );

    \I__11474\ : InMux
    port map (
            O => \N__51000\,
            I => \N__50997\
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__50997\,
            I => \pid_side.error_d_reg_prev_esr_RNIBAGJ2Z0Z_12\
        );

    \I__11472\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50989\
        );

    \I__11471\ : InMux
    port map (
            O => \N__50993\,
            I => \N__50984\
        );

    \I__11470\ : InMux
    port map (
            O => \N__50992\,
            I => \N__50984\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__50989\,
            I => \pid_side.un1_pid_prereg_29\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__50984\,
            I => \pid_side.un1_pid_prereg_29\
        );

    \I__11467\ : InMux
    port map (
            O => \N__50979\,
            I => \N__50973\
        );

    \I__11466\ : InMux
    port map (
            O => \N__50978\,
            I => \N__50973\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__50973\,
            I => \pid_side.error_d_reg_prevZ0Z_1\
        );

    \I__11464\ : CascadeMux
    port map (
            O => \N__50970\,
            I => \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1_cascade_\
        );

    \I__11463\ : CascadeMux
    port map (
            O => \N__50967\,
            I => \N__50963\
        );

    \I__11462\ : InMux
    port map (
            O => \N__50966\,
            I => \N__50960\
        );

    \I__11461\ : InMux
    port map (
            O => \N__50963\,
            I => \N__50957\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__50960\,
            I => \pid_side.un1_pid_prereg\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__50957\,
            I => \pid_side.un1_pid_prereg\
        );

    \I__11458\ : InMux
    port map (
            O => \N__50952\,
            I => \N__50943\
        );

    \I__11457\ : InMux
    port map (
            O => \N__50951\,
            I => \N__50943\
        );

    \I__11456\ : InMux
    port map (
            O => \N__50950\,
            I => \N__50943\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__50943\,
            I => \pid_side.error_d_reg_prevZ0Z_0\
        );

    \I__11454\ : InMux
    port map (
            O => \N__50940\,
            I => \N__50937\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__50937\,
            I => \N__50933\
        );

    \I__11452\ : InMux
    port map (
            O => \N__50936\,
            I => \N__50930\
        );

    \I__11451\ : Odrv12
    port map (
            O => \N__50933\,
            I => \pid_side.un1_pid_prereg_axb_0\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__50930\,
            I => \pid_side.un1_pid_prereg_axb_0\
        );

    \I__11449\ : InMux
    port map (
            O => \N__50925\,
            I => \N__50922\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__50922\,
            I => \pid_side.error_p_reg_esr_RNIAVKD1Z0Z_1\
        );

    \I__11447\ : CascadeMux
    port map (
            O => \N__50919\,
            I => \pid_side.un1_pid_prereg_18_cascade_\
        );

    \I__11446\ : CascadeMux
    port map (
            O => \N__50916\,
            I => \N__50913\
        );

    \I__11445\ : InMux
    port map (
            O => \N__50913\,
            I => \N__50910\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__50910\,
            I => \N__50907\
        );

    \I__11443\ : Odrv4
    port map (
            O => \N__50907\,
            I => \pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13\
        );

    \I__11442\ : CascadeMux
    port map (
            O => \N__50904\,
            I => \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13_cascade_\
        );

    \I__11441\ : InMux
    port map (
            O => \N__50901\,
            I => \N__50895\
        );

    \I__11440\ : InMux
    port map (
            O => \N__50900\,
            I => \N__50895\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__50895\,
            I => \pid_side.error_d_reg_prevZ0Z_13\
        );

    \I__11438\ : CascadeMux
    port map (
            O => \N__50892\,
            I => \N__50889\
        );

    \I__11437\ : InMux
    port map (
            O => \N__50889\,
            I => \N__50883\
        );

    \I__11436\ : InMux
    port map (
            O => \N__50888\,
            I => \N__50883\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__50883\,
            I => \N__50880\
        );

    \I__11434\ : Odrv4
    port map (
            O => \N__50880\,
            I => side_command_7
        );

    \I__11433\ : InMux
    port map (
            O => \N__50877\,
            I => \N__50874\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__50874\,
            I => \N__50871\
        );

    \I__11431\ : Odrv12
    port map (
            O => \N__50871\,
            I => \pid_front.O_7\
        );

    \I__11430\ : InMux
    port map (
            O => \N__50868\,
            I => \N__50859\
        );

    \I__11429\ : InMux
    port map (
            O => \N__50867\,
            I => \N__50859\
        );

    \I__11428\ : InMux
    port map (
            O => \N__50866\,
            I => \N__50859\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__50859\,
            I => \N__50856\
        );

    \I__11426\ : Span4Mux_h
    port map (
            O => \N__50856\,
            I => \N__50853\
        );

    \I__11425\ : Span4Mux_h
    port map (
            O => \N__50853\,
            I => \N__50850\
        );

    \I__11424\ : Odrv4
    port map (
            O => \N__50850\,
            I => \pid_front.error_d_regZ0Z_3\
        );

    \I__11423\ : CascadeMux
    port map (
            O => \N__50847\,
            I => \N__50844\
        );

    \I__11422\ : InMux
    port map (
            O => \N__50844\,
            I => \N__50841\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__50841\,
            I => \N__50838\
        );

    \I__11420\ : Span4Mux_h
    port map (
            O => \N__50838\,
            I => \N__50835\
        );

    \I__11419\ : Odrv4
    port map (
            O => \N__50835\,
            I => \pid_side.error_p_reg_esr_RNI5QI23Z0Z_5\
        );

    \I__11418\ : InMux
    port map (
            O => \N__50832\,
            I => \N__50829\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__50829\,
            I => \N__50825\
        );

    \I__11416\ : InMux
    port map (
            O => \N__50828\,
            I => \N__50822\
        );

    \I__11415\ : Odrv12
    port map (
            O => \N__50825\,
            I => \pid_side.un1_pid_prereg_axb_1\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__50822\,
            I => \pid_side.un1_pid_prereg_axb_1\
        );

    \I__11413\ : CascadeMux
    port map (
            O => \N__50817\,
            I => \pid_side.error_p_reg_esr_RNISH6JZ0Z_0_cascade_\
        );

    \I__11412\ : InMux
    port map (
            O => \N__50814\,
            I => \N__50811\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__50811\,
            I => \pid_side.error_d_reg_esr_RNIFP9R2Z0Z_1\
        );

    \I__11410\ : InMux
    port map (
            O => \N__50808\,
            I => \N__50802\
        );

    \I__11409\ : InMux
    port map (
            O => \N__50807\,
            I => \N__50802\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__50802\,
            I => \pid_side.N_1546_i\
        );

    \I__11407\ : InMux
    port map (
            O => \N__50799\,
            I => \N__50796\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__50796\,
            I => \N__50793\
        );

    \I__11405\ : Span4Mux_h
    port map (
            O => \N__50793\,
            I => \N__50790\
        );

    \I__11404\ : Span4Mux_h
    port map (
            O => \N__50790\,
            I => \N__50787\
        );

    \I__11403\ : Span4Mux_v
    port map (
            O => \N__50787\,
            I => \N__50784\
        );

    \I__11402\ : Odrv4
    port map (
            O => \N__50784\,
            I => \drone_H_disp_front_i_9\
        );

    \I__11401\ : InMux
    port map (
            O => \N__50781\,
            I => \N__50776\
        );

    \I__11400\ : InMux
    port map (
            O => \N__50780\,
            I => \N__50773\
        );

    \I__11399\ : InMux
    port map (
            O => \N__50779\,
            I => \N__50769\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__50776\,
            I => \N__50762\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__50773\,
            I => \N__50762\
        );

    \I__11396\ : InMux
    port map (
            O => \N__50772\,
            I => \N__50759\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__50769\,
            I => \N__50756\
        );

    \I__11394\ : InMux
    port map (
            O => \N__50768\,
            I => \N__50753\
        );

    \I__11393\ : InMux
    port map (
            O => \N__50767\,
            I => \N__50750\
        );

    \I__11392\ : Span4Mux_v
    port map (
            O => \N__50762\,
            I => \N__50746\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__50759\,
            I => \N__50743\
        );

    \I__11390\ : Span4Mux_h
    port map (
            O => \N__50756\,
            I => \N__50738\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__50753\,
            I => \N__50738\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__50750\,
            I => \N__50735\
        );

    \I__11387\ : InMux
    port map (
            O => \N__50749\,
            I => \N__50732\
        );

    \I__11386\ : Sp12to4
    port map (
            O => \N__50746\,
            I => \N__50728\
        );

    \I__11385\ : Span4Mux_h
    port map (
            O => \N__50743\,
            I => \N__50725\
        );

    \I__11384\ : Span4Mux_v
    port map (
            O => \N__50738\,
            I => \N__50718\
        );

    \I__11383\ : Span4Mux_h
    port map (
            O => \N__50735\,
            I => \N__50718\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__50732\,
            I => \N__50718\
        );

    \I__11381\ : InMux
    port map (
            O => \N__50731\,
            I => \N__50715\
        );

    \I__11380\ : Span12Mux_h
    port map (
            O => \N__50728\,
            I => \N__50706\
        );

    \I__11379\ : Sp12to4
    port map (
            O => \N__50725\,
            I => \N__50706\
        );

    \I__11378\ : Sp12to4
    port map (
            O => \N__50718\,
            I => \N__50706\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__50715\,
            I => \N__50706\
        );

    \I__11376\ : Odrv12
    port map (
            O => \N__50706\,
            I => uart_drone_data_1
        );

    \I__11375\ : InMux
    port map (
            O => \N__50703\,
            I => \N__50700\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__50700\,
            I => \dron_frame_decoder_1.drone_H_disp_front_9\
        );

    \I__11373\ : CEMux
    port map (
            O => \N__50697\,
            I => \N__50693\
        );

    \I__11372\ : CEMux
    port map (
            O => \N__50696\,
            I => \N__50689\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__50693\,
            I => \N__50686\
        );

    \I__11370\ : CEMux
    port map (
            O => \N__50692\,
            I => \N__50683\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__50689\,
            I => \N__50680\
        );

    \I__11368\ : Span4Mux_h
    port map (
            O => \N__50686\,
            I => \N__50677\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__50683\,
            I => \N__50674\
        );

    \I__11366\ : Sp12to4
    port map (
            O => \N__50680\,
            I => \N__50671\
        );

    \I__11365\ : Sp12to4
    port map (
            O => \N__50677\,
            I => \N__50668\
        );

    \I__11364\ : Span4Mux_h
    port map (
            O => \N__50674\,
            I => \N__50665\
        );

    \I__11363\ : Span12Mux_v
    port map (
            O => \N__50671\,
            I => \N__50662\
        );

    \I__11362\ : Span12Mux_v
    port map (
            O => \N__50668\,
            I => \N__50659\
        );

    \I__11361\ : Sp12to4
    port map (
            O => \N__50665\,
            I => \N__50656\
        );

    \I__11360\ : Odrv12
    port map (
            O => \N__50662\,
            I => \dron_frame_decoder_1.N_481_0\
        );

    \I__11359\ : Odrv12
    port map (
            O => \N__50659\,
            I => \dron_frame_decoder_1.N_481_0\
        );

    \I__11358\ : Odrv12
    port map (
            O => \N__50656\,
            I => \dron_frame_decoder_1.N_481_0\
        );

    \I__11357\ : InMux
    port map (
            O => \N__50649\,
            I => \N__50646\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__50646\,
            I => \dron_frame_decoder_1.drone_H_disp_side_4\
        );

    \I__11355\ : InMux
    port map (
            O => \N__50643\,
            I => \N__50640\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__50640\,
            I => \N__50637\
        );

    \I__11353\ : Odrv4
    port map (
            O => \N__50637\,
            I => \dron_frame_decoder_1.drone_H_disp_side_6\
        );

    \I__11352\ : InMux
    port map (
            O => \N__50634\,
            I => \N__50631\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__50631\,
            I => \N__50628\
        );

    \I__11350\ : Odrv4
    port map (
            O => \N__50628\,
            I => \dron_frame_decoder_1.drone_H_disp_side_7\
        );

    \I__11349\ : InMux
    port map (
            O => \N__50625\,
            I => \N__50619\
        );

    \I__11348\ : InMux
    port map (
            O => \N__50624\,
            I => \N__50612\
        );

    \I__11347\ : InMux
    port map (
            O => \N__50623\,
            I => \N__50612\
        );

    \I__11346\ : InMux
    port map (
            O => \N__50622\,
            I => \N__50612\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__50619\,
            I => \N__50602\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__50612\,
            I => \N__50599\
        );

    \I__11343\ : InMux
    port map (
            O => \N__50611\,
            I => \N__50596\
        );

    \I__11342\ : InMux
    port map (
            O => \N__50610\,
            I => \N__50583\
        );

    \I__11341\ : InMux
    port map (
            O => \N__50609\,
            I => \N__50583\
        );

    \I__11340\ : InMux
    port map (
            O => \N__50608\,
            I => \N__50583\
        );

    \I__11339\ : InMux
    port map (
            O => \N__50607\,
            I => \N__50583\
        );

    \I__11338\ : InMux
    port map (
            O => \N__50606\,
            I => \N__50583\
        );

    \I__11337\ : InMux
    port map (
            O => \N__50605\,
            I => \N__50583\
        );

    \I__11336\ : Span4Mux_h
    port map (
            O => \N__50602\,
            I => \N__50580\
        );

    \I__11335\ : Span4Mux_h
    port map (
            O => \N__50599\,
            I => \N__50577\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__50596\,
            I => \N__50574\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__50583\,
            I => \N__50571\
        );

    \I__11332\ : Span4Mux_h
    port map (
            O => \N__50580\,
            I => \N__50568\
        );

    \I__11331\ : Span4Mux_h
    port map (
            O => \N__50577\,
            I => \N__50565\
        );

    \I__11330\ : Span12Mux_h
    port map (
            O => \N__50574\,
            I => \N__50562\
        );

    \I__11329\ : Span12Mux_h
    port map (
            O => \N__50571\,
            I => \N__50559\
        );

    \I__11328\ : Span4Mux_v
    port map (
            O => \N__50568\,
            I => \N__50556\
        );

    \I__11327\ : Span4Mux_h
    port map (
            O => \N__50565\,
            I => \N__50553\
        );

    \I__11326\ : Odrv12
    port map (
            O => \N__50562\,
            I => \pid_front.stateZ0Z_1\
        );

    \I__11325\ : Odrv12
    port map (
            O => \N__50559\,
            I => \pid_front.stateZ0Z_1\
        );

    \I__11324\ : Odrv4
    port map (
            O => \N__50556\,
            I => \pid_front.stateZ0Z_1\
        );

    \I__11323\ : Odrv4
    port map (
            O => \N__50553\,
            I => \pid_front.stateZ0Z_1\
        );

    \I__11322\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50541\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__50541\,
            I => \N__50538\
        );

    \I__11320\ : Span4Mux_h
    port map (
            O => \N__50538\,
            I => \N__50535\
        );

    \I__11319\ : Span4Mux_h
    port map (
            O => \N__50535\,
            I => \N__50532\
        );

    \I__11318\ : Odrv4
    port map (
            O => \N__50532\,
            I => \pid_front.un1_pid_prereg_cry_0_THRU_CO\
        );

    \I__11317\ : InMux
    port map (
            O => \N__50529\,
            I => \N__50526\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__50526\,
            I => \N__50523\
        );

    \I__11315\ : Span4Mux_v
    port map (
            O => \N__50523\,
            I => \N__50520\
        );

    \I__11314\ : Span4Mux_h
    port map (
            O => \N__50520\,
            I => \N__50516\
        );

    \I__11313\ : InMux
    port map (
            O => \N__50519\,
            I => \N__50513\
        );

    \I__11312\ : Odrv4
    port map (
            O => \N__50516\,
            I => \pid_front.un1_pid_prereg_axb_1\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__50513\,
            I => \pid_front.un1_pid_prereg_axb_1\
        );

    \I__11310\ : InMux
    port map (
            O => \N__50508\,
            I => \N__50502\
        );

    \I__11309\ : CascadeMux
    port map (
            O => \N__50507\,
            I => \N__50499\
        );

    \I__11308\ : InMux
    port map (
            O => \N__50506\,
            I => \N__50494\
        );

    \I__11307\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50494\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__50502\,
            I => \N__50490\
        );

    \I__11305\ : InMux
    port map (
            O => \N__50499\,
            I => \N__50487\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__50494\,
            I => \N__50484\
        );

    \I__11303\ : InMux
    port map (
            O => \N__50493\,
            I => \N__50481\
        );

    \I__11302\ : Span4Mux_v
    port map (
            O => \N__50490\,
            I => \N__50477\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__50487\,
            I => \N__50474\
        );

    \I__11300\ : Span12Mux_v
    port map (
            O => \N__50484\,
            I => \N__50471\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__50481\,
            I => \N__50468\
        );

    \I__11298\ : InMux
    port map (
            O => \N__50480\,
            I => \N__50465\
        );

    \I__11297\ : Span4Mux_h
    port map (
            O => \N__50477\,
            I => \N__50462\
        );

    \I__11296\ : Span4Mux_v
    port map (
            O => \N__50474\,
            I => \N__50459\
        );

    \I__11295\ : Span12Mux_h
    port map (
            O => \N__50471\,
            I => \N__50454\
        );

    \I__11294\ : Span12Mux_s4_v
    port map (
            O => \N__50468\,
            I => \N__50454\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__50465\,
            I => \N__50447\
        );

    \I__11292\ : Span4Mux_h
    port map (
            O => \N__50462\,
            I => \N__50447\
        );

    \I__11291\ : Span4Mux_v
    port map (
            O => \N__50459\,
            I => \N__50447\
        );

    \I__11290\ : Odrv12
    port map (
            O => \N__50454\,
            I => \pid_front.stateZ0Z_0\
        );

    \I__11289\ : Odrv4
    port map (
            O => \N__50447\,
            I => \pid_front.stateZ0Z_0\
        );

    \I__11288\ : InMux
    port map (
            O => \N__50442\,
            I => \N__50438\
        );

    \I__11287\ : InMux
    port map (
            O => \N__50441\,
            I => \N__50435\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__50438\,
            I => \N__50431\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__50435\,
            I => \N__50428\
        );

    \I__11284\ : CascadeMux
    port map (
            O => \N__50434\,
            I => \N__50425\
        );

    \I__11283\ : Span4Mux_v
    port map (
            O => \N__50431\,
            I => \N__50420\
        );

    \I__11282\ : Span4Mux_v
    port map (
            O => \N__50428\,
            I => \N__50420\
        );

    \I__11281\ : InMux
    port map (
            O => \N__50425\,
            I => \N__50417\
        );

    \I__11280\ : Sp12to4
    port map (
            O => \N__50420\,
            I => \N__50414\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__50417\,
            I => \pid_front.pid_preregZ0Z_1\
        );

    \I__11278\ : Odrv12
    port map (
            O => \N__50414\,
            I => \pid_front.pid_preregZ0Z_1\
        );

    \I__11277\ : InMux
    port map (
            O => \N__50409\,
            I => \N__50406\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__50406\,
            I => \drone_H_disp_side_1\
        );

    \I__11275\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50399\
        );

    \I__11274\ : InMux
    port map (
            O => \N__50402\,
            I => \N__50395\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__50399\,
            I => \N__50391\
        );

    \I__11272\ : InMux
    port map (
            O => \N__50398\,
            I => \N__50388\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__50395\,
            I => \N__50385\
        );

    \I__11270\ : InMux
    port map (
            O => \N__50394\,
            I => \N__50380\
        );

    \I__11269\ : Span4Mux_v
    port map (
            O => \N__50391\,
            I => \N__50375\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__50388\,
            I => \N__50375\
        );

    \I__11267\ : Span4Mux_h
    port map (
            O => \N__50385\,
            I => \N__50372\
        );

    \I__11266\ : InMux
    port map (
            O => \N__50384\,
            I => \N__50369\
        );

    \I__11265\ : InMux
    port map (
            O => \N__50383\,
            I => \N__50366\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__50380\,
            I => \N__50363\
        );

    \I__11263\ : Span4Mux_v
    port map (
            O => \N__50375\,
            I => \N__50360\
        );

    \I__11262\ : Span4Mux_h
    port map (
            O => \N__50372\,
            I => \N__50357\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__50369\,
            I => \N__50354\
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__50366\,
            I => \N__50351\
        );

    \I__11259\ : Span12Mux_s4_h
    port map (
            O => \N__50363\,
            I => \N__50348\
        );

    \I__11258\ : Span4Mux_v
    port map (
            O => \N__50360\,
            I => \N__50345\
        );

    \I__11257\ : Span4Mux_h
    port map (
            O => \N__50357\,
            I => \N__50340\
        );

    \I__11256\ : Span4Mux_v
    port map (
            O => \N__50354\,
            I => \N__50340\
        );

    \I__11255\ : Span4Mux_v
    port map (
            O => \N__50351\,
            I => \N__50337\
        );

    \I__11254\ : Span12Mux_v
    port map (
            O => \N__50348\,
            I => \N__50333\
        );

    \I__11253\ : Span4Mux_v
    port map (
            O => \N__50345\,
            I => \N__50330\
        );

    \I__11252\ : Span4Mux_v
    port map (
            O => \N__50340\,
            I => \N__50327\
        );

    \I__11251\ : Span4Mux_v
    port map (
            O => \N__50337\,
            I => \N__50324\
        );

    \I__11250\ : InMux
    port map (
            O => \N__50336\,
            I => \N__50321\
        );

    \I__11249\ : Odrv12
    port map (
            O => \N__50333\,
            I => uart_drone_data_2
        );

    \I__11248\ : Odrv4
    port map (
            O => \N__50330\,
            I => uart_drone_data_2
        );

    \I__11247\ : Odrv4
    port map (
            O => \N__50327\,
            I => uart_drone_data_2
        );

    \I__11246\ : Odrv4
    port map (
            O => \N__50324\,
            I => uart_drone_data_2
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__50321\,
            I => uart_drone_data_2
        );

    \I__11244\ : InMux
    port map (
            O => \N__50310\,
            I => \N__50307\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__50307\,
            I => \drone_H_disp_side_2\
        );

    \I__11242\ : InMux
    port map (
            O => \N__50304\,
            I => \N__50301\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__50301\,
            I => \drone_H_disp_side_3\
        );

    \I__11240\ : CEMux
    port map (
            O => \N__50298\,
            I => \N__50294\
        );

    \I__11239\ : CEMux
    port map (
            O => \N__50297\,
            I => \N__50291\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__50294\,
            I => \N__50288\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__50291\,
            I => \N__50285\
        );

    \I__11236\ : Span4Mux_h
    port map (
            O => \N__50288\,
            I => \N__50280\
        );

    \I__11235\ : Span4Mux_v
    port map (
            O => \N__50285\,
            I => \N__50280\
        );

    \I__11234\ : Sp12to4
    port map (
            O => \N__50280\,
            I => \N__50277\
        );

    \I__11233\ : Odrv12
    port map (
            O => \N__50277\,
            I => \dron_frame_decoder_1.N_505_0\
        );

    \I__11232\ : InMux
    port map (
            O => \N__50274\,
            I => \N__50271\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__50271\,
            I => \N__50268\
        );

    \I__11230\ : Odrv12
    port map (
            O => \N__50268\,
            I => \pid_side.error_d_reg_prev_esr_RNIGJM23Z0Z_20\
        );

    \I__11229\ : InMux
    port map (
            O => \N__50265\,
            I => \N__50262\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__50262\,
            I => \N__50259\
        );

    \I__11227\ : Odrv12
    port map (
            O => \N__50259\,
            I => \pid_side.un1_pid_prereg_axb_21\
        );

    \I__11226\ : InMux
    port map (
            O => \N__50256\,
            I => \N__50253\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__50253\,
            I => \N__50250\
        );

    \I__11224\ : Span4Mux_v
    port map (
            O => \N__50250\,
            I => \N__50247\
        );

    \I__11223\ : Odrv4
    port map (
            O => \N__50247\,
            I => \ppm_encoder_1.N_286\
        );

    \I__11222\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50241\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__50241\,
            I => \N__50237\
        );

    \I__11220\ : InMux
    port map (
            O => \N__50240\,
            I => \N__50234\
        );

    \I__11219\ : Span4Mux_v
    port map (
            O => \N__50237\,
            I => \N__50230\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__50234\,
            I => \N__50227\
        );

    \I__11217\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50224\
        );

    \I__11216\ : Span4Mux_h
    port map (
            O => \N__50230\,
            I => \N__50219\
        );

    \I__11215\ : Span4Mux_v
    port map (
            O => \N__50227\,
            I => \N__50219\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__50224\,
            I => \ppm_encoder_1.aileronZ0Z_0\
        );

    \I__11213\ : Odrv4
    port map (
            O => \N__50219\,
            I => \ppm_encoder_1.aileronZ0Z_0\
        );

    \I__11212\ : InMux
    port map (
            O => \N__50214\,
            I => \N__50211\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__50211\,
            I => \N__50208\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__50208\,
            I => \N__50205\
        );

    \I__11209\ : Span4Mux_v
    port map (
            O => \N__50205\,
            I => \N__50202\
        );

    \I__11208\ : Span4Mux_v
    port map (
            O => \N__50202\,
            I => \N__50199\
        );

    \I__11207\ : Odrv4
    port map (
            O => \N__50199\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\
        );

    \I__11206\ : CascadeMux
    port map (
            O => \N__50196\,
            I => \N__50193\
        );

    \I__11205\ : InMux
    port map (
            O => \N__50193\,
            I => \N__50190\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__50190\,
            I => \N__50187\
        );

    \I__11203\ : Odrv12
    port map (
            O => \N__50187\,
            I => \pid_side.error_d_reg_prev_esr_RNIGV8H1Z0Z_19\
        );

    \I__11202\ : CascadeMux
    port map (
            O => \N__50184\,
            I => \pid_side.un1_pid_prereg_30_cascade_\
        );

    \I__11201\ : CascadeMux
    port map (
            O => \N__50181\,
            I => \N__50178\
        );

    \I__11200\ : InMux
    port map (
            O => \N__50178\,
            I => \N__50175\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__50175\,
            I => \pid_side.error_d_reg_prev_esr_RNI0PB23Z0Z_14\
        );

    \I__11198\ : InMux
    port map (
            O => \N__50172\,
            I => \N__50169\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__50169\,
            I => \pid_side.error_d_reg_prev_esr_RNI4UC23Z0Z_17\
        );

    \I__11196\ : CascadeMux
    port map (
            O => \N__50166\,
            I => \N__50163\
        );

    \I__11195\ : InMux
    port map (
            O => \N__50163\,
            I => \N__50160\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__50160\,
            I => \pid_side.error_d_reg_prev_esr_RNI5I6H1Z0Z_18\
        );

    \I__11193\ : InMux
    port map (
            O => \N__50157\,
            I => \N__50154\
        );

    \I__11192\ : LocalMux
    port map (
            O => \N__50154\,
            I => \N__50151\
        );

    \I__11191\ : Odrv4
    port map (
            O => \N__50151\,
            I => \pid_side.error_d_reg_prev_esr_RNIP56H1Z0Z_16\
        );

    \I__11190\ : CascadeMux
    port map (
            O => \N__50148\,
            I => \N__50145\
        );

    \I__11189\ : InMux
    port map (
            O => \N__50145\,
            I => \N__50139\
        );

    \I__11188\ : InMux
    port map (
            O => \N__50144\,
            I => \N__50139\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__50139\,
            I => \pid_side.error_d_reg_prevZ0Z_16\
        );

    \I__11186\ : InMux
    port map (
            O => \N__50136\,
            I => \N__50131\
        );

    \I__11185\ : InMux
    port map (
            O => \N__50135\,
            I => \N__50126\
        );

    \I__11184\ : InMux
    port map (
            O => \N__50134\,
            I => \N__50126\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__50131\,
            I => \pid_side.un1_pid_prereg_35\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__50126\,
            I => \pid_side.un1_pid_prereg_35\
        );

    \I__11181\ : CascadeMux
    port map (
            O => \N__50121\,
            I => \pid_side.un1_pid_prereg_36_cascade_\
        );

    \I__11180\ : InMux
    port map (
            O => \N__50118\,
            I => \N__50114\
        );

    \I__11179\ : InMux
    port map (
            O => \N__50117\,
            I => \N__50111\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__50114\,
            I => \pid_side.un1_pid_prereg_30\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__50111\,
            I => \pid_side.un1_pid_prereg_30\
        );

    \I__11176\ : CascadeMux
    port map (
            O => \N__50106\,
            I => \N__50103\
        );

    \I__11175\ : InMux
    port map (
            O => \N__50103\,
            I => \N__50100\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__50100\,
            I => \N__50097\
        );

    \I__11173\ : Odrv4
    port map (
            O => \N__50097\,
            I => \pid_side.error_d_reg_prev_esr_RNIC5C23Z0Z_15\
        );

    \I__11172\ : InMux
    port map (
            O => \N__50094\,
            I => \N__50091\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__50091\,
            I => \N__50088\
        );

    \I__11170\ : Odrv4
    port map (
            O => \N__50088\,
            I => \pid_side.error_d_reg_prev_esr_RNI89K23Z0Z_19\
        );

    \I__11169\ : InMux
    port map (
            O => \N__50085\,
            I => \N__50082\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__50082\,
            I => \N__50079\
        );

    \I__11167\ : Span4Mux_h
    port map (
            O => \N__50079\,
            I => \N__50076\
        );

    \I__11166\ : Odrv4
    port map (
            O => \N__50076\,
            I => \pid_side.pid_preregZ0Z_19\
        );

    \I__11165\ : InMux
    port map (
            O => \N__50073\,
            I => \pid_side.un1_pid_prereg_cry_16\
        );

    \I__11164\ : InMux
    port map (
            O => \N__50070\,
            I => \N__50067\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__50067\,
            I => \N__50064\
        );

    \I__11162\ : Odrv4
    port map (
            O => \N__50064\,
            I => \pid_side.pid_preregZ0Z_20\
        );

    \I__11161\ : InMux
    port map (
            O => \N__50061\,
            I => \pid_side.un1_pid_prereg_cry_17\
        );

    \I__11160\ : InMux
    port map (
            O => \N__50058\,
            I => \N__50055\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__50055\,
            I => \N__50052\
        );

    \I__11158\ : Odrv4
    port map (
            O => \N__50052\,
            I => \pid_side.pid_preregZ0Z_21\
        );

    \I__11157\ : InMux
    port map (
            O => \N__50049\,
            I => \pid_side.un1_pid_prereg_cry_18\
        );

    \I__11156\ : InMux
    port map (
            O => \N__50046\,
            I => \N__50043\
        );

    \I__11155\ : LocalMux
    port map (
            O => \N__50043\,
            I => \N__50040\
        );

    \I__11154\ : Span4Mux_h
    port map (
            O => \N__50040\,
            I => \N__50037\
        );

    \I__11153\ : Odrv4
    port map (
            O => \N__50037\,
            I => \pid_side.pid_preregZ0Z_22\
        );

    \I__11152\ : InMux
    port map (
            O => \N__50034\,
            I => \pid_side.un1_pid_prereg_cry_19\
        );

    \I__11151\ : InMux
    port map (
            O => \N__50031\,
            I => \pid_side.un1_pid_prereg_cry_20\
        );

    \I__11150\ : CascadeMux
    port map (
            O => \N__50028\,
            I => \N__50025\
        );

    \I__11149\ : InMux
    port map (
            O => \N__50025\,
            I => \N__50021\
        );

    \I__11148\ : InMux
    port map (
            O => \N__50024\,
            I => \N__50017\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__50021\,
            I => \N__50011\
        );

    \I__11146\ : InMux
    port map (
            O => \N__50020\,
            I => \N__50008\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__50017\,
            I => \N__50005\
        );

    \I__11144\ : InMux
    port map (
            O => \N__50016\,
            I => \N__49998\
        );

    \I__11143\ : InMux
    port map (
            O => \N__50015\,
            I => \N__49998\
        );

    \I__11142\ : InMux
    port map (
            O => \N__50014\,
            I => \N__49998\
        );

    \I__11141\ : Span4Mux_v
    port map (
            O => \N__50011\,
            I => \N__49993\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__50008\,
            I => \N__49993\
        );

    \I__11139\ : Span4Mux_h
    port map (
            O => \N__50005\,
            I => \N__49990\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__49998\,
            I => \N__49987\
        );

    \I__11137\ : Odrv4
    port map (
            O => \N__49993\,
            I => \pid_side.pid_preregZ0Z_23\
        );

    \I__11136\ : Odrv4
    port map (
            O => \N__49990\,
            I => \pid_side.pid_preregZ0Z_23\
        );

    \I__11135\ : Odrv12
    port map (
            O => \N__49987\,
            I => \pid_side.pid_preregZ0Z_23\
        );

    \I__11134\ : InMux
    port map (
            O => \N__49980\,
            I => \N__49977\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__49977\,
            I => \pid_side.error_d_reg_prev_esr_RNILHF23Z0Z_18\
        );

    \I__11132\ : InMux
    port map (
            O => \N__49974\,
            I => \N__49971\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__49971\,
            I => \pid_side.error_d_reg_prev_esr_RNIJV5H1Z0Z_15\
        );

    \I__11130\ : InMux
    port map (
            O => \N__49968\,
            I => \N__49962\
        );

    \I__11129\ : InMux
    port map (
            O => \N__49967\,
            I => \N__49959\
        );

    \I__11128\ : InMux
    port map (
            O => \N__49966\,
            I => \N__49956\
        );

    \I__11127\ : InMux
    port map (
            O => \N__49965\,
            I => \N__49953\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__49962\,
            I => \N__49950\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__49959\,
            I => \N__49947\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__49956\,
            I => \N__49942\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__49953\,
            I => \N__49942\
        );

    \I__11122\ : Span4Mux_h
    port map (
            O => \N__49950\,
            I => \N__49939\
        );

    \I__11121\ : Odrv12
    port map (
            O => \N__49947\,
            I => \pid_side.pid_preregZ0Z_10\
        );

    \I__11120\ : Odrv4
    port map (
            O => \N__49942\,
            I => \pid_side.pid_preregZ0Z_10\
        );

    \I__11119\ : Odrv4
    port map (
            O => \N__49939\,
            I => \pid_side.pid_preregZ0Z_10\
        );

    \I__11118\ : InMux
    port map (
            O => \N__49932\,
            I => \pid_side.un1_pid_prereg_cry_7\
        );

    \I__11117\ : InMux
    port map (
            O => \N__49929\,
            I => \N__49923\
        );

    \I__11116\ : InMux
    port map (
            O => \N__49928\,
            I => \N__49920\
        );

    \I__11115\ : InMux
    port map (
            O => \N__49927\,
            I => \N__49917\
        );

    \I__11114\ : InMux
    port map (
            O => \N__49926\,
            I => \N__49914\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__49923\,
            I => \N__49911\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__49920\,
            I => \N__49904\
        );

    \I__11111\ : LocalMux
    port map (
            O => \N__49917\,
            I => \N__49904\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__49914\,
            I => \N__49904\
        );

    \I__11109\ : Span4Mux_h
    port map (
            O => \N__49911\,
            I => \N__49901\
        );

    \I__11108\ : Odrv12
    port map (
            O => \N__49904\,
            I => \pid_side.pid_preregZ0Z_11\
        );

    \I__11107\ : Odrv4
    port map (
            O => \N__49901\,
            I => \pid_side.pid_preregZ0Z_11\
        );

    \I__11106\ : InMux
    port map (
            O => \N__49896\,
            I => \pid_side.un1_pid_prereg_cry_8\
        );

    \I__11105\ : CascadeMux
    port map (
            O => \N__49893\,
            I => \N__49889\
        );

    \I__11104\ : InMux
    port map (
            O => \N__49892\,
            I => \N__49886\
        );

    \I__11103\ : InMux
    port map (
            O => \N__49889\,
            I => \N__49883\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__49886\,
            I => \N__49876\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__49883\,
            I => \N__49876\
        );

    \I__11100\ : InMux
    port map (
            O => \N__49882\,
            I => \N__49871\
        );

    \I__11099\ : InMux
    port map (
            O => \N__49881\,
            I => \N__49871\
        );

    \I__11098\ : Span4Mux_v
    port map (
            O => \N__49876\,
            I => \N__49868\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__49871\,
            I => \N__49865\
        );

    \I__11096\ : Odrv4
    port map (
            O => \N__49868\,
            I => \pid_side.pid_preregZ0Z_12\
        );

    \I__11095\ : Odrv4
    port map (
            O => \N__49865\,
            I => \pid_side.pid_preregZ0Z_12\
        );

    \I__11094\ : InMux
    port map (
            O => \N__49860\,
            I => \pid_side.un1_pid_prereg_cry_9\
        );

    \I__11093\ : InMux
    port map (
            O => \N__49857\,
            I => \N__49851\
        );

    \I__11092\ : InMux
    port map (
            O => \N__49856\,
            I => \N__49848\
        );

    \I__11091\ : InMux
    port map (
            O => \N__49855\,
            I => \N__49843\
        );

    \I__11090\ : InMux
    port map (
            O => \N__49854\,
            I => \N__49843\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__49851\,
            I => \N__49835\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__49848\,
            I => \N__49835\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__49843\,
            I => \N__49835\
        );

    \I__11086\ : InMux
    port map (
            O => \N__49842\,
            I => \N__49832\
        );

    \I__11085\ : Span4Mux_v
    port map (
            O => \N__49835\,
            I => \N__49827\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__49832\,
            I => \N__49827\
        );

    \I__11083\ : Odrv4
    port map (
            O => \N__49827\,
            I => \pid_side.pid_preregZ0Z_13\
        );

    \I__11082\ : InMux
    port map (
            O => \N__49824\,
            I => \pid_side.un1_pid_prereg_cry_10\
        );

    \I__11081\ : InMux
    port map (
            O => \N__49821\,
            I => \N__49818\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__49818\,
            I => \N__49815\
        );

    \I__11079\ : Span4Mux_h
    port map (
            O => \N__49815\,
            I => \N__49812\
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__49812\,
            I => \pid_side.pid_preregZ0Z_14\
        );

    \I__11077\ : InMux
    port map (
            O => \N__49809\,
            I => \pid_side.un1_pid_prereg_cry_11\
        );

    \I__11076\ : InMux
    port map (
            O => \N__49806\,
            I => \N__49803\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__49803\,
            I => \N__49800\
        );

    \I__11074\ : Odrv4
    port map (
            O => \N__49800\,
            I => \pid_side.pid_preregZ0Z_15\
        );

    \I__11073\ : InMux
    port map (
            O => \N__49797\,
            I => \pid_side.un1_pid_prereg_cry_12\
        );

    \I__11072\ : InMux
    port map (
            O => \N__49794\,
            I => \N__49791\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__49791\,
            I => \N__49788\
        );

    \I__11070\ : Odrv4
    port map (
            O => \N__49788\,
            I => \pid_side.pid_preregZ0Z_16\
        );

    \I__11069\ : InMux
    port map (
            O => \N__49785\,
            I => \bfn_20_11_0_\
        );

    \I__11068\ : InMux
    port map (
            O => \N__49782\,
            I => \N__49779\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__49779\,
            I => \N__49776\
        );

    \I__11066\ : Odrv4
    port map (
            O => \N__49776\,
            I => \pid_side.pid_preregZ0Z_17\
        );

    \I__11065\ : InMux
    port map (
            O => \N__49773\,
            I => \pid_side.un1_pid_prereg_cry_14\
        );

    \I__11064\ : CascadeMux
    port map (
            O => \N__49770\,
            I => \N__49767\
        );

    \I__11063\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49764\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__49764\,
            I => \N__49761\
        );

    \I__11061\ : Odrv4
    port map (
            O => \N__49761\,
            I => \pid_side.pid_preregZ0Z_18\
        );

    \I__11060\ : InMux
    port map (
            O => \N__49758\,
            I => \pid_side.un1_pid_prereg_cry_15\
        );

    \I__11059\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49752\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__49752\,
            I => \N__49749\
        );

    \I__11057\ : Span4Mux_v
    port map (
            O => \N__49749\,
            I => \N__49745\
        );

    \I__11056\ : InMux
    port map (
            O => \N__49748\,
            I => \N__49742\
        );

    \I__11055\ : Span4Mux_h
    port map (
            O => \N__49745\,
            I => \N__49739\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__49742\,
            I => \N__49736\
        );

    \I__11053\ : Odrv4
    port map (
            O => \N__49739\,
            I => \pid_side.pid_preregZ0Z_2\
        );

    \I__11052\ : Odrv4
    port map (
            O => \N__49736\,
            I => \pid_side.pid_preregZ0Z_2\
        );

    \I__11051\ : InMux
    port map (
            O => \N__49731\,
            I => \pid_side.un1_pid_prereg_cry_1\
        );

    \I__11050\ : InMux
    port map (
            O => \N__49728\,
            I => \N__49725\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__49725\,
            I => \N__49721\
        );

    \I__11048\ : CascadeMux
    port map (
            O => \N__49724\,
            I => \N__49718\
        );

    \I__11047\ : Span4Mux_v
    port map (
            O => \N__49721\,
            I => \N__49715\
        );

    \I__11046\ : InMux
    port map (
            O => \N__49718\,
            I => \N__49712\
        );

    \I__11045\ : Span4Mux_h
    port map (
            O => \N__49715\,
            I => \N__49709\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__49712\,
            I => \N__49706\
        );

    \I__11043\ : Odrv4
    port map (
            O => \N__49709\,
            I => \pid_side.pid_preregZ0Z_3\
        );

    \I__11042\ : Odrv4
    port map (
            O => \N__49706\,
            I => \pid_side.pid_preregZ0Z_3\
        );

    \I__11041\ : InMux
    port map (
            O => \N__49701\,
            I => \pid_side.un1_pid_prereg_cry_0_0\
        );

    \I__11040\ : InMux
    port map (
            O => \N__49698\,
            I => \N__49691\
        );

    \I__11039\ : CascadeMux
    port map (
            O => \N__49697\,
            I => \N__49688\
        );

    \I__11038\ : CascadeMux
    port map (
            O => \N__49696\,
            I => \N__49685\
        );

    \I__11037\ : CascadeMux
    port map (
            O => \N__49695\,
            I => \N__49682\
        );

    \I__11036\ : CascadeMux
    port map (
            O => \N__49694\,
            I => \N__49678\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__49691\,
            I => \N__49675\
        );

    \I__11034\ : InMux
    port map (
            O => \N__49688\,
            I => \N__49672\
        );

    \I__11033\ : InMux
    port map (
            O => \N__49685\,
            I => \N__49665\
        );

    \I__11032\ : InMux
    port map (
            O => \N__49682\,
            I => \N__49665\
        );

    \I__11031\ : InMux
    port map (
            O => \N__49681\,
            I => \N__49665\
        );

    \I__11030\ : InMux
    port map (
            O => \N__49678\,
            I => \N__49661\
        );

    \I__11029\ : Span4Mux_h
    port map (
            O => \N__49675\,
            I => \N__49656\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__49672\,
            I => \N__49656\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__49665\,
            I => \N__49653\
        );

    \I__11026\ : InMux
    port map (
            O => \N__49664\,
            I => \N__49650\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__49661\,
            I => \N__49647\
        );

    \I__11024\ : Span4Mux_v
    port map (
            O => \N__49656\,
            I => \N__49642\
        );

    \I__11023\ : Span4Mux_v
    port map (
            O => \N__49653\,
            I => \N__49642\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__49650\,
            I => \N__49639\
        );

    \I__11021\ : Span4Mux_v
    port map (
            O => \N__49647\,
            I => \N__49636\
        );

    \I__11020\ : Span4Mux_h
    port map (
            O => \N__49642\,
            I => \N__49633\
        );

    \I__11019\ : Span4Mux_v
    port map (
            O => \N__49639\,
            I => \N__49628\
        );

    \I__11018\ : Span4Mux_h
    port map (
            O => \N__49636\,
            I => \N__49628\
        );

    \I__11017\ : Odrv4
    port map (
            O => \N__49633\,
            I => \pid_side.pid_preregZ0Z_4\
        );

    \I__11016\ : Odrv4
    port map (
            O => \N__49628\,
            I => \pid_side.pid_preregZ0Z_4\
        );

    \I__11015\ : InMux
    port map (
            O => \N__49623\,
            I => \pid_side.un1_pid_prereg_cry_1_0\
        );

    \I__11014\ : CascadeMux
    port map (
            O => \N__49620\,
            I => \N__49615\
        );

    \I__11013\ : CascadeMux
    port map (
            O => \N__49619\,
            I => \N__49612\
        );

    \I__11012\ : CascadeMux
    port map (
            O => \N__49618\,
            I => \N__49608\
        );

    \I__11011\ : InMux
    port map (
            O => \N__49615\,
            I => \N__49605\
        );

    \I__11010\ : InMux
    port map (
            O => \N__49612\,
            I => \N__49602\
        );

    \I__11009\ : InMux
    port map (
            O => \N__49611\,
            I => \N__49599\
        );

    \I__11008\ : InMux
    port map (
            O => \N__49608\,
            I => \N__49596\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__49605\,
            I => \N__49593\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__49602\,
            I => \N__49590\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__49599\,
            I => \N__49585\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__49596\,
            I => \N__49585\
        );

    \I__11003\ : Span4Mux_v
    port map (
            O => \N__49593\,
            I => \N__49580\
        );

    \I__11002\ : Span4Mux_v
    port map (
            O => \N__49590\,
            I => \N__49580\
        );

    \I__11001\ : Span4Mux_v
    port map (
            O => \N__49585\,
            I => \N__49577\
        );

    \I__11000\ : Odrv4
    port map (
            O => \N__49580\,
            I => \pid_side.pid_preregZ0Z_5\
        );

    \I__10999\ : Odrv4
    port map (
            O => \N__49577\,
            I => \pid_side.pid_preregZ0Z_5\
        );

    \I__10998\ : InMux
    port map (
            O => \N__49572\,
            I => \pid_side.un1_pid_prereg_cry_2\
        );

    \I__10997\ : CascadeMux
    port map (
            O => \N__49569\,
            I => \N__49565\
        );

    \I__10996\ : InMux
    port map (
            O => \N__49568\,
            I => \N__49561\
        );

    \I__10995\ : InMux
    port map (
            O => \N__49565\,
            I => \N__49556\
        );

    \I__10994\ : InMux
    port map (
            O => \N__49564\,
            I => \N__49556\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__49561\,
            I => \N__49551\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__49556\,
            I => \N__49551\
        );

    \I__10991\ : Span4Mux_h
    port map (
            O => \N__49551\,
            I => \N__49548\
        );

    \I__10990\ : Odrv4
    port map (
            O => \N__49548\,
            I => \pid_side.pid_preregZ0Z_6\
        );

    \I__10989\ : InMux
    port map (
            O => \N__49545\,
            I => \pid_side.un1_pid_prereg_cry_3\
        );

    \I__10988\ : InMux
    port map (
            O => \N__49542\,
            I => \N__49538\
        );

    \I__10987\ : CascadeMux
    port map (
            O => \N__49541\,
            I => \N__49534\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__49538\,
            I => \N__49531\
        );

    \I__10985\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49528\
        );

    \I__10984\ : InMux
    port map (
            O => \N__49534\,
            I => \N__49525\
        );

    \I__10983\ : Span4Mux_h
    port map (
            O => \N__49531\,
            I => \N__49518\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__49528\,
            I => \N__49518\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__49525\,
            I => \N__49518\
        );

    \I__10980\ : Span4Mux_h
    port map (
            O => \N__49518\,
            I => \N__49515\
        );

    \I__10979\ : Odrv4
    port map (
            O => \N__49515\,
            I => \pid_side.pid_preregZ0Z_7\
        );

    \I__10978\ : InMux
    port map (
            O => \N__49512\,
            I => \pid_side.un1_pid_prereg_cry_4\
        );

    \I__10977\ : InMux
    port map (
            O => \N__49509\,
            I => \N__49504\
        );

    \I__10976\ : InMux
    port map (
            O => \N__49508\,
            I => \N__49499\
        );

    \I__10975\ : InMux
    port map (
            O => \N__49507\,
            I => \N__49499\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__49504\,
            I => \N__49494\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__49499\,
            I => \N__49494\
        );

    \I__10972\ : Odrv12
    port map (
            O => \N__49494\,
            I => \pid_side.pid_preregZ0Z_8\
        );

    \I__10971\ : InMux
    port map (
            O => \N__49491\,
            I => \bfn_20_10_0_\
        );

    \I__10970\ : InMux
    port map (
            O => \N__49488\,
            I => \N__49483\
        );

    \I__10969\ : InMux
    port map (
            O => \N__49487\,
            I => \N__49480\
        );

    \I__10968\ : InMux
    port map (
            O => \N__49486\,
            I => \N__49477\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__49483\,
            I => \N__49470\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__49480\,
            I => \N__49470\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__49477\,
            I => \N__49470\
        );

    \I__10964\ : Span4Mux_h
    port map (
            O => \N__49470\,
            I => \N__49467\
        );

    \I__10963\ : Odrv4
    port map (
            O => \N__49467\,
            I => \pid_side.pid_preregZ0Z_9\
        );

    \I__10962\ : InMux
    port map (
            O => \N__49464\,
            I => \pid_side.un1_pid_prereg_cry_6\
        );

    \I__10961\ : InMux
    port map (
            O => \N__49461\,
            I => \N__49457\
        );

    \I__10960\ : InMux
    port map (
            O => \N__49460\,
            I => \N__49454\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__49457\,
            I => \N__49451\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__49454\,
            I => \N__49448\
        );

    \I__10957\ : Span4Mux_v
    port map (
            O => \N__49451\,
            I => \N__49445\
        );

    \I__10956\ : Span4Mux_v
    port map (
            O => \N__49448\,
            I => \N__49442\
        );

    \I__10955\ : Sp12to4
    port map (
            O => \N__49445\,
            I => \N__49439\
        );

    \I__10954\ : Span4Mux_h
    port map (
            O => \N__49442\,
            I => \N__49436\
        );

    \I__10953\ : Odrv12
    port map (
            O => \N__49439\,
            I => \pid_front.un1_pid_prereg_axb_0\
        );

    \I__10952\ : Odrv4
    port map (
            O => \N__49436\,
            I => \pid_front.un1_pid_prereg_axb_0\
        );

    \I__10951\ : InMux
    port map (
            O => \N__49431\,
            I => \N__49428\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__49428\,
            I => \N__49424\
        );

    \I__10949\ : InMux
    port map (
            O => \N__49427\,
            I => \N__49420\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__49424\,
            I => \N__49417\
        );

    \I__10947\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49414\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__49420\,
            I => \N__49411\
        );

    \I__10945\ : Odrv4
    port map (
            O => \N__49417\,
            I => \pid_front.pid_preregZ0Z_0\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__49414\,
            I => \pid_front.pid_preregZ0Z_0\
        );

    \I__10943\ : Odrv12
    port map (
            O => \N__49411\,
            I => \pid_front.pid_preregZ0Z_0\
        );

    \I__10942\ : CascadeMux
    port map (
            O => \N__49404\,
            I => \N__49401\
        );

    \I__10941\ : InMux
    port map (
            O => \N__49401\,
            I => \N__49397\
        );

    \I__10940\ : InMux
    port map (
            O => \N__49400\,
            I => \N__49394\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__49397\,
            I => \N__49389\
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__49394\,
            I => \N__49389\
        );

    \I__10937\ : Span4Mux_v
    port map (
            O => \N__49389\,
            I => \N__49386\
        );

    \I__10936\ : Span4Mux_h
    port map (
            O => \N__49386\,
            I => \N__49383\
        );

    \I__10935\ : Span4Mux_h
    port map (
            O => \N__49383\,
            I => \N__49380\
        );

    \I__10934\ : Odrv4
    port map (
            O => \N__49380\,
            I => \pid_front.error_d_reg_prevZ0Z_18\
        );

    \I__10933\ : CEMux
    port map (
            O => \N__49377\,
            I => \N__49317\
        );

    \I__10932\ : CEMux
    port map (
            O => \N__49376\,
            I => \N__49317\
        );

    \I__10931\ : CEMux
    port map (
            O => \N__49375\,
            I => \N__49317\
        );

    \I__10930\ : CEMux
    port map (
            O => \N__49374\,
            I => \N__49317\
        );

    \I__10929\ : CEMux
    port map (
            O => \N__49373\,
            I => \N__49317\
        );

    \I__10928\ : CEMux
    port map (
            O => \N__49372\,
            I => \N__49317\
        );

    \I__10927\ : CEMux
    port map (
            O => \N__49371\,
            I => \N__49317\
        );

    \I__10926\ : CEMux
    port map (
            O => \N__49370\,
            I => \N__49317\
        );

    \I__10925\ : CEMux
    port map (
            O => \N__49369\,
            I => \N__49317\
        );

    \I__10924\ : CEMux
    port map (
            O => \N__49368\,
            I => \N__49317\
        );

    \I__10923\ : CEMux
    port map (
            O => \N__49367\,
            I => \N__49317\
        );

    \I__10922\ : CEMux
    port map (
            O => \N__49366\,
            I => \N__49317\
        );

    \I__10921\ : CEMux
    port map (
            O => \N__49365\,
            I => \N__49317\
        );

    \I__10920\ : CEMux
    port map (
            O => \N__49364\,
            I => \N__49317\
        );

    \I__10919\ : CEMux
    port map (
            O => \N__49363\,
            I => \N__49317\
        );

    \I__10918\ : CEMux
    port map (
            O => \N__49362\,
            I => \N__49317\
        );

    \I__10917\ : CEMux
    port map (
            O => \N__49361\,
            I => \N__49317\
        );

    \I__10916\ : CEMux
    port map (
            O => \N__49360\,
            I => \N__49317\
        );

    \I__10915\ : CEMux
    port map (
            O => \N__49359\,
            I => \N__49317\
        );

    \I__10914\ : CEMux
    port map (
            O => \N__49358\,
            I => \N__49317\
        );

    \I__10913\ : GlobalMux
    port map (
            O => \N__49317\,
            I => \N__49314\
        );

    \I__10912\ : gio2CtrlBuf
    port map (
            O => \N__49314\,
            I => \pid_front.state_0_g_0\
        );

    \I__10911\ : InMux
    port map (
            O => \N__49311\,
            I => \N__49308\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__49308\,
            I => \N__49305\
        );

    \I__10909\ : Odrv12
    port map (
            O => \N__49305\,
            I => \pid_front.O_6\
        );

    \I__10908\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49296\
        );

    \I__10907\ : InMux
    port map (
            O => \N__49301\,
            I => \N__49296\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__49296\,
            I => \N__49292\
        );

    \I__10905\ : InMux
    port map (
            O => \N__49295\,
            I => \N__49289\
        );

    \I__10904\ : Span4Mux_h
    port map (
            O => \N__49292\,
            I => \N__49286\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__49289\,
            I => \N__49283\
        );

    \I__10902\ : Span4Mux_h
    port map (
            O => \N__49286\,
            I => \N__49280\
        );

    \I__10901\ : Span12Mux_v
    port map (
            O => \N__49283\,
            I => \N__49277\
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__49280\,
            I => \pid_front.error_d_regZ0Z_2\
        );

    \I__10899\ : Odrv12
    port map (
            O => \N__49277\,
            I => \pid_front.error_d_regZ0Z_2\
        );

    \I__10898\ : IoInMux
    port map (
            O => \N__49272\,
            I => \N__49269\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__49269\,
            I => \GB_BUFFER_reset_system_g_THRU_CO\
        );

    \I__10896\ : InMux
    port map (
            O => \N__49266\,
            I => \N__49263\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__49263\,
            I => \N__49260\
        );

    \I__10894\ : Odrv4
    port map (
            O => \N__49260\,
            I => \pid_side.un1_pid_prereg_cry_0_THRU_CO\
        );

    \I__10893\ : InMux
    port map (
            O => \N__49257\,
            I => \pid_side.un1_pid_prereg_cry_0\
        );

    \I__10892\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49251\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__49251\,
            I => \N__49248\
        );

    \I__10890\ : Odrv4
    port map (
            O => \N__49248\,
            I => \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13\
        );

    \I__10889\ : CascadeMux
    port map (
            O => \N__49245\,
            I => \N__49242\
        );

    \I__10888\ : InMux
    port map (
            O => \N__49242\,
            I => \N__49239\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__49239\,
            I => \N__49236\
        );

    \I__10886\ : Odrv4
    port map (
            O => \N__49236\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02\
        );

    \I__10885\ : InMux
    port map (
            O => \N__49233\,
            I => \N__49230\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__49230\,
            I => \N__49227\
        );

    \I__10883\ : Span4Mux_h
    port map (
            O => \N__49227\,
            I => \N__49224\
        );

    \I__10882\ : Odrv4
    port map (
            O => \N__49224\,
            I => \ppm_encoder_1.un1_init_pulses_11_13\
        );

    \I__10881\ : InMux
    port map (
            O => \N__49221\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_12\
        );

    \I__10880\ : InMux
    port map (
            O => \N__49218\,
            I => \N__49215\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__49215\,
            I => \N__49212\
        );

    \I__10878\ : Span4Mux_h
    port map (
            O => \N__49212\,
            I => \N__49209\
        );

    \I__10877\ : Odrv4
    port map (
            O => \N__49209\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__10876\ : InMux
    port map (
            O => \N__49206\,
            I => \N__49203\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__49203\,
            I => \N__49200\
        );

    \I__10874\ : Span4Mux_v
    port map (
            O => \N__49200\,
            I => \N__49197\
        );

    \I__10873\ : Odrv4
    port map (
            O => \N__49197\,
            I => \ppm_encoder_1.un1_init_pulses_11_14\
        );

    \I__10872\ : InMux
    port map (
            O => \N__49194\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13\
        );

    \I__10871\ : InMux
    port map (
            O => \N__49191\,
            I => \N__49188\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__49188\,
            I => \N__49185\
        );

    \I__10869\ : Odrv12
    port map (
            O => \N__49185\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_15\
        );

    \I__10868\ : InMux
    port map (
            O => \N__49182\,
            I => \N__49179\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__49179\,
            I => \N__49176\
        );

    \I__10866\ : Span4Mux_v
    port map (
            O => \N__49176\,
            I => \N__49173\
        );

    \I__10865\ : Odrv4
    port map (
            O => \N__49173\,
            I => \ppm_encoder_1.un1_init_pulses_11_15\
        );

    \I__10864\ : InMux
    port map (
            O => \N__49170\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_14\
        );

    \I__10863\ : InMux
    port map (
            O => \N__49167\,
            I => \N__49164\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__49164\,
            I => \N__49161\
        );

    \I__10861\ : Span4Mux_h
    port map (
            O => \N__49161\,
            I => \N__49158\
        );

    \I__10860\ : Odrv4
    port map (
            O => \N__49158\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_16\
        );

    \I__10859\ : InMux
    port map (
            O => \N__49155\,
            I => \N__49152\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__49152\,
            I => \N__49149\
        );

    \I__10857\ : Span4Mux_v
    port map (
            O => \N__49149\,
            I => \N__49146\
        );

    \I__10856\ : Odrv4
    port map (
            O => \N__49146\,
            I => \ppm_encoder_1.un1_init_pulses_11_16\
        );

    \I__10855\ : InMux
    port map (
            O => \N__49143\,
            I => \bfn_18_17_0_\
        );

    \I__10854\ : InMux
    port map (
            O => \N__49140\,
            I => \N__49137\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__49137\,
            I => \N__49134\
        );

    \I__10852\ : Span4Mux_h
    port map (
            O => \N__49134\,
            I => \N__49131\
        );

    \I__10851\ : Odrv4
    port map (
            O => \N__49131\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_17\
        );

    \I__10850\ : InMux
    port map (
            O => \N__49128\,
            I => \N__49125\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__49125\,
            I => \N__49122\
        );

    \I__10848\ : Span4Mux_h
    port map (
            O => \N__49122\,
            I => \N__49119\
        );

    \I__10847\ : Odrv4
    port map (
            O => \N__49119\,
            I => \ppm_encoder_1.un1_init_pulses_11_17\
        );

    \I__10846\ : InMux
    port map (
            O => \N__49116\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_16\
        );

    \I__10845\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49109\
        );

    \I__10844\ : InMux
    port map (
            O => \N__49112\,
            I => \N__49106\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__49109\,
            I => \N__49102\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__49106\,
            I => \N__49099\
        );

    \I__10841\ : CascadeMux
    port map (
            O => \N__49105\,
            I => \N__49096\
        );

    \I__10840\ : Span4Mux_v
    port map (
            O => \N__49102\,
            I => \N__49091\
        );

    \I__10839\ : Span4Mux_h
    port map (
            O => \N__49099\,
            I => \N__49091\
        );

    \I__10838\ : InMux
    port map (
            O => \N__49096\,
            I => \N__49088\
        );

    \I__10837\ : Odrv4
    port map (
            O => \N__49091\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__49088\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__10835\ : InMux
    port map (
            O => \N__49083\,
            I => \N__49070\
        );

    \I__10834\ : CascadeMux
    port map (
            O => \N__49082\,
            I => \N__49062\
        );

    \I__10833\ : InMux
    port map (
            O => \N__49081\,
            I => \N__49053\
        );

    \I__10832\ : InMux
    port map (
            O => \N__49080\,
            I => \N__49053\
        );

    \I__10831\ : InMux
    port map (
            O => \N__49079\,
            I => \N__49053\
        );

    \I__10830\ : InMux
    port map (
            O => \N__49078\,
            I => \N__49044\
        );

    \I__10829\ : InMux
    port map (
            O => \N__49077\,
            I => \N__49044\
        );

    \I__10828\ : InMux
    port map (
            O => \N__49076\,
            I => \N__49044\
        );

    \I__10827\ : InMux
    port map (
            O => \N__49075\,
            I => \N__49044\
        );

    \I__10826\ : InMux
    port map (
            O => \N__49074\,
            I => \N__49040\
        );

    \I__10825\ : InMux
    port map (
            O => \N__49073\,
            I => \N__49037\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__49070\,
            I => \N__49034\
        );

    \I__10823\ : InMux
    port map (
            O => \N__49069\,
            I => \N__49027\
        );

    \I__10822\ : InMux
    port map (
            O => \N__49068\,
            I => \N__49027\
        );

    \I__10821\ : InMux
    port map (
            O => \N__49067\,
            I => \N__49027\
        );

    \I__10820\ : CascadeMux
    port map (
            O => \N__49066\,
            I => \N__49018\
        );

    \I__10819\ : CascadeMux
    port map (
            O => \N__49065\,
            I => \N__49015\
        );

    \I__10818\ : InMux
    port map (
            O => \N__49062\,
            I => \N__49008\
        );

    \I__10817\ : InMux
    port map (
            O => \N__49061\,
            I => \N__49008\
        );

    \I__10816\ : InMux
    port map (
            O => \N__49060\,
            I => \N__49005\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__49053\,
            I => \N__49000\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__49044\,
            I => \N__49000\
        );

    \I__10813\ : CascadeMux
    port map (
            O => \N__49043\,
            I => \N__48991\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__49040\,
            I => \N__48977\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__49037\,
            I => \N__48977\
        );

    \I__10810\ : Span4Mux_v
    port map (
            O => \N__49034\,
            I => \N__48977\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__49027\,
            I => \N__48977\
        );

    \I__10808\ : InMux
    port map (
            O => \N__49026\,
            I => \N__48972\
        );

    \I__10807\ : InMux
    port map (
            O => \N__49025\,
            I => \N__48972\
        );

    \I__10806\ : InMux
    port map (
            O => \N__49024\,
            I => \N__48967\
        );

    \I__10805\ : InMux
    port map (
            O => \N__49023\,
            I => \N__48967\
        );

    \I__10804\ : InMux
    port map (
            O => \N__49022\,
            I => \N__48956\
        );

    \I__10803\ : InMux
    port map (
            O => \N__49021\,
            I => \N__48956\
        );

    \I__10802\ : InMux
    port map (
            O => \N__49018\,
            I => \N__48956\
        );

    \I__10801\ : InMux
    port map (
            O => \N__49015\,
            I => \N__48956\
        );

    \I__10800\ : InMux
    port map (
            O => \N__49014\,
            I => \N__48956\
        );

    \I__10799\ : InMux
    port map (
            O => \N__49013\,
            I => \N__48953\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__49008\,
            I => \N__48950\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__49005\,
            I => \N__48945\
        );

    \I__10796\ : Span4Mux_h
    port map (
            O => \N__49000\,
            I => \N__48945\
        );

    \I__10795\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48936\
        );

    \I__10794\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48936\
        );

    \I__10793\ : InMux
    port map (
            O => \N__48997\,
            I => \N__48936\
        );

    \I__10792\ : InMux
    port map (
            O => \N__48996\,
            I => \N__48936\
        );

    \I__10791\ : CascadeMux
    port map (
            O => \N__48995\,
            I => \N__48932\
        );

    \I__10790\ : InMux
    port map (
            O => \N__48994\,
            I => \N__48928\
        );

    \I__10789\ : InMux
    port map (
            O => \N__48991\,
            I => \N__48923\
        );

    \I__10788\ : InMux
    port map (
            O => \N__48990\,
            I => \N__48923\
        );

    \I__10787\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48914\
        );

    \I__10786\ : InMux
    port map (
            O => \N__48988\,
            I => \N__48914\
        );

    \I__10785\ : InMux
    port map (
            O => \N__48987\,
            I => \N__48914\
        );

    \I__10784\ : InMux
    port map (
            O => \N__48986\,
            I => \N__48914\
        );

    \I__10783\ : Span4Mux_v
    port map (
            O => \N__48977\,
            I => \N__48909\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__48972\,
            I => \N__48909\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__48967\,
            I => \N__48904\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__48956\,
            I => \N__48904\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__48953\,
            I => \N__48895\
        );

    \I__10778\ : Span4Mux_v
    port map (
            O => \N__48950\,
            I => \N__48895\
        );

    \I__10777\ : Span4Mux_v
    port map (
            O => \N__48945\,
            I => \N__48895\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__48936\,
            I => \N__48895\
        );

    \I__10775\ : InMux
    port map (
            O => \N__48935\,
            I => \N__48888\
        );

    \I__10774\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48888\
        );

    \I__10773\ : InMux
    port map (
            O => \N__48931\,
            I => \N__48888\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__48928\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__48923\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__48914\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__48909\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__48904\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10767\ : Odrv4
    port map (
            O => \N__48895\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__48888\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10765\ : InMux
    port map (
            O => \N__48873\,
            I => \N__48858\
        );

    \I__10764\ : CascadeMux
    port map (
            O => \N__48872\,
            I => \N__48855\
        );

    \I__10763\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48848\
        );

    \I__10762\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48841\
        );

    \I__10761\ : InMux
    port map (
            O => \N__48869\,
            I => \N__48841\
        );

    \I__10760\ : InMux
    port map (
            O => \N__48868\,
            I => \N__48841\
        );

    \I__10759\ : CascadeMux
    port map (
            O => \N__48867\,
            I => \N__48838\
        );

    \I__10758\ : CascadeMux
    port map (
            O => \N__48866\,
            I => \N__48835\
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__48865\,
            I => \N__48829\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__48864\,
            I => \N__48826\
        );

    \I__10755\ : CascadeMux
    port map (
            O => \N__48863\,
            I => \N__48816\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__48862\,
            I => \N__48812\
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__48861\,
            I => \N__48809\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__48858\,
            I => \N__48805\
        );

    \I__10751\ : InMux
    port map (
            O => \N__48855\,
            I => \N__48802\
        );

    \I__10750\ : InMux
    port map (
            O => \N__48854\,
            I => \N__48799\
        );

    \I__10749\ : InMux
    port map (
            O => \N__48853\,
            I => \N__48786\
        );

    \I__10748\ : InMux
    port map (
            O => \N__48852\,
            I => \N__48781\
        );

    \I__10747\ : InMux
    port map (
            O => \N__48851\,
            I => \N__48781\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__48848\,
            I => \N__48776\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__48841\,
            I => \N__48776\
        );

    \I__10744\ : InMux
    port map (
            O => \N__48838\,
            I => \N__48769\
        );

    \I__10743\ : InMux
    port map (
            O => \N__48835\,
            I => \N__48769\
        );

    \I__10742\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48769\
        );

    \I__10741\ : InMux
    port map (
            O => \N__48833\,
            I => \N__48764\
        );

    \I__10740\ : InMux
    port map (
            O => \N__48832\,
            I => \N__48764\
        );

    \I__10739\ : InMux
    port map (
            O => \N__48829\,
            I => \N__48759\
        );

    \I__10738\ : InMux
    port map (
            O => \N__48826\,
            I => \N__48759\
        );

    \I__10737\ : InMux
    port map (
            O => \N__48825\,
            I => \N__48744\
        );

    \I__10736\ : InMux
    port map (
            O => \N__48824\,
            I => \N__48744\
        );

    \I__10735\ : InMux
    port map (
            O => \N__48823\,
            I => \N__48744\
        );

    \I__10734\ : InMux
    port map (
            O => \N__48822\,
            I => \N__48744\
        );

    \I__10733\ : InMux
    port map (
            O => \N__48821\,
            I => \N__48744\
        );

    \I__10732\ : InMux
    port map (
            O => \N__48820\,
            I => \N__48744\
        );

    \I__10731\ : InMux
    port map (
            O => \N__48819\,
            I => \N__48744\
        );

    \I__10730\ : InMux
    port map (
            O => \N__48816\,
            I => \N__48730\
        );

    \I__10729\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48730\
        );

    \I__10728\ : InMux
    port map (
            O => \N__48812\,
            I => \N__48723\
        );

    \I__10727\ : InMux
    port map (
            O => \N__48809\,
            I => \N__48723\
        );

    \I__10726\ : InMux
    port map (
            O => \N__48808\,
            I => \N__48723\
        );

    \I__10725\ : Span4Mux_v
    port map (
            O => \N__48805\,
            I => \N__48718\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__48802\,
            I => \N__48718\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__48799\,
            I => \N__48715\
        );

    \I__10722\ : InMux
    port map (
            O => \N__48798\,
            I => \N__48710\
        );

    \I__10721\ : InMux
    port map (
            O => \N__48797\,
            I => \N__48710\
        );

    \I__10720\ : CascadeMux
    port map (
            O => \N__48796\,
            I => \N__48706\
        );

    \I__10719\ : CascadeMux
    port map (
            O => \N__48795\,
            I => \N__48703\
        );

    \I__10718\ : InMux
    port map (
            O => \N__48794\,
            I => \N__48687\
        );

    \I__10717\ : InMux
    port map (
            O => \N__48793\,
            I => \N__48687\
        );

    \I__10716\ : InMux
    port map (
            O => \N__48792\,
            I => \N__48687\
        );

    \I__10715\ : InMux
    port map (
            O => \N__48791\,
            I => \N__48687\
        );

    \I__10714\ : InMux
    port map (
            O => \N__48790\,
            I => \N__48682\
        );

    \I__10713\ : InMux
    port map (
            O => \N__48789\,
            I => \N__48682\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__48786\,
            I => \N__48671\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__48781\,
            I => \N__48671\
        );

    \I__10710\ : Span4Mux_v
    port map (
            O => \N__48776\,
            I => \N__48671\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__48769\,
            I => \N__48671\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__48764\,
            I => \N__48671\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__48759\,
            I => \N__48666\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__48744\,
            I => \N__48666\
        );

    \I__10705\ : InMux
    port map (
            O => \N__48743\,
            I => \N__48663\
        );

    \I__10704\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48654\
        );

    \I__10703\ : InMux
    port map (
            O => \N__48741\,
            I => \N__48654\
        );

    \I__10702\ : InMux
    port map (
            O => \N__48740\,
            I => \N__48654\
        );

    \I__10701\ : InMux
    port map (
            O => \N__48739\,
            I => \N__48654\
        );

    \I__10700\ : InMux
    port map (
            O => \N__48738\,
            I => \N__48647\
        );

    \I__10699\ : InMux
    port map (
            O => \N__48737\,
            I => \N__48647\
        );

    \I__10698\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48647\
        );

    \I__10697\ : CascadeMux
    port map (
            O => \N__48735\,
            I => \N__48632\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__48730\,
            I => \N__48627\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__48723\,
            I => \N__48627\
        );

    \I__10694\ : Span4Mux_v
    port map (
            O => \N__48718\,
            I => \N__48622\
        );

    \I__10693\ : Span4Mux_v
    port map (
            O => \N__48715\,
            I => \N__48622\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__48710\,
            I => \N__48619\
        );

    \I__10691\ : InMux
    port map (
            O => \N__48709\,
            I => \N__48610\
        );

    \I__10690\ : InMux
    port map (
            O => \N__48706\,
            I => \N__48610\
        );

    \I__10689\ : InMux
    port map (
            O => \N__48703\,
            I => \N__48610\
        );

    \I__10688\ : InMux
    port map (
            O => \N__48702\,
            I => \N__48610\
        );

    \I__10687\ : InMux
    port map (
            O => \N__48701\,
            I => \N__48599\
        );

    \I__10686\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48599\
        );

    \I__10685\ : InMux
    port map (
            O => \N__48699\,
            I => \N__48599\
        );

    \I__10684\ : InMux
    port map (
            O => \N__48698\,
            I => \N__48599\
        );

    \I__10683\ : InMux
    port map (
            O => \N__48697\,
            I => \N__48599\
        );

    \I__10682\ : InMux
    port map (
            O => \N__48696\,
            I => \N__48596\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__48687\,
            I => \N__48587\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__48682\,
            I => \N__48587\
        );

    \I__10679\ : Span4Mux_v
    port map (
            O => \N__48671\,
            I => \N__48587\
        );

    \I__10678\ : Span4Mux_h
    port map (
            O => \N__48666\,
            I => \N__48587\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__48663\,
            I => \N__48580\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__48654\,
            I => \N__48580\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__48647\,
            I => \N__48580\
        );

    \I__10674\ : InMux
    port map (
            O => \N__48646\,
            I => \N__48571\
        );

    \I__10673\ : InMux
    port map (
            O => \N__48645\,
            I => \N__48571\
        );

    \I__10672\ : InMux
    port map (
            O => \N__48644\,
            I => \N__48571\
        );

    \I__10671\ : InMux
    port map (
            O => \N__48643\,
            I => \N__48571\
        );

    \I__10670\ : InMux
    port map (
            O => \N__48642\,
            I => \N__48568\
        );

    \I__10669\ : InMux
    port map (
            O => \N__48641\,
            I => \N__48557\
        );

    \I__10668\ : InMux
    port map (
            O => \N__48640\,
            I => \N__48557\
        );

    \I__10667\ : InMux
    port map (
            O => \N__48639\,
            I => \N__48557\
        );

    \I__10666\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48557\
        );

    \I__10665\ : InMux
    port map (
            O => \N__48637\,
            I => \N__48557\
        );

    \I__10664\ : InMux
    port map (
            O => \N__48636\,
            I => \N__48554\
        );

    \I__10663\ : InMux
    port map (
            O => \N__48635\,
            I => \N__48549\
        );

    \I__10662\ : InMux
    port map (
            O => \N__48632\,
            I => \N__48549\
        );

    \I__10661\ : Odrv4
    port map (
            O => \N__48627\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10660\ : Odrv4
    port map (
            O => \N__48622\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__48619\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__48610\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__48599\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__48596\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10655\ : Odrv4
    port map (
            O => \N__48587\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__48580\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__48571\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__48568\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__48557\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__48554\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__48549\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10648\ : InMux
    port map (
            O => \N__48522\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_17\
        );

    \I__10647\ : InMux
    port map (
            O => \N__48519\,
            I => \N__48516\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__48516\,
            I => \N__48513\
        );

    \I__10645\ : Span4Mux_v
    port map (
            O => \N__48513\,
            I => \N__48510\
        );

    \I__10644\ : Odrv4
    port map (
            O => \N__48510\,
            I => \ppm_encoder_1.un1_init_pulses_11_18\
        );

    \I__10643\ : InMux
    port map (
            O => \N__48507\,
            I => \N__48504\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__48504\,
            I => \dron_frame_decoder_1.drone_H_disp_side_5\
        );

    \I__10641\ : InMux
    port map (
            O => \N__48501\,
            I => \N__48498\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__48498\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_5\
        );

    \I__10639\ : InMux
    port map (
            O => \N__48495\,
            I => \N__48492\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__48492\,
            I => \ppm_encoder_1.un1_init_pulses_11_5\
        );

    \I__10637\ : InMux
    port map (
            O => \N__48489\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_4\
        );

    \I__10636\ : InMux
    port map (
            O => \N__48486\,
            I => \N__48483\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__48483\,
            I => \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6\
        );

    \I__10634\ : CascadeMux
    port map (
            O => \N__48480\,
            I => \N__48477\
        );

    \I__10633\ : InMux
    port map (
            O => \N__48477\,
            I => \N__48474\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__48474\,
            I => \N__48471\
        );

    \I__10631\ : Span4Mux_h
    port map (
            O => \N__48471\,
            I => \N__48468\
        );

    \I__10630\ : Odrv4
    port map (
            O => \N__48468\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0\
        );

    \I__10629\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48462\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__48462\,
            I => \N__48459\
        );

    \I__10627\ : Span4Mux_h
    port map (
            O => \N__48459\,
            I => \N__48456\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__48456\,
            I => \ppm_encoder_1.un1_init_pulses_11_6\
        );

    \I__10625\ : InMux
    port map (
            O => \N__48453\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_5\
        );

    \I__10624\ : CascadeMux
    port map (
            O => \N__48450\,
            I => \N__48447\
        );

    \I__10623\ : InMux
    port map (
            O => \N__48447\,
            I => \N__48444\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__48444\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_7\
        );

    \I__10621\ : InMux
    port map (
            O => \N__48441\,
            I => \N__48438\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__48438\,
            I => \ppm_encoder_1.un1_init_pulses_11_7\
        );

    \I__10619\ : InMux
    port map (
            O => \N__48435\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_6\
        );

    \I__10618\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48429\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__48429\,
            I => \N__48426\
        );

    \I__10616\ : Odrv4
    port map (
            O => \N__48426\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_8\
        );

    \I__10615\ : InMux
    port map (
            O => \N__48423\,
            I => \N__48420\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__48420\,
            I => \ppm_encoder_1.un1_init_pulses_11_8\
        );

    \I__10613\ : InMux
    port map (
            O => \N__48417\,
            I => \bfn_18_16_0_\
        );

    \I__10612\ : InMux
    port map (
            O => \N__48414\,
            I => \N__48411\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__48411\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_9\
        );

    \I__10610\ : InMux
    port map (
            O => \N__48408\,
            I => \N__48405\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__48405\,
            I => \ppm_encoder_1.un1_init_pulses_11_9\
        );

    \I__10608\ : InMux
    port map (
            O => \N__48402\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_8\
        );

    \I__10607\ : InMux
    port map (
            O => \N__48399\,
            I => \N__48396\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__48396\,
            I => \N__48393\
        );

    \I__10605\ : Odrv4
    port map (
            O => \N__48393\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_10\
        );

    \I__10604\ : CascadeMux
    port map (
            O => \N__48390\,
            I => \N__48387\
        );

    \I__10603\ : InMux
    port map (
            O => \N__48387\,
            I => \N__48384\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__48384\,
            I => \N__48381\
        );

    \I__10601\ : Odrv4
    port map (
            O => \N__48381\,
            I => \ppm_encoder_1.un1_init_pulses_11_10\
        );

    \I__10600\ : InMux
    port map (
            O => \N__48378\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_9\
        );

    \I__10599\ : InMux
    port map (
            O => \N__48375\,
            I => \N__48372\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__48372\,
            I => \N__48369\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__48369\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_11\
        );

    \I__10596\ : CascadeMux
    port map (
            O => \N__48366\,
            I => \N__48363\
        );

    \I__10595\ : InMux
    port map (
            O => \N__48363\,
            I => \N__48360\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__48360\,
            I => \N__48357\
        );

    \I__10593\ : Odrv4
    port map (
            O => \N__48357\,
            I => \ppm_encoder_1.un1_init_pulses_11_11\
        );

    \I__10592\ : InMux
    port map (
            O => \N__48354\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_10\
        );

    \I__10591\ : InMux
    port map (
            O => \N__48351\,
            I => \N__48348\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__48348\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_12\
        );

    \I__10589\ : CascadeMux
    port map (
            O => \N__48345\,
            I => \N__48342\
        );

    \I__10588\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48339\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__48339\,
            I => \N__48336\
        );

    \I__10586\ : Odrv4
    port map (
            O => \N__48336\,
            I => \ppm_encoder_1.un1_init_pulses_11_12\
        );

    \I__10585\ : InMux
    port map (
            O => \N__48333\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_11\
        );

    \I__10584\ : InMux
    port map (
            O => \N__48330\,
            I => \N__48327\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__48327\,
            I => \N__48323\
        );

    \I__10582\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48320\
        );

    \I__10581\ : Span4Mux_h
    port map (
            O => \N__48323\,
            I => \N__48317\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__48320\,
            I => \N__48314\
        );

    \I__10579\ : Span4Mux_v
    port map (
            O => \N__48317\,
            I => \N__48310\
        );

    \I__10578\ : Span4Mux_h
    port map (
            O => \N__48314\,
            I => \N__48307\
        );

    \I__10577\ : InMux
    port map (
            O => \N__48313\,
            I => \N__48304\
        );

    \I__10576\ : Odrv4
    port map (
            O => \N__48310\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__10575\ : Odrv4
    port map (
            O => \N__48307\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__48304\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__10573\ : CascadeMux
    port map (
            O => \N__48297\,
            I => \N__48293\
        );

    \I__10572\ : CascadeMux
    port map (
            O => \N__48296\,
            I => \N__48287\
        );

    \I__10571\ : InMux
    port map (
            O => \N__48293\,
            I => \N__48282\
        );

    \I__10570\ : InMux
    port map (
            O => \N__48292\,
            I => \N__48279\
        );

    \I__10569\ : InMux
    port map (
            O => \N__48291\,
            I => \N__48276\
        );

    \I__10568\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48269\
        );

    \I__10567\ : InMux
    port map (
            O => \N__48287\,
            I => \N__48269\
        );

    \I__10566\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48264\
        );

    \I__10565\ : InMux
    port map (
            O => \N__48285\,
            I => \N__48264\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__48282\,
            I => \N__48259\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__48279\,
            I => \N__48259\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__48276\,
            I => \N__48256\
        );

    \I__10561\ : InMux
    port map (
            O => \N__48275\,
            I => \N__48251\
        );

    \I__10560\ : InMux
    port map (
            O => \N__48274\,
            I => \N__48251\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__48269\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__48264\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__10557\ : Odrv4
    port map (
            O => \N__48259\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__10556\ : Odrv12
    port map (
            O => \N__48256\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__48251\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__10554\ : InMux
    port map (
            O => \N__48240\,
            I => \N__48237\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__48237\,
            I => \N__48233\
        );

    \I__10552\ : InMux
    port map (
            O => \N__48236\,
            I => \N__48229\
        );

    \I__10551\ : Span4Mux_h
    port map (
            O => \N__48233\,
            I => \N__48226\
        );

    \I__10550\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48223\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__48229\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__10548\ : Odrv4
    port map (
            O => \N__48226\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__48223\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__10546\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48213\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__48213\,
            I => \N__48210\
        );

    \I__10544\ : Span4Mux_v
    port map (
            O => \N__48210\,
            I => \N__48207\
        );

    \I__10543\ : Odrv4
    port map (
            O => \N__48207\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2\
        );

    \I__10542\ : CascadeMux
    port map (
            O => \N__48204\,
            I => \N__48201\
        );

    \I__10541\ : InMux
    port map (
            O => \N__48201\,
            I => \N__48198\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__48198\,
            I => \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0\
        );

    \I__10539\ : InMux
    port map (
            O => \N__48195\,
            I => \N__48192\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__48192\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_1\
        );

    \I__10537\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48186\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__48186\,
            I => \N__48183\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__48183\,
            I => \N__48180\
        );

    \I__10534\ : Odrv4
    port map (
            O => \N__48180\,
            I => \ppm_encoder_1.un1_init_pulses_11_1\
        );

    \I__10533\ : InMux
    port map (
            O => \N__48177\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_0\
        );

    \I__10532\ : InMux
    port map (
            O => \N__48174\,
            I => \N__48171\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__48171\,
            I => \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2\
        );

    \I__10530\ : CascadeMux
    port map (
            O => \N__48168\,
            I => \N__48165\
        );

    \I__10529\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48162\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__48162\,
            I => \N__48159\
        );

    \I__10527\ : Span4Mux_v
    port map (
            O => \N__48159\,
            I => \N__48156\
        );

    \I__10526\ : Odrv4
    port map (
            O => \N__48156\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1\
        );

    \I__10525\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48150\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__48150\,
            I => \N__48147\
        );

    \I__10523\ : Span4Mux_v
    port map (
            O => \N__48147\,
            I => \N__48144\
        );

    \I__10522\ : Odrv4
    port map (
            O => \N__48144\,
            I => \ppm_encoder_1.un1_init_pulses_11_2\
        );

    \I__10521\ : InMux
    port map (
            O => \N__48141\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_1\
        );

    \I__10520\ : InMux
    port map (
            O => \N__48138\,
            I => \N__48135\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__48135\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_3\
        );

    \I__10518\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48129\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__48129\,
            I => \N__48126\
        );

    \I__10516\ : Span4Mux_h
    port map (
            O => \N__48126\,
            I => \N__48123\
        );

    \I__10515\ : Odrv4
    port map (
            O => \N__48123\,
            I => \ppm_encoder_1.un1_init_pulses_11_3\
        );

    \I__10514\ : InMux
    port map (
            O => \N__48120\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_2\
        );

    \I__10513\ : InMux
    port map (
            O => \N__48117\,
            I => \N__48114\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__48114\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_4\
        );

    \I__10511\ : InMux
    port map (
            O => \N__48111\,
            I => \N__48108\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__48108\,
            I => \N__48105\
        );

    \I__10509\ : Span4Mux_h
    port map (
            O => \N__48105\,
            I => \N__48102\
        );

    \I__10508\ : Odrv4
    port map (
            O => \N__48102\,
            I => \ppm_encoder_1.un1_init_pulses_11_4\
        );

    \I__10507\ : InMux
    port map (
            O => \N__48099\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_3\
        );

    \I__10506\ : InMux
    port map (
            O => \N__48096\,
            I => \N__48093\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__48093\,
            I => \pid_side.m9_e_4\
        );

    \I__10504\ : CascadeMux
    port map (
            O => \N__48090\,
            I => \pid_side.m9_e_5_cascade_\
        );

    \I__10503\ : InMux
    port map (
            O => \N__48087\,
            I => \N__48081\
        );

    \I__10502\ : InMux
    port map (
            O => \N__48086\,
            I => \N__48074\
        );

    \I__10501\ : InMux
    port map (
            O => \N__48085\,
            I => \N__48074\
        );

    \I__10500\ : InMux
    port map (
            O => \N__48084\,
            I => \N__48074\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__48081\,
            I => \pid_side.pid_prereg_esr_RNIFB07Z0Z_20\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__48074\,
            I => \pid_side.pid_prereg_esr_RNIFB07Z0Z_20\
        );

    \I__10497\ : CascadeMux
    port map (
            O => \N__48069\,
            I => \pid_side.pid_prereg_esr_RNIFB07Z0Z_20_cascade_\
        );

    \I__10496\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48063\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__48063\,
            I => \N__48059\
        );

    \I__10494\ : InMux
    port map (
            O => \N__48062\,
            I => \N__48056\
        );

    \I__10493\ : Span4Mux_h
    port map (
            O => \N__48059\,
            I => \N__48053\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__48056\,
            I => \N__48050\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__48053\,
            I => \N__48047\
        );

    \I__10490\ : Span12Mux_v
    port map (
            O => \N__48050\,
            I => \N__48044\
        );

    \I__10489\ : Span4Mux_v
    port map (
            O => \N__48047\,
            I => \N__48041\
        );

    \I__10488\ : Odrv12
    port map (
            O => \N__48044\,
            I => side_order_13
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__48041\,
            I => side_order_13
        );

    \I__10486\ : CEMux
    port map (
            O => \N__48036\,
            I => \N__48032\
        );

    \I__10485\ : CEMux
    port map (
            O => \N__48035\,
            I => \N__48029\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__48032\,
            I => \N__48026\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__48029\,
            I => \N__48022\
        );

    \I__10482\ : Span4Mux_h
    port map (
            O => \N__48026\,
            I => \N__48017\
        );

    \I__10481\ : CEMux
    port map (
            O => \N__48025\,
            I => \N__48014\
        );

    \I__10480\ : Span4Mux_h
    port map (
            O => \N__48022\,
            I => \N__48011\
        );

    \I__10479\ : CEMux
    port map (
            O => \N__48021\,
            I => \N__48008\
        );

    \I__10478\ : CEMux
    port map (
            O => \N__48020\,
            I => \N__48005\
        );

    \I__10477\ : Odrv4
    port map (
            O => \N__48017\,
            I => \pid_side.state_0_1\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__48014\,
            I => \pid_side.state_0_1\
        );

    \I__10475\ : Odrv4
    port map (
            O => \N__48011\,
            I => \pid_side.state_0_1\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__48008\,
            I => \pid_side.state_0_1\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__48005\,
            I => \pid_side.state_0_1\
        );

    \I__10472\ : SRMux
    port map (
            O => \N__47994\,
            I => \N__47991\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__47991\,
            I => \N__47988\
        );

    \I__10470\ : Span4Mux_v
    port map (
            O => \N__47988\,
            I => \N__47979\
        );

    \I__10469\ : SRMux
    port map (
            O => \N__47987\,
            I => \N__47976\
        );

    \I__10468\ : SRMux
    port map (
            O => \N__47986\,
            I => \N__47973\
        );

    \I__10467\ : SRMux
    port map (
            O => \N__47985\,
            I => \N__47970\
        );

    \I__10466\ : SRMux
    port map (
            O => \N__47984\,
            I => \N__47967\
        );

    \I__10465\ : SRMux
    port map (
            O => \N__47983\,
            I => \N__47964\
        );

    \I__10464\ : InMux
    port map (
            O => \N__47982\,
            I => \N__47961\
        );

    \I__10463\ : Odrv4
    port map (
            O => \N__47979\,
            I => \pid_side.un1_reset_0_i\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__47976\,
            I => \pid_side.un1_reset_0_i\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__47973\,
            I => \pid_side.un1_reset_0_i\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__47970\,
            I => \pid_side.un1_reset_0_i\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__47967\,
            I => \pid_side.un1_reset_0_i\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__47964\,
            I => \pid_side.un1_reset_0_i\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__47961\,
            I => \pid_side.un1_reset_0_i\
        );

    \I__10456\ : CascadeMux
    port map (
            O => \N__47946\,
            I => \N__47942\
        );

    \I__10455\ : InMux
    port map (
            O => \N__47945\,
            I => \N__47939\
        );

    \I__10454\ : InMux
    port map (
            O => \N__47942\,
            I => \N__47936\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__47939\,
            I => \N__47933\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__47936\,
            I => \N__47930\
        );

    \I__10451\ : Span4Mux_v
    port map (
            O => \N__47933\,
            I => \N__47927\
        );

    \I__10450\ : Span4Mux_v
    port map (
            O => \N__47930\,
            I => \N__47924\
        );

    \I__10449\ : Sp12to4
    port map (
            O => \N__47927\,
            I => \N__47921\
        );

    \I__10448\ : Sp12to4
    port map (
            O => \N__47924\,
            I => \N__47916\
        );

    \I__10447\ : Span12Mux_h
    port map (
            O => \N__47921\,
            I => \N__47916\
        );

    \I__10446\ : Odrv12
    port map (
            O => \N__47916\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__10445\ : InMux
    port map (
            O => \N__47913\,
            I => \N__47909\
        );

    \I__10444\ : InMux
    port map (
            O => \N__47912\,
            I => \N__47906\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__47909\,
            I => \N__47900\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__47906\,
            I => \N__47900\
        );

    \I__10441\ : InMux
    port map (
            O => \N__47905\,
            I => \N__47897\
        );

    \I__10440\ : Span4Mux_v
    port map (
            O => \N__47900\,
            I => \N__47894\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__47897\,
            I => \N__47891\
        );

    \I__10438\ : Span4Mux_v
    port map (
            O => \N__47894\,
            I => \N__47888\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__47891\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__10436\ : Odrv4
    port map (
            O => \N__47888\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__10435\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47880\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__47880\,
            I => \N__47877\
        );

    \I__10433\ : Span4Mux_h
    port map (
            O => \N__47877\,
            I => \N__47874\
        );

    \I__10432\ : Span4Mux_v
    port map (
            O => \N__47874\,
            I => \N__47866\
        );

    \I__10431\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47863\
        );

    \I__10430\ : InMux
    port map (
            O => \N__47872\,
            I => \N__47854\
        );

    \I__10429\ : InMux
    port map (
            O => \N__47871\,
            I => \N__47854\
        );

    \I__10428\ : InMux
    port map (
            O => \N__47870\,
            I => \N__47854\
        );

    \I__10427\ : InMux
    port map (
            O => \N__47869\,
            I => \N__47854\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__47866\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__47863\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__47854\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__10423\ : InMux
    port map (
            O => \N__47847\,
            I => \N__47844\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__47844\,
            I => \N__47841\
        );

    \I__10421\ : Span4Mux_h
    port map (
            O => \N__47841\,
            I => \N__47838\
        );

    \I__10420\ : Span4Mux_v
    port map (
            O => \N__47838\,
            I => \N__47833\
        );

    \I__10419\ : InMux
    port map (
            O => \N__47837\,
            I => \N__47828\
        );

    \I__10418\ : InMux
    port map (
            O => \N__47836\,
            I => \N__47828\
        );

    \I__10417\ : Odrv4
    port map (
            O => \N__47833\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__47828\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__10415\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47819\
        );

    \I__10414\ : CascadeMux
    port map (
            O => \N__47822\,
            I => \N__47816\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__47819\,
            I => \N__47812\
        );

    \I__10412\ : InMux
    port map (
            O => \N__47816\,
            I => \N__47809\
        );

    \I__10411\ : InMux
    port map (
            O => \N__47815\,
            I => \N__47806\
        );

    \I__10410\ : Span4Mux_h
    port map (
            O => \N__47812\,
            I => \N__47803\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__47809\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__47806\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__10407\ : Odrv4
    port map (
            O => \N__47803\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__10406\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47793\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__47793\,
            I => \N__47790\
        );

    \I__10404\ : Span4Mux_h
    port map (
            O => \N__47790\,
            I => \N__47787\
        );

    \I__10403\ : Span4Mux_h
    port map (
            O => \N__47787\,
            I => \N__47784\
        );

    \I__10402\ : Odrv4
    port map (
            O => \N__47784\,
            I => \pid_alt.state_RNIFCSD1Z0Z_0\
        );

    \I__10401\ : IoInMux
    port map (
            O => \N__47781\,
            I => \N__47778\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__47778\,
            I => \N__47775\
        );

    \I__10399\ : Span4Mux_s1_v
    port map (
            O => \N__47775\,
            I => \N__47772\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__47772\,
            I => \pid_alt.N_664_0\
        );

    \I__10397\ : InMux
    port map (
            O => \N__47769\,
            I => \N__47766\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__47766\,
            I => \N__47763\
        );

    \I__10395\ : Span4Mux_h
    port map (
            O => \N__47763\,
            I => \N__47758\
        );

    \I__10394\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47755\
        );

    \I__10393\ : InMux
    port map (
            O => \N__47761\,
            I => \N__47752\
        );

    \I__10392\ : Odrv4
    port map (
            O => \N__47758\,
            I => \pid_side.pid_preregZ0Z_0\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__47755\,
            I => \pid_side.pid_preregZ0Z_0\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__47752\,
            I => \pid_side.pid_preregZ0Z_0\
        );

    \I__10389\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47742\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__47742\,
            I => \N__47738\
        );

    \I__10387\ : CascadeMux
    port map (
            O => \N__47741\,
            I => \N__47735\
        );

    \I__10386\ : Span4Mux_h
    port map (
            O => \N__47738\,
            I => \N__47732\
        );

    \I__10385\ : InMux
    port map (
            O => \N__47735\,
            I => \N__47728\
        );

    \I__10384\ : Span4Mux_v
    port map (
            O => \N__47732\,
            I => \N__47725\
        );

    \I__10383\ : InMux
    port map (
            O => \N__47731\,
            I => \N__47722\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__47728\,
            I => \pid_side.pid_preregZ0Z_1\
        );

    \I__10381\ : Odrv4
    port map (
            O => \N__47725\,
            I => \pid_side.pid_preregZ0Z_1\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__47722\,
            I => \pid_side.pid_preregZ0Z_1\
        );

    \I__10379\ : IoInMux
    port map (
            O => \N__47715\,
            I => \N__47712\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__47712\,
            I => \N__47706\
        );

    \I__10377\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47700\
        );

    \I__10376\ : InMux
    port map (
            O => \N__47710\,
            I => \N__47700\
        );

    \I__10375\ : InMux
    port map (
            O => \N__47709\,
            I => \N__47697\
        );

    \I__10374\ : IoSpan4Mux
    port map (
            O => \N__47706\,
            I => \N__47694\
        );

    \I__10373\ : InMux
    port map (
            O => \N__47705\,
            I => \N__47691\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__47700\,
            I => \N__47688\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__47697\,
            I => \N__47685\
        );

    \I__10370\ : Span4Mux_s2_v
    port map (
            O => \N__47694\,
            I => \N__47681\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__47691\,
            I => \N__47678\
        );

    \I__10368\ : Span4Mux_v
    port map (
            O => \N__47688\,
            I => \N__47674\
        );

    \I__10367\ : Span4Mux_h
    port map (
            O => \N__47685\,
            I => \N__47671\
        );

    \I__10366\ : InMux
    port map (
            O => \N__47684\,
            I => \N__47668\
        );

    \I__10365\ : Span4Mux_v
    port map (
            O => \N__47681\,
            I => \N__47665\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__47678\,
            I => \N__47662\
        );

    \I__10363\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47658\
        );

    \I__10362\ : Sp12to4
    port map (
            O => \N__47674\,
            I => \N__47655\
        );

    \I__10361\ : Sp12to4
    port map (
            O => \N__47671\,
            I => \N__47652\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__47668\,
            I => \N__47649\
        );

    \I__10359\ : Span4Mux_v
    port map (
            O => \N__47665\,
            I => \N__47644\
        );

    \I__10358\ : Span4Mux_h
    port map (
            O => \N__47662\,
            I => \N__47644\
        );

    \I__10357\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47641\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__47658\,
            I => \N__47636\
        );

    \I__10355\ : Span12Mux_h
    port map (
            O => \N__47655\,
            I => \N__47636\
        );

    \I__10354\ : Span12Mux_v
    port map (
            O => \N__47652\,
            I => \N__47631\
        );

    \I__10353\ : Span12Mux_v
    port map (
            O => \N__47649\,
            I => \N__47631\
        );

    \I__10352\ : Odrv4
    port map (
            O => \N__47644\,
            I => \debug_CH1_0A_c\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__47641\,
            I => \debug_CH1_0A_c\
        );

    \I__10350\ : Odrv12
    port map (
            O => \N__47636\,
            I => \debug_CH1_0A_c\
        );

    \I__10349\ : Odrv12
    port map (
            O => \N__47631\,
            I => \debug_CH1_0A_c\
        );

    \I__10348\ : CascadeMux
    port map (
            O => \N__47622\,
            I => \N__47614\
        );

    \I__10347\ : InMux
    port map (
            O => \N__47621\,
            I => \N__47611\
        );

    \I__10346\ : InMux
    port map (
            O => \N__47620\,
            I => \N__47600\
        );

    \I__10345\ : InMux
    port map (
            O => \N__47619\,
            I => \N__47600\
        );

    \I__10344\ : InMux
    port map (
            O => \N__47618\,
            I => \N__47600\
        );

    \I__10343\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47600\
        );

    \I__10342\ : InMux
    port map (
            O => \N__47614\,
            I => \N__47600\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__47611\,
            I => \N__47597\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__47600\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__10339\ : Odrv12
    port map (
            O => \N__47597\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__10338\ : InMux
    port map (
            O => \N__47592\,
            I => \N__47589\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__47589\,
            I => \N__47586\
        );

    \I__10336\ : Odrv4
    port map (
            O => \N__47586\,
            I => \pid_side.m18_s_5\
        );

    \I__10335\ : InMux
    port map (
            O => \N__47583\,
            I => \N__47564\
        );

    \I__10334\ : InMux
    port map (
            O => \N__47582\,
            I => \N__47564\
        );

    \I__10333\ : InMux
    port map (
            O => \N__47581\,
            I => \N__47564\
        );

    \I__10332\ : InMux
    port map (
            O => \N__47580\,
            I => \N__47564\
        );

    \I__10331\ : InMux
    port map (
            O => \N__47579\,
            I => \N__47564\
        );

    \I__10330\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47564\
        );

    \I__10329\ : InMux
    port map (
            O => \N__47577\,
            I => \N__47561\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__47564\,
            I => \N__47558\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__47561\,
            I => \N__47555\
        );

    \I__10326\ : Span4Mux_h
    port map (
            O => \N__47558\,
            I => \N__47548\
        );

    \I__10325\ : Span4Mux_h
    port map (
            O => \N__47555\,
            I => \N__47545\
        );

    \I__10324\ : InMux
    port map (
            O => \N__47554\,
            I => \N__47540\
        );

    \I__10323\ : InMux
    port map (
            O => \N__47553\,
            I => \N__47540\
        );

    \I__10322\ : InMux
    port map (
            O => \N__47552\,
            I => \N__47537\
        );

    \I__10321\ : InMux
    port map (
            O => \N__47551\,
            I => \N__47534\
        );

    \I__10320\ : Odrv4
    port map (
            O => \N__47548\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__10319\ : Odrv4
    port map (
            O => \N__47545\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__47540\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__47537\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__47534\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__10315\ : InMux
    port map (
            O => \N__47523\,
            I => \N__47520\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__47520\,
            I => \pid_side.un1_reset_0_i_rn_0\
        );

    \I__10313\ : InMux
    port map (
            O => \N__47517\,
            I => \N__47514\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__47514\,
            I => \pid_side.m26_e_1\
        );

    \I__10311\ : InMux
    port map (
            O => \N__47511\,
            I => \N__47508\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__47508\,
            I => \N__47505\
        );

    \I__10309\ : Span4Mux_v
    port map (
            O => \N__47505\,
            I => \N__47502\
        );

    \I__10308\ : Odrv4
    port map (
            O => \N__47502\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\
        );

    \I__10307\ : InMux
    port map (
            O => \N__47499\,
            I => \N__47496\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__47496\,
            I => \N__47493\
        );

    \I__10305\ : Odrv4
    port map (
            O => \N__47493\,
            I => \ppm_encoder_1.un1_init_pulses_10_11\
        );

    \I__10304\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47487\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__47487\,
            I => \N__47484\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__47484\,
            I => \N__47480\
        );

    \I__10301\ : InMux
    port map (
            O => \N__47483\,
            I => \N__47477\
        );

    \I__10300\ : Span4Mux_v
    port map (
            O => \N__47480\,
            I => \N__47472\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__47477\,
            I => \N__47472\
        );

    \I__10298\ : Odrv4
    port map (
            O => \N__47472\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__10297\ : InMux
    port map (
            O => \N__47469\,
            I => \N__47458\
        );

    \I__10296\ : InMux
    port map (
            O => \N__47468\,
            I => \N__47453\
        );

    \I__10295\ : InMux
    port map (
            O => \N__47467\,
            I => \N__47448\
        );

    \I__10294\ : InMux
    port map (
            O => \N__47466\,
            I => \N__47448\
        );

    \I__10293\ : InMux
    port map (
            O => \N__47465\,
            I => \N__47441\
        );

    \I__10292\ : InMux
    port map (
            O => \N__47464\,
            I => \N__47441\
        );

    \I__10291\ : InMux
    port map (
            O => \N__47463\,
            I => \N__47441\
        );

    \I__10290\ : InMux
    port map (
            O => \N__47462\,
            I => \N__47436\
        );

    \I__10289\ : InMux
    port map (
            O => \N__47461\,
            I => \N__47436\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__47458\,
            I => \N__47433\
        );

    \I__10287\ : InMux
    port map (
            O => \N__47457\,
            I => \N__47428\
        );

    \I__10286\ : InMux
    port map (
            O => \N__47456\,
            I => \N__47428\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__47453\,
            I => \N__47425\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__47448\,
            I => \N__47410\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__47441\,
            I => \N__47410\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__47436\,
            I => \N__47410\
        );

    \I__10281\ : Span4Mux_h
    port map (
            O => \N__47433\,
            I => \N__47407\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__47428\,
            I => \N__47404\
        );

    \I__10279\ : Span4Mux_h
    port map (
            O => \N__47425\,
            I => \N__47401\
        );

    \I__10278\ : InMux
    port map (
            O => \N__47424\,
            I => \N__47394\
        );

    \I__10277\ : InMux
    port map (
            O => \N__47423\,
            I => \N__47394\
        );

    \I__10276\ : InMux
    port map (
            O => \N__47422\,
            I => \N__47394\
        );

    \I__10275\ : InMux
    port map (
            O => \N__47421\,
            I => \N__47387\
        );

    \I__10274\ : InMux
    port map (
            O => \N__47420\,
            I => \N__47387\
        );

    \I__10273\ : InMux
    port map (
            O => \N__47419\,
            I => \N__47387\
        );

    \I__10272\ : InMux
    port map (
            O => \N__47418\,
            I => \N__47384\
        );

    \I__10271\ : InMux
    port map (
            O => \N__47417\,
            I => \N__47381\
        );

    \I__10270\ : Span4Mux_v
    port map (
            O => \N__47410\,
            I => \N__47378\
        );

    \I__10269\ : Span4Mux_v
    port map (
            O => \N__47407\,
            I => \N__47375\
        );

    \I__10268\ : Span4Mux_h
    port map (
            O => \N__47404\,
            I => \N__47372\
        );

    \I__10267\ : Span4Mux_v
    port map (
            O => \N__47401\,
            I => \N__47369\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__47394\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__47387\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__47384\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__47381\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10262\ : Odrv4
    port map (
            O => \N__47378\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10261\ : Odrv4
    port map (
            O => \N__47375\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10260\ : Odrv4
    port map (
            O => \N__47372\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10259\ : Odrv4
    port map (
            O => \N__47369\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__10258\ : CascadeMux
    port map (
            O => \N__47352\,
            I => \N__47340\
        );

    \I__10257\ : CascadeMux
    port map (
            O => \N__47351\,
            I => \N__47337\
        );

    \I__10256\ : CascadeMux
    port map (
            O => \N__47350\,
            I => \N__47334\
        );

    \I__10255\ : CascadeMux
    port map (
            O => \N__47349\,
            I => \N__47331\
        );

    \I__10254\ : CascadeMux
    port map (
            O => \N__47348\,
            I => \N__47328\
        );

    \I__10253\ : CascadeMux
    port map (
            O => \N__47347\,
            I => \N__47324\
        );

    \I__10252\ : CascadeMux
    port map (
            O => \N__47346\,
            I => \N__47321\
        );

    \I__10251\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47308\
        );

    \I__10250\ : InMux
    port map (
            O => \N__47344\,
            I => \N__47308\
        );

    \I__10249\ : InMux
    port map (
            O => \N__47343\,
            I => \N__47308\
        );

    \I__10248\ : InMux
    port map (
            O => \N__47340\,
            I => \N__47301\
        );

    \I__10247\ : InMux
    port map (
            O => \N__47337\,
            I => \N__47301\
        );

    \I__10246\ : InMux
    port map (
            O => \N__47334\,
            I => \N__47301\
        );

    \I__10245\ : InMux
    port map (
            O => \N__47331\,
            I => \N__47298\
        );

    \I__10244\ : InMux
    port map (
            O => \N__47328\,
            I => \N__47295\
        );

    \I__10243\ : InMux
    port map (
            O => \N__47327\,
            I => \N__47292\
        );

    \I__10242\ : InMux
    port map (
            O => \N__47324\,
            I => \N__47287\
        );

    \I__10241\ : InMux
    port map (
            O => \N__47321\,
            I => \N__47287\
        );

    \I__10240\ : CascadeMux
    port map (
            O => \N__47320\,
            I => \N__47284\
        );

    \I__10239\ : CascadeMux
    port map (
            O => \N__47319\,
            I => \N__47281\
        );

    \I__10238\ : CascadeMux
    port map (
            O => \N__47318\,
            I => \N__47278\
        );

    \I__10237\ : CascadeMux
    port map (
            O => \N__47317\,
            I => \N__47274\
        );

    \I__10236\ : CascadeMux
    port map (
            O => \N__47316\,
            I => \N__47271\
        );

    \I__10235\ : CascadeMux
    port map (
            O => \N__47315\,
            I => \N__47268\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__47308\,
            I => \N__47265\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__47301\,
            I => \N__47256\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__47298\,
            I => \N__47256\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__47295\,
            I => \N__47256\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__47292\,
            I => \N__47256\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__47287\,
            I => \N__47253\
        );

    \I__10228\ : InMux
    port map (
            O => \N__47284\,
            I => \N__47248\
        );

    \I__10227\ : InMux
    port map (
            O => \N__47281\,
            I => \N__47248\
        );

    \I__10226\ : InMux
    port map (
            O => \N__47278\,
            I => \N__47245\
        );

    \I__10225\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47242\
        );

    \I__10224\ : InMux
    port map (
            O => \N__47274\,
            I => \N__47236\
        );

    \I__10223\ : InMux
    port map (
            O => \N__47271\,
            I => \N__47236\
        );

    \I__10222\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47233\
        );

    \I__10221\ : Span4Mux_v
    port map (
            O => \N__47265\,
            I => \N__47230\
        );

    \I__10220\ : Span4Mux_v
    port map (
            O => \N__47256\,
            I => \N__47225\
        );

    \I__10219\ : Span4Mux_h
    port map (
            O => \N__47253\,
            I => \N__47225\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__47248\,
            I => \N__47218\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__47245\,
            I => \N__47218\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__47242\,
            I => \N__47218\
        );

    \I__10215\ : InMux
    port map (
            O => \N__47241\,
            I => \N__47215\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__47236\,
            I => \N__47210\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__47233\,
            I => \N__47210\
        );

    \I__10212\ : Odrv4
    port map (
            O => \N__47230\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__10211\ : Odrv4
    port map (
            O => \N__47225\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__10210\ : Odrv12
    port map (
            O => \N__47218\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__47215\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__10208\ : Odrv4
    port map (
            O => \N__47210\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__10207\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47196\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__47196\,
            I => \N__47193\
        );

    \I__10205\ : Odrv4
    port map (
            O => \N__47193\,
            I => \ppm_encoder_1.un1_init_pulses_10_12\
        );

    \I__10204\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47181\
        );

    \I__10203\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47181\
        );

    \I__10202\ : InMux
    port map (
            O => \N__47188\,
            I => \N__47181\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__47181\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__10200\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47174\
        );

    \I__10199\ : InMux
    port map (
            O => \N__47177\,
            I => \N__47166\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__47174\,
            I => \N__47158\
        );

    \I__10197\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47153\
        );

    \I__10196\ : InMux
    port map (
            O => \N__47172\,
            I => \N__47153\
        );

    \I__10195\ : InMux
    port map (
            O => \N__47171\,
            I => \N__47147\
        );

    \I__10194\ : InMux
    port map (
            O => \N__47170\,
            I => \N__47144\
        );

    \I__10193\ : InMux
    port map (
            O => \N__47169\,
            I => \N__47141\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__47166\,
            I => \N__47138\
        );

    \I__10191\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47135\
        );

    \I__10190\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47132\
        );

    \I__10189\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47129\
        );

    \I__10188\ : InMux
    port map (
            O => \N__47162\,
            I => \N__47123\
        );

    \I__10187\ : InMux
    port map (
            O => \N__47161\,
            I => \N__47120\
        );

    \I__10186\ : Span4Mux_h
    port map (
            O => \N__47158\,
            I => \N__47115\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__47153\,
            I => \N__47115\
        );

    \I__10184\ : InMux
    port map (
            O => \N__47152\,
            I => \N__47110\
        );

    \I__10183\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47110\
        );

    \I__10182\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47106\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__47147\,
            I => \N__47093\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__47144\,
            I => \N__47093\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__47141\,
            I => \N__47093\
        );

    \I__10178\ : Span4Mux_v
    port map (
            O => \N__47138\,
            I => \N__47093\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__47135\,
            I => \N__47093\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__47132\,
            I => \N__47093\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__47129\,
            I => \N__47090\
        );

    \I__10174\ : InMux
    port map (
            O => \N__47128\,
            I => \N__47087\
        );

    \I__10173\ : InMux
    port map (
            O => \N__47127\,
            I => \N__47084\
        );

    \I__10172\ : InMux
    port map (
            O => \N__47126\,
            I => \N__47081\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__47123\,
            I => \N__47072\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__47120\,
            I => \N__47072\
        );

    \I__10169\ : Span4Mux_v
    port map (
            O => \N__47115\,
            I => \N__47072\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__47110\,
            I => \N__47072\
        );

    \I__10167\ : InMux
    port map (
            O => \N__47109\,
            I => \N__47069\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__47106\,
            I => \N__47064\
        );

    \I__10165\ : Span4Mux_v
    port map (
            O => \N__47093\,
            I => \N__47064\
        );

    \I__10164\ : Span4Mux_h
    port map (
            O => \N__47090\,
            I => \N__47061\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__47087\,
            I => \N__47054\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__47084\,
            I => \N__47054\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__47081\,
            I => \N__47054\
        );

    \I__10160\ : Span4Mux_v
    port map (
            O => \N__47072\,
            I => \N__47051\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__47069\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10158\ : Odrv4
    port map (
            O => \N__47064\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10157\ : Odrv4
    port map (
            O => \N__47061\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10156\ : Odrv4
    port map (
            O => \N__47054\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10155\ : Odrv4
    port map (
            O => \N__47051\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10154\ : InMux
    port map (
            O => \N__47040\,
            I => \N__47036\
        );

    \I__10153\ : InMux
    port map (
            O => \N__47039\,
            I => \N__47033\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__47036\,
            I => \N__47029\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__47033\,
            I => \N__47026\
        );

    \I__10150\ : CascadeMux
    port map (
            O => \N__47032\,
            I => \N__47023\
        );

    \I__10149\ : Span4Mux_h
    port map (
            O => \N__47029\,
            I => \N__47020\
        );

    \I__10148\ : Span4Mux_h
    port map (
            O => \N__47026\,
            I => \N__47017\
        );

    \I__10147\ : InMux
    port map (
            O => \N__47023\,
            I => \N__47014\
        );

    \I__10146\ : Span4Mux_h
    port map (
            O => \N__47020\,
            I => \N__47009\
        );

    \I__10145\ : Span4Mux_h
    port map (
            O => \N__47017\,
            I => \N__47009\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__47014\,
            I => \ppm_encoder_1.elevatorZ0Z_2\
        );

    \I__10143\ : Odrv4
    port map (
            O => \N__47009\,
            I => \ppm_encoder_1.elevatorZ0Z_2\
        );

    \I__10142\ : InMux
    port map (
            O => \N__47004\,
            I => \N__47001\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__47001\,
            I => \N__46997\
        );

    \I__10140\ : InMux
    port map (
            O => \N__47000\,
            I => \N__46994\
        );

    \I__10139\ : Span4Mux_v
    port map (
            O => \N__46997\,
            I => \N__46988\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__46994\,
            I => \N__46988\
        );

    \I__10137\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46985\
        );

    \I__10136\ : Span4Mux_h
    port map (
            O => \N__46988\,
            I => \N__46982\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__46985\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__10134\ : Odrv4
    port map (
            O => \N__46982\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__10133\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46974\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__46974\,
            I => \N__46971\
        );

    \I__10131\ : Odrv12
    port map (
            O => \N__46971\,
            I => \ppm_encoder_1.N_288\
        );

    \I__10130\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46965\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__46965\,
            I => \N__46962\
        );

    \I__10128\ : Odrv4
    port map (
            O => \N__46962\,
            I => \ppm_encoder_1.N_290\
        );

    \I__10127\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46956\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__46956\,
            I => \N__46953\
        );

    \I__10125\ : Span4Mux_h
    port map (
            O => \N__46953\,
            I => \N__46948\
        );

    \I__10124\ : InMux
    port map (
            O => \N__46952\,
            I => \N__46945\
        );

    \I__10123\ : InMux
    port map (
            O => \N__46951\,
            I => \N__46942\
        );

    \I__10122\ : Span4Mux_v
    port map (
            O => \N__46948\,
            I => \N__46937\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__46945\,
            I => \N__46937\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__46942\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__10119\ : Odrv4
    port map (
            O => \N__46937\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__10118\ : InMux
    port map (
            O => \N__46932\,
            I => \N__46929\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__46929\,
            I => \N__46926\
        );

    \I__10116\ : Span4Mux_v
    port map (
            O => \N__46926\,
            I => \N__46923\
        );

    \I__10115\ : Odrv4
    port map (
            O => \N__46923\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\
        );

    \I__10114\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46914\
        );

    \I__10113\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46914\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__46914\,
            I => \N__46911\
        );

    \I__10111\ : Odrv12
    port map (
            O => \N__46911\,
            I => \pid_front.error_d_reg_prevZ0Z_1\
        );

    \I__10110\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46901\
        );

    \I__10109\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46901\
        );

    \I__10108\ : CascadeMux
    port map (
            O => \N__46906\,
            I => \N__46897\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__46901\,
            I => \N__46894\
        );

    \I__10106\ : InMux
    port map (
            O => \N__46900\,
            I => \N__46891\
        );

    \I__10105\ : InMux
    port map (
            O => \N__46897\,
            I => \N__46888\
        );

    \I__10104\ : Span4Mux_h
    port map (
            O => \N__46894\,
            I => \N__46885\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__46891\,
            I => \N__46880\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__46888\,
            I => \N__46880\
        );

    \I__10101\ : Span4Mux_v
    port map (
            O => \N__46885\,
            I => \N__46875\
        );

    \I__10100\ : Span4Mux_v
    port map (
            O => \N__46880\,
            I => \N__46875\
        );

    \I__10099\ : Span4Mux_v
    port map (
            O => \N__46875\,
            I => \N__46872\
        );

    \I__10098\ : Odrv4
    port map (
            O => \N__46872\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_153_d\
        );

    \I__10097\ : CascadeMux
    port map (
            O => \N__46869\,
            I => \N__46866\
        );

    \I__10096\ : InMux
    port map (
            O => \N__46866\,
            I => \N__46862\
        );

    \I__10095\ : InMux
    port map (
            O => \N__46865\,
            I => \N__46859\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__46862\,
            I => \N__46856\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__46859\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__10092\ : Odrv12
    port map (
            O => \N__46856\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__10091\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46847\
        );

    \I__10090\ : InMux
    port map (
            O => \N__46850\,
            I => \N__46844\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__46847\,
            I => \N__46841\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__46844\,
            I => \N__46838\
        );

    \I__10087\ : Span4Mux_v
    port map (
            O => \N__46841\,
            I => \N__46835\
        );

    \I__10086\ : Span12Mux_v
    port map (
            O => \N__46838\,
            I => \N__46832\
        );

    \I__10085\ : Span4Mux_h
    port map (
            O => \N__46835\,
            I => \N__46829\
        );

    \I__10084\ : Odrv12
    port map (
            O => \N__46832\,
            I => \pid_front.error_d_reg_prevZ0Z_11\
        );

    \I__10083\ : Odrv4
    port map (
            O => \N__46829\,
            I => \pid_front.error_d_reg_prevZ0Z_11\
        );

    \I__10082\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46821\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__46821\,
            I => \N__46818\
        );

    \I__10080\ : Span4Mux_h
    port map (
            O => \N__46818\,
            I => \N__46814\
        );

    \I__10079\ : CascadeMux
    port map (
            O => \N__46817\,
            I => \N__46811\
        );

    \I__10078\ : Span4Mux_v
    port map (
            O => \N__46814\,
            I => \N__46808\
        );

    \I__10077\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46805\
        );

    \I__10076\ : Odrv4
    port map (
            O => \N__46808\,
            I => scaler_4_data_4
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__46805\,
            I => scaler_4_data_4
        );

    \I__10074\ : InMux
    port map (
            O => \N__46800\,
            I => \N__46797\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__46797\,
            I => \N__46793\
        );

    \I__10072\ : InMux
    port map (
            O => \N__46796\,
            I => \N__46790\
        );

    \I__10071\ : Span4Mux_h
    port map (
            O => \N__46793\,
            I => \N__46787\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__46790\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__10069\ : Odrv4
    port map (
            O => \N__46787\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__10068\ : CEMux
    port map (
            O => \N__46782\,
            I => \N__46778\
        );

    \I__10067\ : CEMux
    port map (
            O => \N__46781\,
            I => \N__46773\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__46778\,
            I => \N__46770\
        );

    \I__10065\ : CEMux
    port map (
            O => \N__46777\,
            I => \N__46767\
        );

    \I__10064\ : CEMux
    port map (
            O => \N__46776\,
            I => \N__46764\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46759\
        );

    \I__10062\ : Span4Mux_h
    port map (
            O => \N__46770\,
            I => \N__46754\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__46767\,
            I => \N__46754\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__46764\,
            I => \N__46751\
        );

    \I__10059\ : CEMux
    port map (
            O => \N__46763\,
            I => \N__46748\
        );

    \I__10058\ : CEMux
    port map (
            O => \N__46762\,
            I => \N__46745\
        );

    \I__10057\ : Span4Mux_v
    port map (
            O => \N__46759\,
            I => \N__46742\
        );

    \I__10056\ : Span4Mux_v
    port map (
            O => \N__46754\,
            I => \N__46735\
        );

    \I__10055\ : Span4Mux_v
    port map (
            O => \N__46751\,
            I => \N__46735\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__46748\,
            I => \N__46735\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__46745\,
            I => \N__46732\
        );

    \I__10052\ : Span4Mux_h
    port map (
            O => \N__46742\,
            I => \N__46727\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__46735\,
            I => \N__46727\
        );

    \I__10050\ : Span4Mux_v
    port map (
            O => \N__46732\,
            I => \N__46724\
        );

    \I__10049\ : Span4Mux_h
    port map (
            O => \N__46727\,
            I => \N__46721\
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__46724\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__10047\ : Odrv4
    port map (
            O => \N__46721\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__10046\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46713\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__46713\,
            I => \N__46709\
        );

    \I__10044\ : InMux
    port map (
            O => \N__46712\,
            I => \N__46705\
        );

    \I__10043\ : Span12Mux_v
    port map (
            O => \N__46709\,
            I => \N__46702\
        );

    \I__10042\ : InMux
    port map (
            O => \N__46708\,
            I => \N__46699\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__46705\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__10040\ : Odrv12
    port map (
            O => \N__46702\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__46699\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__10038\ : CascadeMux
    port map (
            O => \N__46692\,
            I => \ppm_encoder_1.N_314_cascade_\
        );

    \I__10037\ : CascadeMux
    port map (
            O => \N__46689\,
            I => \N__46686\
        );

    \I__10036\ : InMux
    port map (
            O => \N__46686\,
            I => \N__46677\
        );

    \I__10035\ : InMux
    port map (
            O => \N__46685\,
            I => \N__46677\
        );

    \I__10034\ : InMux
    port map (
            O => \N__46684\,
            I => \N__46677\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__46677\,
            I => \N__46673\
        );

    \I__10032\ : InMux
    port map (
            O => \N__46676\,
            I => \N__46670\
        );

    \I__10031\ : Sp12to4
    port map (
            O => \N__46673\,
            I => \N__46665\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__46670\,
            I => \N__46665\
        );

    \I__10029\ : Span12Mux_s10_h
    port map (
            O => \N__46665\,
            I => \N__46661\
        );

    \I__10028\ : InMux
    port map (
            O => \N__46664\,
            I => \N__46658\
        );

    \I__10027\ : Odrv12
    port map (
            O => \N__46661\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__46658\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__10025\ : InMux
    port map (
            O => \N__46653\,
            I => \N__46650\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__46650\,
            I => \N__46647\
        );

    \I__10023\ : Span4Mux_h
    port map (
            O => \N__46647\,
            I => \N__46644\
        );

    \I__10022\ : Odrv4
    port map (
            O => \N__46644\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\
        );

    \I__10021\ : InMux
    port map (
            O => \N__46641\,
            I => \N__46638\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__46638\,
            I => \N__46634\
        );

    \I__10019\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46631\
        );

    \I__10018\ : Span4Mux_h
    port map (
            O => \N__46634\,
            I => \N__46628\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__46631\,
            I => \N__46625\
        );

    \I__10016\ : Span4Mux_v
    port map (
            O => \N__46628\,
            I => \N__46620\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__46625\,
            I => \N__46620\
        );

    \I__10014\ : Odrv4
    port map (
            O => \N__46620\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__10013\ : InMux
    port map (
            O => \N__46617\,
            I => \N__46614\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__46614\,
            I => \N__46611\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__46611\,
            I => \ppm_encoder_1.un1_init_pulses_10_10\
        );

    \I__10010\ : InMux
    port map (
            O => \N__46608\,
            I => \N__46605\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__46605\,
            I => \N__46601\
        );

    \I__10008\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46598\
        );

    \I__10007\ : Span4Mux_h
    port map (
            O => \N__46601\,
            I => \N__46595\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__46598\,
            I => \N__46592\
        );

    \I__10005\ : Odrv4
    port map (
            O => \N__46595\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__10004\ : Odrv4
    port map (
            O => \N__46592\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__10003\ : InMux
    port map (
            O => \N__46587\,
            I => \N__46578\
        );

    \I__10002\ : InMux
    port map (
            O => \N__46586\,
            I => \N__46578\
        );

    \I__10001\ : InMux
    port map (
            O => \N__46585\,
            I => \N__46578\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__46578\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__9999\ : InMux
    port map (
            O => \N__46575\,
            I => \N__46561\
        );

    \I__9998\ : InMux
    port map (
            O => \N__46574\,
            I => \N__46558\
        );

    \I__9997\ : InMux
    port map (
            O => \N__46573\,
            I => \N__46555\
        );

    \I__9996\ : CascadeMux
    port map (
            O => \N__46572\,
            I => \N__46550\
        );

    \I__9995\ : InMux
    port map (
            O => \N__46571\,
            I => \N__46547\
        );

    \I__9994\ : InMux
    port map (
            O => \N__46570\,
            I => \N__46544\
        );

    \I__9993\ : InMux
    port map (
            O => \N__46569\,
            I => \N__46541\
        );

    \I__9992\ : InMux
    port map (
            O => \N__46568\,
            I => \N__46536\
        );

    \I__9991\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46536\
        );

    \I__9990\ : InMux
    port map (
            O => \N__46566\,
            I => \N__46531\
        );

    \I__9989\ : InMux
    port map (
            O => \N__46565\,
            I => \N__46531\
        );

    \I__9988\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46528\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__46561\,
            I => \N__46525\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__46558\,
            I => \N__46520\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__46555\,
            I => \N__46520\
        );

    \I__9984\ : InMux
    port map (
            O => \N__46554\,
            I => \N__46513\
        );

    \I__9983\ : InMux
    port map (
            O => \N__46553\,
            I => \N__46513\
        );

    \I__9982\ : InMux
    port map (
            O => \N__46550\,
            I => \N__46513\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__46547\,
            I => \N__46510\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__46544\,
            I => \N__46505\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__46541\,
            I => \N__46505\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__46536\,
            I => \N__46502\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__46531\,
            I => \N__46498\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__46528\,
            I => \N__46495\
        );

    \I__9975\ : Span4Mux_v
    port map (
            O => \N__46525\,
            I => \N__46492\
        );

    \I__9974\ : Span4Mux_v
    port map (
            O => \N__46520\,
            I => \N__46485\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__46513\,
            I => \N__46485\
        );

    \I__9972\ : Span4Mux_h
    port map (
            O => \N__46510\,
            I => \N__46485\
        );

    \I__9971\ : Span4Mux_v
    port map (
            O => \N__46505\,
            I => \N__46480\
        );

    \I__9970\ : Span4Mux_h
    port map (
            O => \N__46502\,
            I => \N__46480\
        );

    \I__9969\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46477\
        );

    \I__9968\ : Span4Mux_v
    port map (
            O => \N__46498\,
            I => \N__46470\
        );

    \I__9967\ : Span4Mux_v
    port map (
            O => \N__46495\,
            I => \N__46470\
        );

    \I__9966\ : Span4Mux_h
    port map (
            O => \N__46492\,
            I => \N__46470\
        );

    \I__9965\ : Span4Mux_v
    port map (
            O => \N__46485\,
            I => \N__46467\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__46480\,
            I => \N__46464\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__46477\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__46470\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9961\ : Odrv4
    port map (
            O => \N__46467\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9960\ : Odrv4
    port map (
            O => \N__46464\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__46455\,
            I => \N__46450\
        );

    \I__9958\ : CascadeMux
    port map (
            O => \N__46454\,
            I => \N__46441\
        );

    \I__9957\ : CascadeMux
    port map (
            O => \N__46453\,
            I => \N__46438\
        );

    \I__9956\ : InMux
    port map (
            O => \N__46450\,
            I => \N__46433\
        );

    \I__9955\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46426\
        );

    \I__9954\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46426\
        );

    \I__9953\ : InMux
    port map (
            O => \N__46447\,
            I => \N__46426\
        );

    \I__9952\ : CascadeMux
    port map (
            O => \N__46446\,
            I => \N__46423\
        );

    \I__9951\ : CascadeMux
    port map (
            O => \N__46445\,
            I => \N__46420\
        );

    \I__9950\ : CascadeMux
    port map (
            O => \N__46444\,
            I => \N__46417\
        );

    \I__9949\ : InMux
    port map (
            O => \N__46441\,
            I => \N__46414\
        );

    \I__9948\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46411\
        );

    \I__9947\ : CascadeMux
    port map (
            O => \N__46437\,
            I => \N__46408\
        );

    \I__9946\ : InMux
    port map (
            O => \N__46436\,
            I => \N__46404\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__46433\,
            I => \N__46399\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__46426\,
            I => \N__46399\
        );

    \I__9943\ : InMux
    port map (
            O => \N__46423\,
            I => \N__46396\
        );

    \I__9942\ : InMux
    port map (
            O => \N__46420\,
            I => \N__46393\
        );

    \I__9941\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46390\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__46414\,
            I => \N__46383\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__46411\,
            I => \N__46383\
        );

    \I__9938\ : InMux
    port map (
            O => \N__46408\,
            I => \N__46378\
        );

    \I__9937\ : InMux
    port map (
            O => \N__46407\,
            I => \N__46378\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__46404\,
            I => \N__46371\
        );

    \I__9935\ : Span4Mux_v
    port map (
            O => \N__46399\,
            I => \N__46371\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__46396\,
            I => \N__46371\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__46393\,
            I => \N__46366\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46366\
        );

    \I__9931\ : InMux
    port map (
            O => \N__46389\,
            I => \N__46361\
        );

    \I__9930\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46361\
        );

    \I__9929\ : Span4Mux_v
    port map (
            O => \N__46383\,
            I => \N__46357\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__46378\,
            I => \N__46354\
        );

    \I__9927\ : Span4Mux_v
    port map (
            O => \N__46371\,
            I => \N__46349\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__46366\,
            I => \N__46344\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__46361\,
            I => \N__46344\
        );

    \I__9924\ : InMux
    port map (
            O => \N__46360\,
            I => \N__46341\
        );

    \I__9923\ : Span4Mux_h
    port map (
            O => \N__46357\,
            I => \N__46336\
        );

    \I__9922\ : Span4Mux_h
    port map (
            O => \N__46354\,
            I => \N__46336\
        );

    \I__9921\ : CascadeMux
    port map (
            O => \N__46353\,
            I => \N__46333\
        );

    \I__9920\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46329\
        );

    \I__9919\ : Span4Mux_h
    port map (
            O => \N__46349\,
            I => \N__46326\
        );

    \I__9918\ : Sp12to4
    port map (
            O => \N__46344\,
            I => \N__46323\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__46341\,
            I => \N__46318\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__46336\,
            I => \N__46318\
        );

    \I__9915\ : InMux
    port map (
            O => \N__46333\,
            I => \N__46313\
        );

    \I__9914\ : InMux
    port map (
            O => \N__46332\,
            I => \N__46313\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__46329\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9912\ : Odrv4
    port map (
            O => \N__46326\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9911\ : Odrv12
    port map (
            O => \N__46323\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9910\ : Odrv4
    port map (
            O => \N__46318\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__46313\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9908\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46298\
        );

    \I__9907\ : InMux
    port map (
            O => \N__46301\,
            I => \N__46295\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__46298\,
            I => \N__46292\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__46295\,
            I => \N__46288\
        );

    \I__9904\ : Span4Mux_v
    port map (
            O => \N__46292\,
            I => \N__46285\
        );

    \I__9903\ : InMux
    port map (
            O => \N__46291\,
            I => \N__46282\
        );

    \I__9902\ : Span12Mux_v
    port map (
            O => \N__46288\,
            I => \N__46279\
        );

    \I__9901\ : Span4Mux_v
    port map (
            O => \N__46285\,
            I => \N__46276\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__46282\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__9899\ : Odrv12
    port map (
            O => \N__46279\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__9898\ : Odrv4
    port map (
            O => \N__46276\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__9897\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46266\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__46266\,
            I => \N__46263\
        );

    \I__9895\ : Span4Mux_h
    port map (
            O => \N__46263\,
            I => \N__46260\
        );

    \I__9894\ : Odrv4
    port map (
            O => \N__46260\,
            I => \ppm_encoder_1.un1_init_pulses_10_8\
        );

    \I__9893\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46254\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__46254\,
            I => \N__46250\
        );

    \I__9891\ : InMux
    port map (
            O => \N__46253\,
            I => \N__46247\
        );

    \I__9890\ : Span4Mux_v
    port map (
            O => \N__46250\,
            I => \N__46242\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__46247\,
            I => \N__46242\
        );

    \I__9888\ : Span4Mux_h
    port map (
            O => \N__46242\,
            I => \N__46239\
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__46239\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__9886\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46233\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__46233\,
            I => \N__46228\
        );

    \I__9884\ : InMux
    port map (
            O => \N__46232\,
            I => \N__46225\
        );

    \I__9883\ : CascadeMux
    port map (
            O => \N__46231\,
            I => \N__46222\
        );

    \I__9882\ : Span4Mux_v
    port map (
            O => \N__46228\,
            I => \N__46219\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__46225\,
            I => \N__46216\
        );

    \I__9880\ : InMux
    port map (
            O => \N__46222\,
            I => \N__46213\
        );

    \I__9879\ : Span4Mux_h
    port map (
            O => \N__46219\,
            I => \N__46208\
        );

    \I__9878\ : Span4Mux_v
    port map (
            O => \N__46216\,
            I => \N__46208\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__46213\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__9876\ : Odrv4
    port map (
            O => \N__46208\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__9875\ : CascadeMux
    port map (
            O => \N__46203\,
            I => \N__46200\
        );

    \I__9874\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46191\
        );

    \I__9873\ : InMux
    port map (
            O => \N__46199\,
            I => \N__46191\
        );

    \I__9872\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46191\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__46191\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__9870\ : InMux
    port map (
            O => \N__46188\,
            I => \N__46185\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__46185\,
            I => \N__46182\
        );

    \I__9868\ : Span4Mux_v
    port map (
            O => \N__46182\,
            I => \N__46179\
        );

    \I__9867\ : Span4Mux_v
    port map (
            O => \N__46179\,
            I => \N__46176\
        );

    \I__9866\ : Odrv4
    port map (
            O => \N__46176\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\
        );

    \I__9865\ : InMux
    port map (
            O => \N__46173\,
            I => \N__46170\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__46170\,
            I => \N__46167\
        );

    \I__9863\ : Span4Mux_h
    port map (
            O => \N__46167\,
            I => \N__46164\
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__46164\,
            I => \ppm_encoder_1.un1_init_pulses_10_9\
        );

    \I__9861\ : InMux
    port map (
            O => \N__46161\,
            I => \N__46157\
        );

    \I__9860\ : InMux
    port map (
            O => \N__46160\,
            I => \N__46154\
        );

    \I__9859\ : LocalMux
    port map (
            O => \N__46157\,
            I => \N__46151\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__46154\,
            I => \N__46148\
        );

    \I__9857\ : Span4Mux_h
    port map (
            O => \N__46151\,
            I => \N__46143\
        );

    \I__9856\ : Span4Mux_h
    port map (
            O => \N__46148\,
            I => \N__46143\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__46143\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__9854\ : CascadeMux
    port map (
            O => \N__46140\,
            I => \N__46137\
        );

    \I__9853\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46134\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__46134\,
            I => \N__46131\
        );

    \I__9851\ : Span4Mux_h
    port map (
            O => \N__46131\,
            I => \N__46128\
        );

    \I__9850\ : Span4Mux_h
    port map (
            O => \N__46128\,
            I => \N__46123\
        );

    \I__9849\ : InMux
    port map (
            O => \N__46127\,
            I => \N__46118\
        );

    \I__9848\ : InMux
    port map (
            O => \N__46126\,
            I => \N__46118\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__46123\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__46118\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__9845\ : InMux
    port map (
            O => \N__46113\,
            I => \N__46109\
        );

    \I__9844\ : InMux
    port map (
            O => \N__46112\,
            I => \N__46105\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__46109\,
            I => \N__46102\
        );

    \I__9842\ : InMux
    port map (
            O => \N__46108\,
            I => \N__46099\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__46105\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__46102\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__46099\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__9838\ : InMux
    port map (
            O => \N__46092\,
            I => \N__46089\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__46089\,
            I => \N__46086\
        );

    \I__9836\ : Span4Mux_v
    port map (
            O => \N__46086\,
            I => \N__46083\
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__46083\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\
        );

    \I__9834\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46077\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__46077\,
            I => \ppm_encoder_1.un1_init_pulses_10_0\
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__46074\,
            I => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\
        );

    \I__9831\ : CascadeMux
    port map (
            O => \N__46071\,
            I => \N__46067\
        );

    \I__9830\ : InMux
    port map (
            O => \N__46070\,
            I => \N__46064\
        );

    \I__9829\ : InMux
    port map (
            O => \N__46067\,
            I => \N__46059\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__46064\,
            I => \N__46056\
        );

    \I__9827\ : InMux
    port map (
            O => \N__46063\,
            I => \N__46051\
        );

    \I__9826\ : InMux
    port map (
            O => \N__46062\,
            I => \N__46051\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__46059\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__9824\ : Odrv4
    port map (
            O => \N__46056\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__46051\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__9822\ : CascadeMux
    port map (
            O => \N__46044\,
            I => \N__46041\
        );

    \I__9821\ : InMux
    port map (
            O => \N__46041\,
            I => \N__46037\
        );

    \I__9820\ : InMux
    port map (
            O => \N__46040\,
            I => \N__46033\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__46037\,
            I => \N__46030\
        );

    \I__9818\ : InMux
    port map (
            O => \N__46036\,
            I => \N__46027\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__46033\,
            I => \N__46022\
        );

    \I__9816\ : Span4Mux_h
    port map (
            O => \N__46030\,
            I => \N__46022\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__46027\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__9814\ : Odrv4
    port map (
            O => \N__46022\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__9813\ : InMux
    port map (
            O => \N__46017\,
            I => \N__46014\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__46014\,
            I => \N__46011\
        );

    \I__9811\ : Span4Mux_h
    port map (
            O => \N__46011\,
            I => \N__46008\
        );

    \I__9810\ : Odrv4
    port map (
            O => \N__46008\,
            I => \ppm_encoder_1.un1_init_pulses_10_5\
        );

    \I__9809\ : InMux
    port map (
            O => \N__46005\,
            I => \N__46001\
        );

    \I__9808\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45998\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__46001\,
            I => \N__45995\
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__45998\,
            I => \N__45992\
        );

    \I__9805\ : Span4Mux_v
    port map (
            O => \N__45995\,
            I => \N__45989\
        );

    \I__9804\ : Odrv12
    port map (
            O => \N__45992\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__9803\ : Odrv4
    port map (
            O => \N__45989\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__9802\ : InMux
    port map (
            O => \N__45984\,
            I => \N__45975\
        );

    \I__9801\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45975\
        );

    \I__9800\ : InMux
    port map (
            O => \N__45982\,
            I => \N__45975\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__45975\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__9798\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45968\
        );

    \I__9797\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45965\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__45968\,
            I => \N__45960\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45960\
        );

    \I__9794\ : Span4Mux_h
    port map (
            O => \N__45960\,
            I => \N__45957\
        );

    \I__9793\ : Span4Mux_h
    port map (
            O => \N__45957\,
            I => \N__45954\
        );

    \I__9792\ : Odrv4
    port map (
            O => \N__45954\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__9791\ : InMux
    port map (
            O => \N__45951\,
            I => \N__45948\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__45948\,
            I => \N__45945\
        );

    \I__9789\ : Span4Mux_h
    port map (
            O => \N__45945\,
            I => \N__45942\
        );

    \I__9788\ : Span4Mux_v
    port map (
            O => \N__45942\,
            I => \N__45939\
        );

    \I__9787\ : Odrv4
    port map (
            O => \N__45939\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\
        );

    \I__9786\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45933\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__45933\,
            I => \N__45930\
        );

    \I__9784\ : Span4Mux_h
    port map (
            O => \N__45930\,
            I => \N__45927\
        );

    \I__9783\ : Odrv4
    port map (
            O => \N__45927\,
            I => \ppm_encoder_1.un1_init_pulses_10_7\
        );

    \I__9782\ : InMux
    port map (
            O => \N__45924\,
            I => \N__45920\
        );

    \I__9781\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45917\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__45920\,
            I => \N__45914\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__45917\,
            I => \N__45911\
        );

    \I__9778\ : Span4Mux_v
    port map (
            O => \N__45914\,
            I => \N__45908\
        );

    \I__9777\ : Span4Mux_h
    port map (
            O => \N__45911\,
            I => \N__45905\
        );

    \I__9776\ : Odrv4
    port map (
            O => \N__45908\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__9775\ : Odrv4
    port map (
            O => \N__45905\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__9774\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45897\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45894\
        );

    \I__9772\ : Span4Mux_v
    port map (
            O => \N__45894\,
            I => \N__45889\
        );

    \I__9771\ : InMux
    port map (
            O => \N__45893\,
            I => \N__45884\
        );

    \I__9770\ : InMux
    port map (
            O => \N__45892\,
            I => \N__45884\
        );

    \I__9769\ : Odrv4
    port map (
            O => \N__45889\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__45884\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__9767\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45875\
        );

    \I__9766\ : CascadeMux
    port map (
            O => \N__45878\,
            I => \N__45871\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__45875\,
            I => \N__45867\
        );

    \I__9764\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45862\
        );

    \I__9763\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45862\
        );

    \I__9762\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45859\
        );

    \I__9761\ : Span4Mux_h
    port map (
            O => \N__45867\,
            I => \N__45856\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__45862\,
            I => \ppm_encoder_1.elevatorZ0Z_0\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__45859\,
            I => \ppm_encoder_1.elevatorZ0Z_0\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__45856\,
            I => \ppm_encoder_1.elevatorZ0Z_0\
        );

    \I__9757\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45846\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__45846\,
            I => \N__45843\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__45843\,
            I => \N__45840\
        );

    \I__9754\ : Span4Mux_v
    port map (
            O => \N__45840\,
            I => \N__45837\
        );

    \I__9753\ : Odrv4
    port map (
            O => \N__45837\,
            I => \ppm_encoder_1.un1_init_pulses_10_6\
        );

    \I__9752\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45830\
        );

    \I__9751\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45827\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45822\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__45827\,
            I => \N__45822\
        );

    \I__9748\ : Span4Mux_v
    port map (
            O => \N__45822\,
            I => \N__45819\
        );

    \I__9747\ : Odrv4
    port map (
            O => \N__45819\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__9746\ : CascadeMux
    port map (
            O => \N__45816\,
            I => \N__45813\
        );

    \I__9745\ : InMux
    port map (
            O => \N__45813\,
            I => \N__45810\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__45807\,
            I => \N__45804\
        );

    \I__9742\ : Span4Mux_v
    port map (
            O => \N__45804\,
            I => \N__45801\
        );

    \I__9741\ : Odrv4
    port map (
            O => \N__45801\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3\
        );

    \I__9740\ : CascadeMux
    port map (
            O => \N__45798\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_\
        );

    \I__9739\ : InMux
    port map (
            O => \N__45795\,
            I => \N__45792\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__45792\,
            I => \N__45789\
        );

    \I__9737\ : Span4Mux_v
    port map (
            O => \N__45789\,
            I => \N__45786\
        );

    \I__9736\ : Odrv4
    port map (
            O => \N__45786\,
            I => \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15\
        );

    \I__9735\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45780\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__45780\,
            I => \N__45775\
        );

    \I__9733\ : InMux
    port map (
            O => \N__45779\,
            I => \N__45772\
        );

    \I__9732\ : InMux
    port map (
            O => \N__45778\,
            I => \N__45769\
        );

    \I__9731\ : Span4Mux_v
    port map (
            O => \N__45775\,
            I => \N__45766\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__45772\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__45769\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__9728\ : Odrv4
    port map (
            O => \N__45766\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__9727\ : InMux
    port map (
            O => \N__45759\,
            I => \N__45756\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__45756\,
            I => \N__45753\
        );

    \I__9725\ : Span12Mux_h
    port map (
            O => \N__45753\,
            I => \N__45748\
        );

    \I__9724\ : InMux
    port map (
            O => \N__45752\,
            I => \N__45745\
        );

    \I__9723\ : InMux
    port map (
            O => \N__45751\,
            I => \N__45742\
        );

    \I__9722\ : Odrv12
    port map (
            O => \N__45748\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__45745\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__45742\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__45735\,
            I => \N__45732\
        );

    \I__9718\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45729\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__45729\,
            I => \pid_side.m26_e_5\
        );

    \I__9716\ : CascadeMux
    port map (
            O => \N__45726\,
            I => \pid_side.pid_prereg_esr_RNIGJDR1Z0Z_10_cascade_\
        );

    \I__9715\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45720\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__45720\,
            I => \pid_side.m18_s_4\
        );

    \I__9713\ : CascadeMux
    port map (
            O => \N__45717\,
            I => \pid_side.pid_prereg_esr_RNIQBAH2Z0Z_23_cascade_\
        );

    \I__9712\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45711\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__45711\,
            I => \N__45708\
        );

    \I__9710\ : Odrv4
    port map (
            O => \N__45708\,
            I => \pid_side.un1_reset_0_i_sn\
        );

    \I__9709\ : CascadeMux
    port map (
            O => \N__45705\,
            I => \pid_side.i19_mux_cascade_\
        );

    \I__9708\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45691\
        );

    \I__9707\ : InMux
    port map (
            O => \N__45701\,
            I => \N__45688\
        );

    \I__9706\ : InMux
    port map (
            O => \N__45700\,
            I => \N__45675\
        );

    \I__9705\ : InMux
    port map (
            O => \N__45699\,
            I => \N__45675\
        );

    \I__9704\ : InMux
    port map (
            O => \N__45698\,
            I => \N__45675\
        );

    \I__9703\ : InMux
    port map (
            O => \N__45697\,
            I => \N__45675\
        );

    \I__9702\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45675\
        );

    \I__9701\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45675\
        );

    \I__9700\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45672\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__45691\,
            I => \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__45688\,
            I => \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__45675\,
            I => \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__45672\,
            I => \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12\
        );

    \I__9695\ : InMux
    port map (
            O => \N__45663\,
            I => \N__45658\
        );

    \I__9694\ : InMux
    port map (
            O => \N__45662\,
            I => \N__45653\
        );

    \I__9693\ : InMux
    port map (
            O => \N__45661\,
            I => \N__45653\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__45658\,
            I => \pid_side.N_11_0\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__45653\,
            I => \pid_side.N_11_0\
        );

    \I__9690\ : CascadeMux
    port map (
            O => \N__45648\,
            I => \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12_cascade_\
        );

    \I__9689\ : InMux
    port map (
            O => \N__45645\,
            I => \N__45638\
        );

    \I__9688\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45638\
        );

    \I__9687\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45635\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__45638\,
            I => \N__45632\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__45635\,
            I => \pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10\
        );

    \I__9684\ : Odrv4
    port map (
            O => \N__45632\,
            I => \pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10\
        );

    \I__9683\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45618\
        );

    \I__9682\ : InMux
    port map (
            O => \N__45626\,
            I => \N__45618\
        );

    \I__9681\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45618\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__45618\,
            I => \N__45615\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__45615\,
            I => \N__45610\
        );

    \I__9678\ : InMux
    port map (
            O => \N__45614\,
            I => \N__45607\
        );

    \I__9677\ : InMux
    port map (
            O => \N__45613\,
            I => \N__45604\
        );

    \I__9676\ : Odrv4
    port map (
            O => \N__45610\,
            I => \pid_side.N_82_mux\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__45607\,
            I => \pid_side.N_82_mux\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__45604\,
            I => \pid_side.N_82_mux\
        );

    \I__9673\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45594\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__45594\,
            I => \N__45591\
        );

    \I__9671\ : Span4Mux_h
    port map (
            O => \N__45591\,
            I => \N__45587\
        );

    \I__9670\ : InMux
    port map (
            O => \N__45590\,
            I => \N__45584\
        );

    \I__9669\ : Span4Mux_v
    port map (
            O => \N__45587\,
            I => \N__45581\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__45584\,
            I => \N__45578\
        );

    \I__9667\ : Span4Mux_h
    port map (
            O => \N__45581\,
            I => \N__45575\
        );

    \I__9666\ : Odrv4
    port map (
            O => \N__45578\,
            I => side_order_12
        );

    \I__9665\ : Odrv4
    port map (
            O => \N__45575\,
            I => side_order_12
        );

    \I__9664\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45567\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__45567\,
            I => \N__45564\
        );

    \I__9662\ : Odrv4
    port map (
            O => \N__45564\,
            I => \ppm_encoder_1.un2_throttle_iv_0_0\
        );

    \I__9661\ : CascadeMux
    port map (
            O => \N__45561\,
            I => \N__45554\
        );

    \I__9660\ : CascadeMux
    port map (
            O => \N__45560\,
            I => \N__45550\
        );

    \I__9659\ : InMux
    port map (
            O => \N__45559\,
            I => \N__45547\
        );

    \I__9658\ : CascadeMux
    port map (
            O => \N__45558\,
            I => \N__45542\
        );

    \I__9657\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45539\
        );

    \I__9656\ : InMux
    port map (
            O => \N__45554\,
            I => \N__45536\
        );

    \I__9655\ : InMux
    port map (
            O => \N__45553\,
            I => \N__45533\
        );

    \I__9654\ : InMux
    port map (
            O => \N__45550\,
            I => \N__45529\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__45547\,
            I => \N__45526\
        );

    \I__9652\ : InMux
    port map (
            O => \N__45546\,
            I => \N__45523\
        );

    \I__9651\ : CascadeMux
    port map (
            O => \N__45545\,
            I => \N__45520\
        );

    \I__9650\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45517\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__45539\,
            I => \N__45510\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__45536\,
            I => \N__45505\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__45533\,
            I => \N__45505\
        );

    \I__9646\ : CascadeMux
    port map (
            O => \N__45532\,
            I => \N__45500\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__45529\,
            I => \N__45493\
        );

    \I__9644\ : Span4Mux_h
    port map (
            O => \N__45526\,
            I => \N__45493\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__45523\,
            I => \N__45493\
        );

    \I__9642\ : InMux
    port map (
            O => \N__45520\,
            I => \N__45490\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__45517\,
            I => \N__45487\
        );

    \I__9640\ : InMux
    port map (
            O => \N__45516\,
            I => \N__45484\
        );

    \I__9639\ : CascadeMux
    port map (
            O => \N__45515\,
            I => \N__45480\
        );

    \I__9638\ : CascadeMux
    port map (
            O => \N__45514\,
            I => \N__45477\
        );

    \I__9637\ : InMux
    port map (
            O => \N__45513\,
            I => \N__45474\
        );

    \I__9636\ : Span4Mux_v
    port map (
            O => \N__45510\,
            I => \N__45469\
        );

    \I__9635\ : Span4Mux_v
    port map (
            O => \N__45505\,
            I => \N__45469\
        );

    \I__9634\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45464\
        );

    \I__9633\ : InMux
    port map (
            O => \N__45503\,
            I => \N__45464\
        );

    \I__9632\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45461\
        );

    \I__9631\ : Span4Mux_v
    port map (
            O => \N__45493\,
            I => \N__45452\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__45490\,
            I => \N__45452\
        );

    \I__9629\ : Span4Mux_h
    port map (
            O => \N__45487\,
            I => \N__45452\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__45484\,
            I => \N__45452\
        );

    \I__9627\ : InMux
    port map (
            O => \N__45483\,
            I => \N__45449\
        );

    \I__9626\ : InMux
    port map (
            O => \N__45480\,
            I => \N__45444\
        );

    \I__9625\ : InMux
    port map (
            O => \N__45477\,
            I => \N__45444\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__45474\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__9623\ : Odrv4
    port map (
            O => \N__45469\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__45464\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__45461\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__9620\ : Odrv4
    port map (
            O => \N__45452\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__45449\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__45444\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__9617\ : InMux
    port map (
            O => \N__45429\,
            I => \N__45425\
        );

    \I__9616\ : InMux
    port map (
            O => \N__45428\,
            I => \N__45422\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__45425\,
            I => \N__45419\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__45422\,
            I => \N__45416\
        );

    \I__9613\ : Span12Mux_h
    port map (
            O => \N__45419\,
            I => \N__45413\
        );

    \I__9612\ : Span4Mux_h
    port map (
            O => \N__45416\,
            I => \N__45410\
        );

    \I__9611\ : Odrv12
    port map (
            O => \N__45413\,
            I => front_order_0
        );

    \I__9610\ : Odrv4
    port map (
            O => \N__45410\,
            I => front_order_0
        );

    \I__9609\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45391\
        );

    \I__9608\ : CascadeMux
    port map (
            O => \N__45404\,
            I => \N__45382\
        );

    \I__9607\ : CascadeMux
    port map (
            O => \N__45403\,
            I => \N__45377\
        );

    \I__9606\ : CascadeMux
    port map (
            O => \N__45402\,
            I => \N__45367\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__45401\,
            I => \N__45364\
        );

    \I__9604\ : CascadeMux
    port map (
            O => \N__45400\,
            I => \N__45359\
        );

    \I__9603\ : CascadeMux
    port map (
            O => \N__45399\,
            I => \N__45355\
        );

    \I__9602\ : CascadeMux
    port map (
            O => \N__45398\,
            I => \N__45351\
        );

    \I__9601\ : CascadeMux
    port map (
            O => \N__45397\,
            I => \N__45348\
        );

    \I__9600\ : CascadeMux
    port map (
            O => \N__45396\,
            I => \N__45345\
        );

    \I__9599\ : CascadeMux
    port map (
            O => \N__45395\,
            I => \N__45337\
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__45394\,
            I => \N__45334\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__45391\,
            I => \N__45330\
        );

    \I__9596\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45325\
        );

    \I__9595\ : InMux
    port map (
            O => \N__45389\,
            I => \N__45325\
        );

    \I__9594\ : CascadeMux
    port map (
            O => \N__45388\,
            I => \N__45322\
        );

    \I__9593\ : CascadeMux
    port map (
            O => \N__45387\,
            I => \N__45318\
        );

    \I__9592\ : CascadeMux
    port map (
            O => \N__45386\,
            I => \N__45315\
        );

    \I__9591\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45311\
        );

    \I__9590\ : InMux
    port map (
            O => \N__45382\,
            I => \N__45306\
        );

    \I__9589\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45306\
        );

    \I__9588\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45299\
        );

    \I__9587\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45299\
        );

    \I__9586\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45299\
        );

    \I__9585\ : CascadeMux
    port map (
            O => \N__45375\,
            I => \N__45291\
        );

    \I__9584\ : CascadeMux
    port map (
            O => \N__45374\,
            I => \N__45288\
        );

    \I__9583\ : CascadeMux
    port map (
            O => \N__45373\,
            I => \N__45285\
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__45372\,
            I => \N__45282\
        );

    \I__9581\ : CascadeMux
    port map (
            O => \N__45371\,
            I => \N__45279\
        );

    \I__9580\ : CascadeMux
    port map (
            O => \N__45370\,
            I => \N__45276\
        );

    \I__9579\ : InMux
    port map (
            O => \N__45367\,
            I => \N__45273\
        );

    \I__9578\ : InMux
    port map (
            O => \N__45364\,
            I => \N__45270\
        );

    \I__9577\ : InMux
    port map (
            O => \N__45363\,
            I => \N__45267\
        );

    \I__9576\ : InMux
    port map (
            O => \N__45362\,
            I => \N__45262\
        );

    \I__9575\ : InMux
    port map (
            O => \N__45359\,
            I => \N__45262\
        );

    \I__9574\ : InMux
    port map (
            O => \N__45358\,
            I => \N__45257\
        );

    \I__9573\ : InMux
    port map (
            O => \N__45355\,
            I => \N__45257\
        );

    \I__9572\ : InMux
    port map (
            O => \N__45354\,
            I => \N__45252\
        );

    \I__9571\ : InMux
    port map (
            O => \N__45351\,
            I => \N__45252\
        );

    \I__9570\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45241\
        );

    \I__9569\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45241\
        );

    \I__9568\ : InMux
    port map (
            O => \N__45344\,
            I => \N__45241\
        );

    \I__9567\ : InMux
    port map (
            O => \N__45343\,
            I => \N__45241\
        );

    \I__9566\ : InMux
    port map (
            O => \N__45342\,
            I => \N__45241\
        );

    \I__9565\ : InMux
    port map (
            O => \N__45341\,
            I => \N__45230\
        );

    \I__9564\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45230\
        );

    \I__9563\ : InMux
    port map (
            O => \N__45337\,
            I => \N__45230\
        );

    \I__9562\ : InMux
    port map (
            O => \N__45334\,
            I => \N__45230\
        );

    \I__9561\ : InMux
    port map (
            O => \N__45333\,
            I => \N__45230\
        );

    \I__9560\ : Span4Mux_v
    port map (
            O => \N__45330\,
            I => \N__45225\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__45325\,
            I => \N__45225\
        );

    \I__9558\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45222\
        );

    \I__9557\ : InMux
    port map (
            O => \N__45321\,
            I => \N__45215\
        );

    \I__9556\ : InMux
    port map (
            O => \N__45318\,
            I => \N__45215\
        );

    \I__9555\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45215\
        );

    \I__9554\ : CascadeMux
    port map (
            O => \N__45314\,
            I => \N__45212\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__45311\,
            I => \N__45209\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__45306\,
            I => \N__45204\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__45299\,
            I => \N__45204\
        );

    \I__9550\ : CascadeMux
    port map (
            O => \N__45298\,
            I => \N__45197\
        );

    \I__9549\ : CascadeMux
    port map (
            O => \N__45297\,
            I => \N__45194\
        );

    \I__9548\ : CascadeMux
    port map (
            O => \N__45296\,
            I => \N__45191\
        );

    \I__9547\ : CascadeMux
    port map (
            O => \N__45295\,
            I => \N__45187\
        );

    \I__9546\ : InMux
    port map (
            O => \N__45294\,
            I => \N__45181\
        );

    \I__9545\ : InMux
    port map (
            O => \N__45291\,
            I => \N__45181\
        );

    \I__9544\ : InMux
    port map (
            O => \N__45288\,
            I => \N__45174\
        );

    \I__9543\ : InMux
    port map (
            O => \N__45285\,
            I => \N__45174\
        );

    \I__9542\ : InMux
    port map (
            O => \N__45282\,
            I => \N__45174\
        );

    \I__9541\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45169\
        );

    \I__9540\ : InMux
    port map (
            O => \N__45276\,
            I => \N__45169\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__45273\,
            I => \N__45164\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__45270\,
            I => \N__45164\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__45267\,
            I => \N__45159\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__45262\,
            I => \N__45159\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__45257\,
            I => \N__45144\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__45252\,
            I => \N__45144\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__45241\,
            I => \N__45144\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__45230\,
            I => \N__45144\
        );

    \I__9531\ : Span4Mux_h
    port map (
            O => \N__45225\,
            I => \N__45144\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__45222\,
            I => \N__45144\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__45215\,
            I => \N__45144\
        );

    \I__9528\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45141\
        );

    \I__9527\ : Span4Mux_h
    port map (
            O => \N__45209\,
            I => \N__45136\
        );

    \I__9526\ : Span4Mux_v
    port map (
            O => \N__45204\,
            I => \N__45136\
        );

    \I__9525\ : InMux
    port map (
            O => \N__45203\,
            I => \N__45133\
        );

    \I__9524\ : CascadeMux
    port map (
            O => \N__45202\,
            I => \N__45129\
        );

    \I__9523\ : CascadeMux
    port map (
            O => \N__45201\,
            I => \N__45126\
        );

    \I__9522\ : InMux
    port map (
            O => \N__45200\,
            I => \N__45115\
        );

    \I__9521\ : InMux
    port map (
            O => \N__45197\,
            I => \N__45115\
        );

    \I__9520\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45115\
        );

    \I__9519\ : InMux
    port map (
            O => \N__45191\,
            I => \N__45115\
        );

    \I__9518\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45115\
        );

    \I__9517\ : InMux
    port map (
            O => \N__45187\,
            I => \N__45110\
        );

    \I__9516\ : InMux
    port map (
            O => \N__45186\,
            I => \N__45110\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__45181\,
            I => \N__45107\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__45174\,
            I => \N__45098\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__45169\,
            I => \N__45098\
        );

    \I__9512\ : Span4Mux_v
    port map (
            O => \N__45164\,
            I => \N__45098\
        );

    \I__9511\ : Span4Mux_v
    port map (
            O => \N__45159\,
            I => \N__45098\
        );

    \I__9510\ : Span4Mux_v
    port map (
            O => \N__45144\,
            I => \N__45095\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__45141\,
            I => \N__45088\
        );

    \I__9508\ : Span4Mux_h
    port map (
            O => \N__45136\,
            I => \N__45088\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__45133\,
            I => \N__45088\
        );

    \I__9506\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45081\
        );

    \I__9505\ : InMux
    port map (
            O => \N__45129\,
            I => \N__45081\
        );

    \I__9504\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45081\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__45115\,
            I => \N__45076\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__45110\,
            I => \N__45076\
        );

    \I__9501\ : Span4Mux_v
    port map (
            O => \N__45107\,
            I => \N__45071\
        );

    \I__9500\ : Span4Mux_v
    port map (
            O => \N__45098\,
            I => \N__45071\
        );

    \I__9499\ : Span4Mux_v
    port map (
            O => \N__45095\,
            I => \N__45066\
        );

    \I__9498\ : Span4Mux_v
    port map (
            O => \N__45088\,
            I => \N__45066\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__45081\,
            I => pid_altitude_dv
        );

    \I__9496\ : Odrv12
    port map (
            O => \N__45076\,
            I => pid_altitude_dv
        );

    \I__9495\ : Odrv4
    port map (
            O => \N__45071\,
            I => pid_altitude_dv
        );

    \I__9494\ : Odrv4
    port map (
            O => \N__45066\,
            I => pid_altitude_dv
        );

    \I__9493\ : InMux
    port map (
            O => \N__45057\,
            I => \N__45053\
        );

    \I__9492\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45050\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__45053\,
            I => \N__45047\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__45050\,
            I => \N__45044\
        );

    \I__9489\ : Span12Mux_h
    port map (
            O => \N__45047\,
            I => \N__45041\
        );

    \I__9488\ : Span12Mux_s9_h
    port map (
            O => \N__45044\,
            I => \N__45038\
        );

    \I__9487\ : Odrv12
    port map (
            O => \N__45041\,
            I => \pid_front.error_d_reg_prevZ0Z_14\
        );

    \I__9486\ : Odrv12
    port map (
            O => \N__45038\,
            I => \pid_front.error_d_reg_prevZ0Z_14\
        );

    \I__9485\ : InMux
    port map (
            O => \N__45033\,
            I => \N__45029\
        );

    \I__9484\ : CascadeMux
    port map (
            O => \N__45032\,
            I => \N__45026\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__45029\,
            I => \N__45022\
        );

    \I__9482\ : InMux
    port map (
            O => \N__45026\,
            I => \N__45017\
        );

    \I__9481\ : InMux
    port map (
            O => \N__45025\,
            I => \N__45017\
        );

    \I__9480\ : Odrv12
    port map (
            O => \N__45022\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__45017\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__9478\ : CascadeMux
    port map (
            O => \N__45012\,
            I => \N__45008\
        );

    \I__9477\ : CascadeMux
    port map (
            O => \N__45011\,
            I => \N__45005\
        );

    \I__9476\ : InMux
    port map (
            O => \N__45008\,
            I => \N__45002\
        );

    \I__9475\ : InMux
    port map (
            O => \N__45005\,
            I => \N__44999\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__45002\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__44999\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__9472\ : InMux
    port map (
            O => \N__44994\,
            I => \N__44991\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__44991\,
            I => \pid_side.m32_1\
        );

    \I__9470\ : InMux
    port map (
            O => \N__44988\,
            I => \N__44985\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__44985\,
            I => \N__44981\
        );

    \I__9468\ : InMux
    port map (
            O => \N__44984\,
            I => \N__44975\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__44981\,
            I => \N__44972\
        );

    \I__9466\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44967\
        );

    \I__9465\ : InMux
    port map (
            O => \N__44979\,
            I => \N__44961\
        );

    \I__9464\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44961\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__44975\,
            I => \N__44958\
        );

    \I__9462\ : Span4Mux_h
    port map (
            O => \N__44972\,
            I => \N__44955\
        );

    \I__9461\ : IoInMux
    port map (
            O => \N__44971\,
            I => \N__44952\
        );

    \I__9460\ : InMux
    port map (
            O => \N__44970\,
            I => \N__44947\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__44967\,
            I => \N__44944\
        );

    \I__9458\ : InMux
    port map (
            O => \N__44966\,
            I => \N__44941\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44938\
        );

    \I__9456\ : Span4Mux_v
    port map (
            O => \N__44958\,
            I => \N__44935\
        );

    \I__9455\ : Span4Mux_v
    port map (
            O => \N__44955\,
            I => \N__44932\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__44952\,
            I => \N__44929\
        );

    \I__9453\ : InMux
    port map (
            O => \N__44951\,
            I => \N__44925\
        );

    \I__9452\ : InMux
    port map (
            O => \N__44950\,
            I => \N__44922\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__44947\,
            I => \N__44919\
        );

    \I__9450\ : Span4Mux_h
    port map (
            O => \N__44944\,
            I => \N__44916\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__44941\,
            I => \N__44913\
        );

    \I__9448\ : Span4Mux_v
    port map (
            O => \N__44938\,
            I => \N__44910\
        );

    \I__9447\ : Span4Mux_v
    port map (
            O => \N__44935\,
            I => \N__44905\
        );

    \I__9446\ : Span4Mux_v
    port map (
            O => \N__44932\,
            I => \N__44905\
        );

    \I__9445\ : Span4Mux_s3_v
    port map (
            O => \N__44929\,
            I => \N__44902\
        );

    \I__9444\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44899\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__44925\,
            I => \N__44896\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__44922\,
            I => \N__44891\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__44919\,
            I => \N__44891\
        );

    \I__9440\ : Span4Mux_h
    port map (
            O => \N__44916\,
            I => \N__44888\
        );

    \I__9439\ : Span4Mux_v
    port map (
            O => \N__44913\,
            I => \N__44881\
        );

    \I__9438\ : Span4Mux_h
    port map (
            O => \N__44910\,
            I => \N__44881\
        );

    \I__9437\ : Span4Mux_v
    port map (
            O => \N__44905\,
            I => \N__44881\
        );

    \I__9436\ : Span4Mux_h
    port map (
            O => \N__44902\,
            I => \N__44878\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__44899\,
            I => reset_system
        );

    \I__9434\ : Odrv4
    port map (
            O => \N__44896\,
            I => reset_system
        );

    \I__9433\ : Odrv4
    port map (
            O => \N__44891\,
            I => reset_system
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__44888\,
            I => reset_system
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__44881\,
            I => reset_system
        );

    \I__9430\ : Odrv4
    port map (
            O => \N__44878\,
            I => reset_system
        );

    \I__9429\ : CascadeMux
    port map (
            O => \N__44865\,
            I => \pid_side.m26_e_5_cascade_\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__44862\,
            I => \pid_side.N_11_0_cascade_\
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__44859\,
            I => \N__44855\
        );

    \I__9426\ : InMux
    port map (
            O => \N__44858\,
            I => \N__44847\
        );

    \I__9425\ : InMux
    port map (
            O => \N__44855\,
            I => \N__44847\
        );

    \I__9424\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44847\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__44847\,
            I => \N__44844\
        );

    \I__9422\ : Span4Mux_v
    port map (
            O => \N__44844\,
            I => \N__44840\
        );

    \I__9421\ : InMux
    port map (
            O => \N__44843\,
            I => \N__44837\
        );

    \I__9420\ : Odrv4
    port map (
            O => \N__44840\,
            I => \pid_side.pid_prereg_esr_RNILRSP2Z0Z_5\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__44837\,
            I => \pid_side.pid_prereg_esr_RNILRSP2Z0Z_5\
        );

    \I__9418\ : InMux
    port map (
            O => \N__44832\,
            I => \N__44823\
        );

    \I__9417\ : InMux
    port map (
            O => \N__44831\,
            I => \N__44823\
        );

    \I__9416\ : InMux
    port map (
            O => \N__44830\,
            I => \N__44823\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__44823\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__9414\ : InMux
    port map (
            O => \N__44820\,
            I => \N__44817\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__44817\,
            I => \N__44813\
        );

    \I__9412\ : InMux
    port map (
            O => \N__44816\,
            I => \N__44810\
        );

    \I__9411\ : Span4Mux_v
    port map (
            O => \N__44813\,
            I => \N__44807\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__44810\,
            I => \N__44804\
        );

    \I__9409\ : Span4Mux_h
    port map (
            O => \N__44807\,
            I => \N__44801\
        );

    \I__9408\ : Span4Mux_v
    port map (
            O => \N__44804\,
            I => \N__44798\
        );

    \I__9407\ : Span4Mux_v
    port map (
            O => \N__44801\,
            I => \N__44795\
        );

    \I__9406\ : Span4Mux_v
    port map (
            O => \N__44798\,
            I => \N__44792\
        );

    \I__9405\ : Odrv4
    port map (
            O => \N__44795\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__9404\ : Odrv4
    port map (
            O => \N__44792\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__9403\ : InMux
    port map (
            O => \N__44787\,
            I => \N__44784\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__44784\,
            I => \N__44781\
        );

    \I__9401\ : Odrv4
    port map (
            O => \N__44781\,
            I => \ppm_encoder_1.un1_init_pulses_10_15\
        );

    \I__9400\ : InMux
    port map (
            O => \N__44778\,
            I => \N__44775\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__44775\,
            I => \ppm_encoder_1.un1_init_pulses_10_16\
        );

    \I__9398\ : InMux
    port map (
            O => \N__44772\,
            I => \N__44766\
        );

    \I__9397\ : InMux
    port map (
            O => \N__44771\,
            I => \N__44766\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__44766\,
            I => \N__44762\
        );

    \I__9395\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44759\
        );

    \I__9394\ : Span4Mux_v
    port map (
            O => \N__44762\,
            I => \N__44756\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__44759\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__44756\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__9391\ : InMux
    port map (
            O => \N__44751\,
            I => \N__44748\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__44748\,
            I => \N__44745\
        );

    \I__9389\ : Span4Mux_h
    port map (
            O => \N__44745\,
            I => \N__44742\
        );

    \I__9388\ : Odrv4
    port map (
            O => \N__44742\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\
        );

    \I__9387\ : InMux
    port map (
            O => \N__44739\,
            I => \N__44736\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__44736\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\
        );

    \I__9385\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44730\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__44730\,
            I => \ppm_encoder_1.pulses2countZ0Z_14\
        );

    \I__9383\ : CascadeMux
    port map (
            O => \N__44727\,
            I => \N__44722\
        );

    \I__9382\ : InMux
    port map (
            O => \N__44726\,
            I => \N__44717\
        );

    \I__9381\ : InMux
    port map (
            O => \N__44725\,
            I => \N__44714\
        );

    \I__9380\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44707\
        );

    \I__9379\ : InMux
    port map (
            O => \N__44721\,
            I => \N__44707\
        );

    \I__9378\ : InMux
    port map (
            O => \N__44720\,
            I => \N__44707\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__44717\,
            I => \N__44698\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__44714\,
            I => \N__44698\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__44707\,
            I => \N__44695\
        );

    \I__9374\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44686\
        );

    \I__9373\ : InMux
    port map (
            O => \N__44705\,
            I => \N__44686\
        );

    \I__9372\ : InMux
    port map (
            O => \N__44704\,
            I => \N__44686\
        );

    \I__9371\ : InMux
    port map (
            O => \N__44703\,
            I => \N__44686\
        );

    \I__9370\ : Span4Mux_v
    port map (
            O => \N__44698\,
            I => \N__44678\
        );

    \I__9369\ : Span4Mux_v
    port map (
            O => \N__44695\,
            I => \N__44675\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__44686\,
            I => \N__44672\
        );

    \I__9367\ : InMux
    port map (
            O => \N__44685\,
            I => \N__44661\
        );

    \I__9366\ : InMux
    port map (
            O => \N__44684\,
            I => \N__44661\
        );

    \I__9365\ : InMux
    port map (
            O => \N__44683\,
            I => \N__44661\
        );

    \I__9364\ : InMux
    port map (
            O => \N__44682\,
            I => \N__44661\
        );

    \I__9363\ : InMux
    port map (
            O => \N__44681\,
            I => \N__44661\
        );

    \I__9362\ : Span4Mux_v
    port map (
            O => \N__44678\,
            I => \N__44657\
        );

    \I__9361\ : Sp12to4
    port map (
            O => \N__44675\,
            I => \N__44650\
        );

    \I__9360\ : Sp12to4
    port map (
            O => \N__44672\,
            I => \N__44650\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__44661\,
            I => \N__44650\
        );

    \I__9358\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44647\
        );

    \I__9357\ : Odrv4
    port map (
            O => \N__44657\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__9356\ : Odrv12
    port map (
            O => \N__44650\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__44647\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__9354\ : InMux
    port map (
            O => \N__44640\,
            I => \N__44637\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__44637\,
            I => \N__44634\
        );

    \I__9352\ : Odrv12
    port map (
            O => \N__44634\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\
        );

    \I__9351\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44628\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__44628\,
            I => \N__44625\
        );

    \I__9349\ : Odrv12
    port map (
            O => \N__44625\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\
        );

    \I__9348\ : CascadeMux
    port map (
            O => \N__44622\,
            I => \N__44619\
        );

    \I__9347\ : InMux
    port map (
            O => \N__44619\,
            I => \N__44616\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__44616\,
            I => \ppm_encoder_1.pulses2countZ0Z_3\
        );

    \I__9345\ : CEMux
    port map (
            O => \N__44613\,
            I => \N__44609\
        );

    \I__9344\ : CEMux
    port map (
            O => \N__44612\,
            I => \N__44606\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__44609\,
            I => \N__44603\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__44606\,
            I => \N__44599\
        );

    \I__9341\ : Span4Mux_h
    port map (
            O => \N__44603\,
            I => \N__44596\
        );

    \I__9340\ : CEMux
    port map (
            O => \N__44602\,
            I => \N__44593\
        );

    \I__9339\ : Span4Mux_v
    port map (
            O => \N__44599\,
            I => \N__44589\
        );

    \I__9338\ : Span4Mux_v
    port map (
            O => \N__44596\,
            I => \N__44584\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__44593\,
            I => \N__44584\
        );

    \I__9336\ : CEMux
    port map (
            O => \N__44592\,
            I => \N__44581\
        );

    \I__9335\ : Span4Mux_h
    port map (
            O => \N__44589\,
            I => \N__44577\
        );

    \I__9334\ : Span4Mux_v
    port map (
            O => \N__44584\,
            I => \N__44572\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__44581\,
            I => \N__44572\
        );

    \I__9332\ : CEMux
    port map (
            O => \N__44580\,
            I => \N__44569\
        );

    \I__9331\ : Span4Mux_v
    port map (
            O => \N__44577\,
            I => \N__44566\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__44572\,
            I => \N__44563\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__44569\,
            I => \N__44560\
        );

    \I__9328\ : Odrv4
    port map (
            O => \N__44566\,
            I => \ppm_encoder_1.N_2150_0\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__44563\,
            I => \ppm_encoder_1.N_2150_0\
        );

    \I__9326\ : Odrv12
    port map (
            O => \N__44560\,
            I => \ppm_encoder_1.N_2150_0\
        );

    \I__9325\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44548\
        );

    \I__9324\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44545\
        );

    \I__9323\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44542\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__44548\,
            I => \N__44539\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__44545\,
            I => \N__44536\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__44542\,
            I => \N__44531\
        );

    \I__9319\ : Span4Mux_v
    port map (
            O => \N__44539\,
            I => \N__44531\
        );

    \I__9318\ : Span4Mux_h
    port map (
            O => \N__44536\,
            I => \N__44528\
        );

    \I__9317\ : Odrv4
    port map (
            O => \N__44531\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__9316\ : Odrv4
    port map (
            O => \N__44528\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__9315\ : InMux
    port map (
            O => \N__44523\,
            I => \N__44520\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__44520\,
            I => \N__44515\
        );

    \I__9313\ : InMux
    port map (
            O => \N__44519\,
            I => \N__44512\
        );

    \I__9312\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44509\
        );

    \I__9311\ : Span4Mux_h
    port map (
            O => \N__44515\,
            I => \N__44506\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__44512\,
            I => \N__44503\
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__44509\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__9308\ : Odrv4
    port map (
            O => \N__44506\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__44503\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__44496\,
            I => \N__44493\
        );

    \I__9305\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44488\
        );

    \I__9304\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44485\
        );

    \I__9303\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44482\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__44488\,
            I => \N__44479\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__44485\,
            I => \N__44476\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__44482\,
            I => \N__44471\
        );

    \I__9299\ : Span4Mux_v
    port map (
            O => \N__44479\,
            I => \N__44471\
        );

    \I__9298\ : Span4Mux_h
    port map (
            O => \N__44476\,
            I => \N__44468\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__44471\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__9296\ : Odrv4
    port map (
            O => \N__44468\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__9295\ : InMux
    port map (
            O => \N__44463\,
            I => \N__44460\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__44460\,
            I => \N__44456\
        );

    \I__9293\ : InMux
    port map (
            O => \N__44459\,
            I => \N__44452\
        );

    \I__9292\ : Span4Mux_v
    port map (
            O => \N__44456\,
            I => \N__44449\
        );

    \I__9291\ : InMux
    port map (
            O => \N__44455\,
            I => \N__44446\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__44452\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__9289\ : Odrv4
    port map (
            O => \N__44449\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__44446\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__9287\ : InMux
    port map (
            O => \N__44439\,
            I => \N__44433\
        );

    \I__9286\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44433\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__44433\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\
        );

    \I__9284\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44427\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__44427\,
            I => \ppm_encoder_1.un1_init_pulses_10_4\
        );

    \I__9282\ : InMux
    port map (
            O => \N__44424\,
            I => \N__44421\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__44421\,
            I => \N__44418\
        );

    \I__9280\ : Span4Mux_v
    port map (
            O => \N__44418\,
            I => \N__44414\
        );

    \I__9279\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44411\
        );

    \I__9278\ : Odrv4
    port map (
            O => \N__44414\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__44411\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__9276\ : InMux
    port map (
            O => \N__44406\,
            I => \N__44403\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__44403\,
            I => \ppm_encoder_1.un1_init_pulses_10_13\
        );

    \I__9274\ : InMux
    port map (
            O => \N__44400\,
            I => \N__44397\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__44397\,
            I => \N__44394\
        );

    \I__9272\ : Span4Mux_h
    port map (
            O => \N__44394\,
            I => \N__44390\
        );

    \I__9271\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44387\
        );

    \I__9270\ : Odrv4
    port map (
            O => \N__44390\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__44387\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__9268\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44379\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__44379\,
            I => \ppm_encoder_1.un1_init_pulses_10_18\
        );

    \I__9266\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44373\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__44373\,
            I => \N__44369\
        );

    \I__9264\ : InMux
    port map (
            O => \N__44372\,
            I => \N__44366\
        );

    \I__9263\ : Span4Mux_h
    port map (
            O => \N__44369\,
            I => \N__44362\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__44366\,
            I => \N__44359\
        );

    \I__9261\ : InMux
    port map (
            O => \N__44365\,
            I => \N__44356\
        );

    \I__9260\ : Sp12to4
    port map (
            O => \N__44362\,
            I => \N__44351\
        );

    \I__9259\ : Sp12to4
    port map (
            O => \N__44359\,
            I => \N__44351\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__44356\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__9257\ : Odrv12
    port map (
            O => \N__44351\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__9256\ : InMux
    port map (
            O => \N__44346\,
            I => \N__44343\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__44343\,
            I => \N__44340\
        );

    \I__9254\ : Span4Mux_h
    port map (
            O => \N__44340\,
            I => \N__44337\
        );

    \I__9253\ : Odrv4
    port map (
            O => \N__44337\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\
        );

    \I__9252\ : InMux
    port map (
            O => \N__44334\,
            I => \N__44331\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__44331\,
            I => \N__44328\
        );

    \I__9250\ : Odrv4
    port map (
            O => \N__44328\,
            I => \ppm_encoder_1.un1_init_pulses_10_14\
        );

    \I__9249\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44322\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__44322\,
            I => \N__44318\
        );

    \I__9247\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44315\
        );

    \I__9246\ : Span4Mux_h
    port map (
            O => \N__44318\,
            I => \N__44312\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__44315\,
            I => \N__44309\
        );

    \I__9244\ : Span4Mux_h
    port map (
            O => \N__44312\,
            I => \N__44304\
        );

    \I__9243\ : Span4Mux_h
    port map (
            O => \N__44309\,
            I => \N__44304\
        );

    \I__9242\ : Odrv4
    port map (
            O => \N__44304\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__9241\ : InMux
    port map (
            O => \N__44301\,
            I => \N__44298\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__44298\,
            I => \N__44295\
        );

    \I__9239\ : Span4Mux_v
    port map (
            O => \N__44295\,
            I => \N__44292\
        );

    \I__9238\ : Span4Mux_v
    port map (
            O => \N__44292\,
            I => \N__44289\
        );

    \I__9237\ : Odrv4
    port map (
            O => \N__44289\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\
        );

    \I__9236\ : InMux
    port map (
            O => \N__44286\,
            I => \N__44283\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__44283\,
            I => \ppm_encoder_1.un1_init_pulses_10_2\
        );

    \I__9234\ : InMux
    port map (
            O => \N__44280\,
            I => \N__44277\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__44277\,
            I => \N__44273\
        );

    \I__9232\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44270\
        );

    \I__9231\ : Odrv12
    port map (
            O => \N__44273\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__44270\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__9229\ : InMux
    port map (
            O => \N__44265\,
            I => \N__44262\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__44262\,
            I => \ppm_encoder_1.un1_init_pulses_10_17\
        );

    \I__9227\ : InMux
    port map (
            O => \N__44259\,
            I => \N__44256\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__44256\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_17\
        );

    \I__9225\ : CascadeMux
    port map (
            O => \N__44253\,
            I => \N__44250\
        );

    \I__9224\ : InMux
    port map (
            O => \N__44250\,
            I => \N__44247\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__44247\,
            I => \N__44244\
        );

    \I__9222\ : Odrv4
    port map (
            O => \N__44244\,
            I => \ppm_encoder_1.un1_init_pulses_10_3\
        );

    \I__9221\ : InMux
    port map (
            O => \N__44241\,
            I => \N__44238\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__44238\,
            I => \N__44234\
        );

    \I__9219\ : InMux
    port map (
            O => \N__44237\,
            I => \N__44231\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__44234\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__44231\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__9216\ : InMux
    port map (
            O => \N__44226\,
            I => \N__44220\
        );

    \I__9215\ : InMux
    port map (
            O => \N__44225\,
            I => \N__44220\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__44220\,
            I => \N__44217\
        );

    \I__9213\ : Span4Mux_v
    port map (
            O => \N__44217\,
            I => \N__44213\
        );

    \I__9212\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44210\
        );

    \I__9211\ : Span4Mux_h
    port map (
            O => \N__44213\,
            I => \N__44207\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__44210\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__9209\ : Odrv4
    port map (
            O => \N__44207\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__9208\ : CascadeMux
    port map (
            O => \N__44202\,
            I => \N__44196\
        );

    \I__9207\ : CascadeMux
    port map (
            O => \N__44201\,
            I => \N__44191\
        );

    \I__9206\ : CascadeMux
    port map (
            O => \N__44200\,
            I => \N__44186\
        );

    \I__9205\ : CascadeMux
    port map (
            O => \N__44199\,
            I => \N__44183\
        );

    \I__9204\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44180\
        );

    \I__9203\ : InMux
    port map (
            O => \N__44195\,
            I => \N__44177\
        );

    \I__9202\ : InMux
    port map (
            O => \N__44194\,
            I => \N__44174\
        );

    \I__9201\ : InMux
    port map (
            O => \N__44191\,
            I => \N__44171\
        );

    \I__9200\ : CascadeMux
    port map (
            O => \N__44190\,
            I => \N__44167\
        );

    \I__9199\ : InMux
    port map (
            O => \N__44189\,
            I => \N__44163\
        );

    \I__9198\ : InMux
    port map (
            O => \N__44186\,
            I => \N__44160\
        );

    \I__9197\ : InMux
    port map (
            O => \N__44183\,
            I => \N__44156\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__44180\,
            I => \N__44153\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__44177\,
            I => \N__44148\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__44174\,
            I => \N__44148\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__44171\,
            I => \N__44145\
        );

    \I__9192\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44142\
        );

    \I__9191\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44139\
        );

    \I__9190\ : InMux
    port map (
            O => \N__44166\,
            I => \N__44136\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__44163\,
            I => \N__44133\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__44160\,
            I => \N__44130\
        );

    \I__9187\ : CascadeMux
    port map (
            O => \N__44159\,
            I => \N__44127\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__44156\,
            I => \N__44120\
        );

    \I__9185\ : Span4Mux_v
    port map (
            O => \N__44153\,
            I => \N__44117\
        );

    \I__9184\ : Span4Mux_v
    port map (
            O => \N__44148\,
            I => \N__44108\
        );

    \I__9183\ : Span4Mux_h
    port map (
            O => \N__44145\,
            I => \N__44108\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__44142\,
            I => \N__44108\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__44139\,
            I => \N__44108\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__44136\,
            I => \N__44101\
        );

    \I__9179\ : Span4Mux_h
    port map (
            O => \N__44133\,
            I => \N__44101\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__44130\,
            I => \N__44101\
        );

    \I__9177\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44096\
        );

    \I__9176\ : InMux
    port map (
            O => \N__44126\,
            I => \N__44096\
        );

    \I__9175\ : InMux
    port map (
            O => \N__44125\,
            I => \N__44093\
        );

    \I__9174\ : InMux
    port map (
            O => \N__44124\,
            I => \N__44088\
        );

    \I__9173\ : InMux
    port map (
            O => \N__44123\,
            I => \N__44088\
        );

    \I__9172\ : Odrv4
    port map (
            O => \N__44120\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__9171\ : Odrv4
    port map (
            O => \N__44117\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__9170\ : Odrv4
    port map (
            O => \N__44108\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__44101\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__44096\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__44093\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__44088\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__9165\ : CascadeMux
    port map (
            O => \N__44073\,
            I => \N__44066\
        );

    \I__9164\ : CascadeMux
    port map (
            O => \N__44072\,
            I => \N__44063\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__44071\,
            I => \N__44060\
        );

    \I__9162\ : CascadeMux
    port map (
            O => \N__44070\,
            I => \N__44055\
        );

    \I__9161\ : InMux
    port map (
            O => \N__44069\,
            I => \N__44050\
        );

    \I__9160\ : InMux
    port map (
            O => \N__44066\,
            I => \N__44045\
        );

    \I__9159\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44042\
        );

    \I__9158\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44039\
        );

    \I__9157\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44034\
        );

    \I__9156\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44034\
        );

    \I__9155\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44031\
        );

    \I__9154\ : InMux
    port map (
            O => \N__44054\,
            I => \N__44028\
        );

    \I__9153\ : InMux
    port map (
            O => \N__44053\,
            I => \N__44025\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__44050\,
            I => \N__44022\
        );

    \I__9151\ : InMux
    port map (
            O => \N__44049\,
            I => \N__44015\
        );

    \I__9150\ : InMux
    port map (
            O => \N__44048\,
            I => \N__44015\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__44045\,
            I => \N__44012\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__44042\,
            I => \N__44005\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__44039\,
            I => \N__44005\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__44034\,
            I => \N__44005\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__44031\,
            I => \N__43998\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__44028\,
            I => \N__43998\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__44025\,
            I => \N__43998\
        );

    \I__9142\ : Span4Mux_v
    port map (
            O => \N__44022\,
            I => \N__43995\
        );

    \I__9141\ : InMux
    port map (
            O => \N__44021\,
            I => \N__43992\
        );

    \I__9140\ : InMux
    port map (
            O => \N__44020\,
            I => \N__43989\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__44015\,
            I => \N__43980\
        );

    \I__9138\ : Span4Mux_h
    port map (
            O => \N__44012\,
            I => \N__43980\
        );

    \I__9137\ : Span4Mux_v
    port map (
            O => \N__44005\,
            I => \N__43980\
        );

    \I__9136\ : Span4Mux_v
    port map (
            O => \N__43998\,
            I => \N__43980\
        );

    \I__9135\ : Odrv4
    port map (
            O => \N__43995\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__43992\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__43989\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__9132\ : Odrv4
    port map (
            O => \N__43980\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__9131\ : CascadeMux
    port map (
            O => \N__43971\,
            I => \ppm_encoder_1.un2_throttle_iv_0_3_cascade_\
        );

    \I__9130\ : CascadeMux
    port map (
            O => \N__43968\,
            I => \N__43965\
        );

    \I__9129\ : InMux
    port map (
            O => \N__43965\,
            I => \N__43962\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__43962\,
            I => \ppm_encoder_1.elevator_RNIT3R05Z0Z_3\
        );

    \I__9127\ : InMux
    port map (
            O => \N__43959\,
            I => \N__43956\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__43956\,
            I => \ppm_encoder_1.N_289\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__43953\,
            I => \N__43949\
        );

    \I__9124\ : InMux
    port map (
            O => \N__43952\,
            I => \N__43946\
        );

    \I__9123\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43943\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__43946\,
            I => \N__43940\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__43943\,
            I => \N__43937\
        );

    \I__9120\ : Span4Mux_h
    port map (
            O => \N__43940\,
            I => \N__43934\
        );

    \I__9119\ : Odrv4
    port map (
            O => \N__43937\,
            I => side_order_3
        );

    \I__9118\ : Odrv4
    port map (
            O => \N__43934\,
            I => side_order_3
        );

    \I__9117\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43926\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__43926\,
            I => \N__43923\
        );

    \I__9115\ : Span12Mux_v
    port map (
            O => \N__43923\,
            I => \N__43920\
        );

    \I__9114\ : Odrv12
    port map (
            O => \N__43920\,
            I => \ppm_encoder_1.un1_aileron_cry_2_THRU_CO\
        );

    \I__9113\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43912\
        );

    \I__9112\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43907\
        );

    \I__9111\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43907\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__43912\,
            I => \ppm_encoder_1.aileronZ0Z_3\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__43907\,
            I => \ppm_encoder_1.aileronZ0Z_3\
        );

    \I__9108\ : InMux
    port map (
            O => \N__43902\,
            I => \N__43899\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__43899\,
            I => \N__43896\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__43896\,
            I => \N__43893\
        );

    \I__9105\ : Odrv4
    port map (
            O => \N__43893\,
            I => \ppm_encoder_1.un1_elevator_cry_2_THRU_CO\
        );

    \I__9104\ : InMux
    port map (
            O => \N__43890\,
            I => \N__43887\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__43887\,
            I => \N__43883\
        );

    \I__9102\ : InMux
    port map (
            O => \N__43886\,
            I => \N__43880\
        );

    \I__9101\ : Span4Mux_h
    port map (
            O => \N__43883\,
            I => \N__43875\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__43880\,
            I => \N__43875\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__43875\,
            I => \N__43872\
        );

    \I__9098\ : Span4Mux_v
    port map (
            O => \N__43872\,
            I => \N__43869\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__43869\,
            I => front_order_3
        );

    \I__9096\ : InMux
    port map (
            O => \N__43866\,
            I => \N__43857\
        );

    \I__9095\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43857\
        );

    \I__9094\ : InMux
    port map (
            O => \N__43864\,
            I => \N__43857\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__43857\,
            I => \ppm_encoder_1.elevatorZ0Z_3\
        );

    \I__9092\ : CascadeMux
    port map (
            O => \N__43854\,
            I => \N__43851\
        );

    \I__9091\ : InMux
    port map (
            O => \N__43851\,
            I => \N__43848\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__43848\,
            I => \ppm_encoder_1.un1_init_pulses_10_1\
        );

    \I__9089\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43842\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__43842\,
            I => \N__43838\
        );

    \I__9087\ : InMux
    port map (
            O => \N__43841\,
            I => \N__43835\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__43838\,
            I => \N__43832\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__43835\,
            I => \N__43829\
        );

    \I__9084\ : Odrv4
    port map (
            O => \N__43832\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__9083\ : Odrv4
    port map (
            O => \N__43829\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__9082\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43821\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__43821\,
            I => \N__43818\
        );

    \I__9080\ : Span4Mux_v
    port map (
            O => \N__43818\,
            I => \N__43815\
        );

    \I__9079\ : Span4Mux_v
    port map (
            O => \N__43815\,
            I => \N__43812\
        );

    \I__9078\ : Odrv4
    port map (
            O => \N__43812\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\
        );

    \I__9077\ : CascadeMux
    port map (
            O => \N__43809\,
            I => \N__43806\
        );

    \I__9076\ : InMux
    port map (
            O => \N__43806\,
            I => \N__43803\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__43803\,
            I => \N__43800\
        );

    \I__9074\ : Span4Mux_h
    port map (
            O => \N__43800\,
            I => \N__43797\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__43797\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0\
        );

    \I__9072\ : InMux
    port map (
            O => \N__43794\,
            I => \N__43789\
        );

    \I__9071\ : InMux
    port map (
            O => \N__43793\,
            I => \N__43786\
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__43792\,
            I => \N__43783\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__43789\,
            I => \N__43780\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__43786\,
            I => \N__43777\
        );

    \I__9067\ : InMux
    port map (
            O => \N__43783\,
            I => \N__43774\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__43780\,
            I => \N__43771\
        );

    \I__9065\ : Span4Mux_v
    port map (
            O => \N__43777\,
            I => \N__43768\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__43774\,
            I => \ppm_encoder_1.aileronZ0Z_2\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__43771\,
            I => \ppm_encoder_1.aileronZ0Z_2\
        );

    \I__9062\ : Odrv4
    port map (
            O => \N__43768\,
            I => \ppm_encoder_1.aileronZ0Z_2\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__43761\,
            I => \ppm_encoder_1.un2_throttle_iv_0_2_cascade_\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__43758\,
            I => \N__43755\
        );

    \I__9059\ : InMux
    port map (
            O => \N__43755\,
            I => \N__43752\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__43752\,
            I => \N__43749\
        );

    \I__9057\ : Odrv4
    port map (
            O => \N__43749\,
            I => \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2\
        );

    \I__9056\ : InMux
    port map (
            O => \N__43746\,
            I => \N__43740\
        );

    \I__9055\ : InMux
    port map (
            O => \N__43745\,
            I => \N__43733\
        );

    \I__9054\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43733\
        );

    \I__9053\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43733\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__43740\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__43733\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__9050\ : CascadeMux
    port map (
            O => \N__43728\,
            I => \N__43725\
        );

    \I__9049\ : InMux
    port map (
            O => \N__43725\,
            I => \N__43719\
        );

    \I__9048\ : InMux
    port map (
            O => \N__43724\,
            I => \N__43716\
        );

    \I__9047\ : InMux
    port map (
            O => \N__43723\,
            I => \N__43711\
        );

    \I__9046\ : InMux
    port map (
            O => \N__43722\,
            I => \N__43711\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__43719\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__43716\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__43711\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__43704\,
            I => \N__43700\
        );

    \I__9041\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43696\
        );

    \I__9040\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43693\
        );

    \I__9039\ : InMux
    port map (
            O => \N__43699\,
            I => \N__43688\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__43696\,
            I => \N__43685\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__43693\,
            I => \N__43682\
        );

    \I__9036\ : InMux
    port map (
            O => \N__43692\,
            I => \N__43677\
        );

    \I__9035\ : InMux
    port map (
            O => \N__43691\,
            I => \N__43677\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__43688\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__43685\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9032\ : Odrv4
    port map (
            O => \N__43682\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__43677\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9030\ : InMux
    port map (
            O => \N__43668\,
            I => \N__43664\
        );

    \I__9029\ : InMux
    port map (
            O => \N__43667\,
            I => \N__43661\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__43664\,
            I => \N__43655\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__43661\,
            I => \N__43655\
        );

    \I__9026\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43652\
        );

    \I__9025\ : Span4Mux_v
    port map (
            O => \N__43655\,
            I => \N__43649\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__43652\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__9023\ : Odrv4
    port map (
            O => \N__43649\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__9022\ : CascadeMux
    port map (
            O => \N__43644\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\
        );

    \I__9021\ : CascadeMux
    port map (
            O => \N__43641\,
            I => \ppm_encoder_1.un2_throttle_iv_0_0_cascade_\
        );

    \I__9020\ : InMux
    port map (
            O => \N__43638\,
            I => \N__43635\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__43635\,
            I => \N__43632\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__43632\,
            I => \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0\
        );

    \I__9017\ : InMux
    port map (
            O => \N__43629\,
            I => \N__43625\
        );

    \I__9016\ : InMux
    port map (
            O => \N__43628\,
            I => \N__43622\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__43625\,
            I => \N__43619\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__43622\,
            I => \N__43615\
        );

    \I__9013\ : Span4Mux_h
    port map (
            O => \N__43619\,
            I => \N__43612\
        );

    \I__9012\ : InMux
    port map (
            O => \N__43618\,
            I => \N__43609\
        );

    \I__9011\ : Span4Mux_v
    port map (
            O => \N__43615\,
            I => \N__43605\
        );

    \I__9010\ : Span4Mux_v
    port map (
            O => \N__43612\,
            I => \N__43600\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__43609\,
            I => \N__43600\
        );

    \I__9008\ : InMux
    port map (
            O => \N__43608\,
            I => \N__43597\
        );

    \I__9007\ : Odrv4
    port map (
            O => \N__43605\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__9006\ : Odrv4
    port map (
            O => \N__43600\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__43597\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__9004\ : InMux
    port map (
            O => \N__43590\,
            I => \N__43587\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__43587\,
            I => \N__43583\
        );

    \I__9002\ : InMux
    port map (
            O => \N__43586\,
            I => \N__43580\
        );

    \I__9001\ : Sp12to4
    port map (
            O => \N__43583\,
            I => \N__43575\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__43580\,
            I => \N__43575\
        );

    \I__8999\ : Span12Mux_v
    port map (
            O => \N__43575\,
            I => \N__43570\
        );

    \I__8998\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43565\
        );

    \I__8997\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43565\
        );

    \I__8996\ : Odrv12
    port map (
            O => \N__43570\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__43565\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__8994\ : CascadeMux
    port map (
            O => \N__43560\,
            I => \N__43557\
        );

    \I__8993\ : InMux
    port map (
            O => \N__43557\,
            I => \N__43551\
        );

    \I__8992\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43551\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__43551\,
            I => \N__43548\
        );

    \I__8990\ : Span4Mux_v
    port map (
            O => \N__43548\,
            I => \N__43545\
        );

    \I__8989\ : Span4Mux_v
    port map (
            O => \N__43545\,
            I => \N__43542\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__43542\,
            I => \ppm_encoder_1.N_232\
        );

    \I__8987\ : CascadeMux
    port map (
            O => \N__43539\,
            I => \N__43533\
        );

    \I__8986\ : InMux
    port map (
            O => \N__43538\,
            I => \N__43530\
        );

    \I__8985\ : InMux
    port map (
            O => \N__43537\,
            I => \N__43527\
        );

    \I__8984\ : InMux
    port map (
            O => \N__43536\,
            I => \N__43524\
        );

    \I__8983\ : InMux
    port map (
            O => \N__43533\,
            I => \N__43521\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__43530\,
            I => \N__43518\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__43527\,
            I => \N__43512\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__43524\,
            I => \N__43512\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__43521\,
            I => \N__43505\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__43518\,
            I => \N__43505\
        );

    \I__8977\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43502\
        );

    \I__8976\ : Sp12to4
    port map (
            O => \N__43512\,
            I => \N__43499\
        );

    \I__8975\ : InMux
    port map (
            O => \N__43511\,
            I => \N__43494\
        );

    \I__8974\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43494\
        );

    \I__8973\ : Odrv4
    port map (
            O => \N__43505\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__43502\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__8971\ : Odrv12
    port map (
            O => \N__43499\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__43494\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__8969\ : InMux
    port map (
            O => \N__43485\,
            I => \N__43476\
        );

    \I__8968\ : InMux
    port map (
            O => \N__43484\,
            I => \N__43473\
        );

    \I__8967\ : InMux
    port map (
            O => \N__43483\,
            I => \N__43468\
        );

    \I__8966\ : InMux
    port map (
            O => \N__43482\,
            I => \N__43468\
        );

    \I__8965\ : InMux
    port map (
            O => \N__43481\,
            I => \N__43463\
        );

    \I__8964\ : InMux
    port map (
            O => \N__43480\,
            I => \N__43463\
        );

    \I__8963\ : InMux
    port map (
            O => \N__43479\,
            I => \N__43460\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__43476\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__43473\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__43468\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__43463\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__43460\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__43449\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_\
        );

    \I__8956\ : CascadeMux
    port map (
            O => \N__43446\,
            I => \N__43442\
        );

    \I__8955\ : CascadeMux
    port map (
            O => \N__43445\,
            I => \N__43439\
        );

    \I__8954\ : InMux
    port map (
            O => \N__43442\,
            I => \N__43432\
        );

    \I__8953\ : InMux
    port map (
            O => \N__43439\,
            I => \N__43429\
        );

    \I__8952\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43424\
        );

    \I__8951\ : InMux
    port map (
            O => \N__43437\,
            I => \N__43424\
        );

    \I__8950\ : InMux
    port map (
            O => \N__43436\,
            I => \N__43419\
        );

    \I__8949\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43419\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__43432\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__43429\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__43424\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__43419\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__43410\,
            I => \N__43405\
        );

    \I__8943\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43402\
        );

    \I__8942\ : InMux
    port map (
            O => \N__43408\,
            I => \N__43399\
        );

    \I__8941\ : InMux
    port map (
            O => \N__43405\,
            I => \N__43396\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__43402\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__43399\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__43396\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__8937\ : InMux
    port map (
            O => \N__43389\,
            I => \N__43384\
        );

    \I__8936\ : InMux
    port map (
            O => \N__43388\,
            I => \N__43379\
        );

    \I__8935\ : InMux
    port map (
            O => \N__43387\,
            I => \N__43376\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43373\
        );

    \I__8933\ : InMux
    port map (
            O => \N__43383\,
            I => \N__43368\
        );

    \I__8932\ : InMux
    port map (
            O => \N__43382\,
            I => \N__43368\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__43379\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__43376\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8929\ : Odrv4
    port map (
            O => \N__43373\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__43368\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__43359\,
            I => \N__43352\
        );

    \I__8926\ : InMux
    port map (
            O => \N__43358\,
            I => \N__43347\
        );

    \I__8925\ : InMux
    port map (
            O => \N__43357\,
            I => \N__43344\
        );

    \I__8924\ : InMux
    port map (
            O => \N__43356\,
            I => \N__43337\
        );

    \I__8923\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43337\
        );

    \I__8922\ : InMux
    port map (
            O => \N__43352\,
            I => \N__43337\
        );

    \I__8921\ : InMux
    port map (
            O => \N__43351\,
            I => \N__43332\
        );

    \I__8920\ : InMux
    port map (
            O => \N__43350\,
            I => \N__43332\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__43347\,
            I => \N__43327\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__43344\,
            I => \N__43327\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__43337\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__43332\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__8915\ : Odrv4
    port map (
            O => \N__43327\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__8914\ : CascadeMux
    port map (
            O => \N__43320\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\
        );

    \I__8913\ : CascadeMux
    port map (
            O => \N__43317\,
            I => \N__43313\
        );

    \I__8912\ : InMux
    port map (
            O => \N__43316\,
            I => \N__43309\
        );

    \I__8911\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43306\
        );

    \I__8910\ : InMux
    port map (
            O => \N__43312\,
            I => \N__43303\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__43309\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_6\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__43306\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_6\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__43303\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_6\
        );

    \I__8906\ : CascadeMux
    port map (
            O => \N__43296\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_\
        );

    \I__8905\ : InMux
    port map (
            O => \N__43293\,
            I => \N__43290\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__43290\,
            I => \N__43286\
        );

    \I__8903\ : InMux
    port map (
            O => \N__43289\,
            I => \N__43283\
        );

    \I__8902\ : Span12Mux_h
    port map (
            O => \N__43286\,
            I => \N__43280\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__43283\,
            I => side_order_0
        );

    \I__8900\ : Odrv12
    port map (
            O => \N__43280\,
            I => side_order_0
        );

    \I__8899\ : InMux
    port map (
            O => \N__43275\,
            I => \N__43271\
        );

    \I__8898\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43268\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43265\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__43268\,
            I => \N__43262\
        );

    \I__8895\ : Span4Mux_v
    port map (
            O => \N__43265\,
            I => \N__43259\
        );

    \I__8894\ : Span4Mux_v
    port map (
            O => \N__43262\,
            I => \N__43256\
        );

    \I__8893\ : Span4Mux_h
    port map (
            O => \N__43259\,
            I => \N__43253\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__43256\,
            I => side_order_5
        );

    \I__8891\ : Odrv4
    port map (
            O => \N__43253\,
            I => side_order_5
        );

    \I__8890\ : InMux
    port map (
            O => \N__43248\,
            I => \N__43244\
        );

    \I__8889\ : InMux
    port map (
            O => \N__43247\,
            I => \N__43241\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__43244\,
            I => \N__43236\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__43241\,
            I => \N__43236\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__43236\,
            I => \N__43233\
        );

    \I__8885\ : Span4Mux_h
    port map (
            O => \N__43233\,
            I => \N__43230\
        );

    \I__8884\ : Odrv4
    port map (
            O => \N__43230\,
            I => side_order_4
        );

    \I__8883\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43224\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__43224\,
            I => \N__43220\
        );

    \I__8881\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43217\
        );

    \I__8880\ : Span4Mux_v
    port map (
            O => \N__43220\,
            I => \N__43211\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__43217\,
            I => \N__43211\
        );

    \I__8878\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43208\
        );

    \I__8877\ : Span4Mux_h
    port map (
            O => \N__43211\,
            I => \N__43205\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__43208\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__43205\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__8874\ : InMux
    port map (
            O => \N__43200\,
            I => \N__43196\
        );

    \I__8873\ : CascadeMux
    port map (
            O => \N__43199\,
            I => \N__43193\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__43196\,
            I => \N__43190\
        );

    \I__8871\ : InMux
    port map (
            O => \N__43193\,
            I => \N__43186\
        );

    \I__8870\ : Span4Mux_v
    port map (
            O => \N__43190\,
            I => \N__43183\
        );

    \I__8869\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43180\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__43186\,
            I => \N__43173\
        );

    \I__8867\ : Span4Mux_h
    port map (
            O => \N__43183\,
            I => \N__43173\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43173\
        );

    \I__8865\ : Odrv4
    port map (
            O => \N__43173\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__8864\ : CascadeMux
    port map (
            O => \N__43170\,
            I => \N__43167\
        );

    \I__8863\ : InMux
    port map (
            O => \N__43167\,
            I => \N__43164\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__43164\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__8861\ : CascadeMux
    port map (
            O => \N__43161\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\
        );

    \I__8860\ : InMux
    port map (
            O => \N__43158\,
            I => \N__43153\
        );

    \I__8859\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43148\
        );

    \I__8858\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43148\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__43153\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__43148\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__8855\ : InMux
    port map (
            O => \N__43143\,
            I => \N__43138\
        );

    \I__8854\ : InMux
    port map (
            O => \N__43142\,
            I => \N__43133\
        );

    \I__8853\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43133\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__43138\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__43133\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__8850\ : CascadeMux
    port map (
            O => \N__43128\,
            I => \N__43125\
        );

    \I__8849\ : InMux
    port map (
            O => \N__43125\,
            I => \N__43121\
        );

    \I__8848\ : InMux
    port map (
            O => \N__43124\,
            I => \N__43117\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__43121\,
            I => \N__43114\
        );

    \I__8846\ : InMux
    port map (
            O => \N__43120\,
            I => \N__43111\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__43117\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__8844\ : Odrv4
    port map (
            O => \N__43114\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__43111\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__8842\ : InMux
    port map (
            O => \N__43104\,
            I => \N__43099\
        );

    \I__8841\ : InMux
    port map (
            O => \N__43103\,
            I => \N__43096\
        );

    \I__8840\ : InMux
    port map (
            O => \N__43102\,
            I => \N__43093\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__43099\,
            I => \N__43090\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__43096\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__43093\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__8836\ : Odrv4
    port map (
            O => \N__43090\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__8835\ : CascadeMux
    port map (
            O => \N__43083\,
            I => \N__43079\
        );

    \I__8834\ : InMux
    port map (
            O => \N__43082\,
            I => \N__43074\
        );

    \I__8833\ : InMux
    port map (
            O => \N__43079\,
            I => \N__43074\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__43074\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\
        );

    \I__8831\ : InMux
    port map (
            O => \N__43071\,
            I => \N__43068\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__43068\,
            I => \N__43065\
        );

    \I__8829\ : Span4Mux_v
    port map (
            O => \N__43065\,
            I => \N__43062\
        );

    \I__8828\ : Odrv4
    port map (
            O => \N__43062\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_16\
        );

    \I__8827\ : CascadeMux
    port map (
            O => \N__43059\,
            I => \N__43056\
        );

    \I__8826\ : InMux
    port map (
            O => \N__43056\,
            I => \N__43050\
        );

    \I__8825\ : InMux
    port map (
            O => \N__43055\,
            I => \N__43050\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__43050\,
            I => \N__43047\
        );

    \I__8823\ : Odrv4
    port map (
            O => \N__43047\,
            I => \pid_front.error_d_reg_prevZ0Z_20\
        );

    \I__8822\ : InMux
    port map (
            O => \N__43044\,
            I => \N__43040\
        );

    \I__8821\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43037\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__43040\,
            I => \N__43034\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__43037\,
            I => \N__43028\
        );

    \I__8818\ : Span4Mux_v
    port map (
            O => \N__43034\,
            I => \N__43028\
        );

    \I__8817\ : CascadeMux
    port map (
            O => \N__43033\,
            I => \N__43025\
        );

    \I__8816\ : Span4Mux_v
    port map (
            O => \N__43028\,
            I => \N__43022\
        );

    \I__8815\ : InMux
    port map (
            O => \N__43025\,
            I => \N__43019\
        );

    \I__8814\ : Span4Mux_h
    port map (
            O => \N__43022\,
            I => \N__43016\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__43019\,
            I => side_order_10
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__43016\,
            I => side_order_10
        );

    \I__8811\ : InMux
    port map (
            O => \N__43011\,
            I => \N__43007\
        );

    \I__8810\ : CascadeMux
    port map (
            O => \N__43010\,
            I => \N__43003\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__43007\,
            I => \N__43000\
        );

    \I__8808\ : CascadeMux
    port map (
            O => \N__43006\,
            I => \N__42997\
        );

    \I__8807\ : InMux
    port map (
            O => \N__43003\,
            I => \N__42994\
        );

    \I__8806\ : Span4Mux_v
    port map (
            O => \N__43000\,
            I => \N__42991\
        );

    \I__8805\ : InMux
    port map (
            O => \N__42997\,
            I => \N__42988\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__42994\,
            I => \N__42983\
        );

    \I__8803\ : Span4Mux_h
    port map (
            O => \N__42991\,
            I => \N__42983\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__42988\,
            I => \N__42978\
        );

    \I__8801\ : Span4Mux_v
    port map (
            O => \N__42983\,
            I => \N__42978\
        );

    \I__8800\ : Odrv4
    port map (
            O => \N__42978\,
            I => side_order_11
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__42975\,
            I => \N__42971\
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__42974\,
            I => \N__42968\
        );

    \I__8797\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42965\
        );

    \I__8796\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42962\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__42965\,
            I => \N__42958\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__42962\,
            I => \N__42955\
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__42961\,
            I => \N__42952\
        );

    \I__8792\ : Span4Mux_v
    port map (
            O => \N__42958\,
            I => \N__42949\
        );

    \I__8791\ : Span4Mux_v
    port map (
            O => \N__42955\,
            I => \N__42946\
        );

    \I__8790\ : InMux
    port map (
            O => \N__42952\,
            I => \N__42943\
        );

    \I__8789\ : Span4Mux_v
    port map (
            O => \N__42949\,
            I => \N__42940\
        );

    \I__8788\ : Span4Mux_h
    port map (
            O => \N__42946\,
            I => \N__42937\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__42943\,
            I => side_order_6
        );

    \I__8786\ : Odrv4
    port map (
            O => \N__42940\,
            I => side_order_6
        );

    \I__8785\ : Odrv4
    port map (
            O => \N__42937\,
            I => side_order_6
        );

    \I__8784\ : CascadeMux
    port map (
            O => \N__42930\,
            I => \N__42926\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__42929\,
            I => \N__42923\
        );

    \I__8782\ : InMux
    port map (
            O => \N__42926\,
            I => \N__42920\
        );

    \I__8781\ : InMux
    port map (
            O => \N__42923\,
            I => \N__42917\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__42920\,
            I => \N__42913\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__42917\,
            I => \N__42910\
        );

    \I__8778\ : CascadeMux
    port map (
            O => \N__42916\,
            I => \N__42907\
        );

    \I__8777\ : Span4Mux_h
    port map (
            O => \N__42913\,
            I => \N__42904\
        );

    \I__8776\ : Span4Mux_v
    port map (
            O => \N__42910\,
            I => \N__42901\
        );

    \I__8775\ : InMux
    port map (
            O => \N__42907\,
            I => \N__42898\
        );

    \I__8774\ : Sp12to4
    port map (
            O => \N__42904\,
            I => \N__42895\
        );

    \I__8773\ : Span4Mux_h
    port map (
            O => \N__42901\,
            I => \N__42892\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__42898\,
            I => side_order_7
        );

    \I__8771\ : Odrv12
    port map (
            O => \N__42895\,
            I => side_order_7
        );

    \I__8770\ : Odrv4
    port map (
            O => \N__42892\,
            I => side_order_7
        );

    \I__8769\ : InMux
    port map (
            O => \N__42885\,
            I => \N__42881\
        );

    \I__8768\ : InMux
    port map (
            O => \N__42884\,
            I => \N__42878\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__42881\,
            I => \N__42875\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__42878\,
            I => \N__42872\
        );

    \I__8765\ : Span4Mux_v
    port map (
            O => \N__42875\,
            I => \N__42866\
        );

    \I__8764\ : Span4Mux_v
    port map (
            O => \N__42872\,
            I => \N__42866\
        );

    \I__8763\ : CascadeMux
    port map (
            O => \N__42871\,
            I => \N__42863\
        );

    \I__8762\ : Span4Mux_h
    port map (
            O => \N__42866\,
            I => \N__42860\
        );

    \I__8761\ : InMux
    port map (
            O => \N__42863\,
            I => \N__42857\
        );

    \I__8760\ : Span4Mux_v
    port map (
            O => \N__42860\,
            I => \N__42854\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__42857\,
            I => side_order_8
        );

    \I__8758\ : Odrv4
    port map (
            O => \N__42854\,
            I => side_order_8
        );

    \I__8757\ : InMux
    port map (
            O => \N__42849\,
            I => \N__42845\
        );

    \I__8756\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42842\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__42845\,
            I => \N__42839\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__42842\,
            I => \N__42836\
        );

    \I__8753\ : Span4Mux_v
    port map (
            O => \N__42839\,
            I => \N__42832\
        );

    \I__8752\ : Span4Mux_h
    port map (
            O => \N__42836\,
            I => \N__42829\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__42835\,
            I => \N__42826\
        );

    \I__8750\ : Span4Mux_h
    port map (
            O => \N__42832\,
            I => \N__42821\
        );

    \I__8749\ : Span4Mux_v
    port map (
            O => \N__42829\,
            I => \N__42821\
        );

    \I__8748\ : InMux
    port map (
            O => \N__42826\,
            I => \N__42818\
        );

    \I__8747\ : Span4Mux_v
    port map (
            O => \N__42821\,
            I => \N__42815\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__42818\,
            I => side_order_9
        );

    \I__8745\ : Odrv4
    port map (
            O => \N__42815\,
            I => side_order_9
        );

    \I__8744\ : InMux
    port map (
            O => \N__42810\,
            I => \N__42805\
        );

    \I__8743\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42802\
        );

    \I__8742\ : InMux
    port map (
            O => \N__42808\,
            I => \N__42799\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__42805\,
            I => \N__42796\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__42802\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__42799\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__8738\ : Odrv4
    port map (
            O => \N__42796\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__8737\ : InMux
    port map (
            O => \N__42789\,
            I => \N__42784\
        );

    \I__8736\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42781\
        );

    \I__8735\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42778\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__42784\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__42781\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__42778\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__8731\ : CascadeMux
    port map (
            O => \N__42771\,
            I => \N__42766\
        );

    \I__8730\ : InMux
    port map (
            O => \N__42770\,
            I => \N__42763\
        );

    \I__8729\ : InMux
    port map (
            O => \N__42769\,
            I => \N__42760\
        );

    \I__8728\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42757\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__42763\,
            I => \N__42754\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__42760\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__42757\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__42754\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__8723\ : CascadeMux
    port map (
            O => \N__42747\,
            I => \N__42742\
        );

    \I__8722\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42739\
        );

    \I__8721\ : InMux
    port map (
            O => \N__42745\,
            I => \N__42736\
        );

    \I__8720\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42733\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__42739\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__42736\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__42733\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__8716\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42723\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__42723\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\
        );

    \I__8714\ : InMux
    port map (
            O => \N__42720\,
            I => \N__42715\
        );

    \I__8713\ : InMux
    port map (
            O => \N__42719\,
            I => \N__42712\
        );

    \I__8712\ : InMux
    port map (
            O => \N__42718\,
            I => \N__42709\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__42715\,
            I => \N__42706\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__42712\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__42709\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__8708\ : Odrv4
    port map (
            O => \N__42706\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__8707\ : CascadeMux
    port map (
            O => \N__42699\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\
        );

    \I__8706\ : CascadeMux
    port map (
            O => \N__42696\,
            I => \N__42693\
        );

    \I__8705\ : InMux
    port map (
            O => \N__42693\,
            I => \N__42688\
        );

    \I__8704\ : InMux
    port map (
            O => \N__42692\,
            I => \N__42685\
        );

    \I__8703\ : InMux
    port map (
            O => \N__42691\,
            I => \N__42682\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__42688\,
            I => \N__42679\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__42685\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__42682\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__8699\ : Odrv4
    port map (
            O => \N__42679\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__8698\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42669\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__42669\,
            I => \ppm_encoder_1.N_139_17\
        );

    \I__8696\ : InMux
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__42663\,
            I => \N__42660\
        );

    \I__8694\ : Odrv4
    port map (
            O => \N__42660\,
            I => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\
        );

    \I__8693\ : CascadeMux
    port map (
            O => \N__42657\,
            I => \ppm_encoder_1.N_139_17_cascade_\
        );

    \I__8692\ : InMux
    port map (
            O => \N__42654\,
            I => \N__42651\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__42651\,
            I => \N__42648\
        );

    \I__8690\ : Span4Mux_h
    port map (
            O => \N__42648\,
            I => \N__42645\
        );

    \I__8689\ : Span4Mux_v
    port map (
            O => \N__42645\,
            I => \N__42642\
        );

    \I__8688\ : Span4Mux_v
    port map (
            O => \N__42642\,
            I => \N__42639\
        );

    \I__8687\ : Odrv4
    port map (
            O => \N__42639\,
            I => \ppm_encoder_1.N_139\
        );

    \I__8686\ : CascadeMux
    port map (
            O => \N__42636\,
            I => \N__42629\
        );

    \I__8685\ : InMux
    port map (
            O => \N__42635\,
            I => \N__42622\
        );

    \I__8684\ : InMux
    port map (
            O => \N__42634\,
            I => \N__42622\
        );

    \I__8683\ : InMux
    port map (
            O => \N__42633\,
            I => \N__42617\
        );

    \I__8682\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42617\
        );

    \I__8681\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42614\
        );

    \I__8680\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42611\
        );

    \I__8679\ : InMux
    port map (
            O => \N__42627\,
            I => \N__42606\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__42622\,
            I => \N__42603\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__42617\,
            I => \N__42598\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__42614\,
            I => \N__42598\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__42611\,
            I => \N__42595\
        );

    \I__8674\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42590\
        );

    \I__8673\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42590\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__42606\,
            I => \N__42587\
        );

    \I__8671\ : Span4Mux_h
    port map (
            O => \N__42603\,
            I => \N__42582\
        );

    \I__8670\ : Span4Mux_h
    port map (
            O => \N__42598\,
            I => \N__42582\
        );

    \I__8669\ : Span4Mux_h
    port map (
            O => \N__42595\,
            I => \N__42579\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__42590\,
            I => \N__42572\
        );

    \I__8667\ : Span4Mux_v
    port map (
            O => \N__42587\,
            I => \N__42572\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__42582\,
            I => \N__42572\
        );

    \I__8665\ : Odrv4
    port map (
            O => \N__42579\,
            I => \pid_front.un1_pid_prereg_92\
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__42572\,
            I => \pid_front.un1_pid_prereg_92\
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__42567\,
            I => \N__42563\
        );

    \I__8662\ : InMux
    port map (
            O => \N__42566\,
            I => \N__42556\
        );

    \I__8661\ : InMux
    port map (
            O => \N__42563\,
            I => \N__42556\
        );

    \I__8660\ : InMux
    port map (
            O => \N__42562\,
            I => \N__42553\
        );

    \I__8659\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42549\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__42556\,
            I => \N__42546\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__42553\,
            I => \N__42543\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__42552\,
            I => \N__42540\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__42549\,
            I => \N__42536\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__42546\,
            I => \N__42531\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__42543\,
            I => \N__42531\
        );

    \I__8652\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42526\
        );

    \I__8651\ : InMux
    port map (
            O => \N__42539\,
            I => \N__42526\
        );

    \I__8650\ : Span4Mux_v
    port map (
            O => \N__42536\,
            I => \N__42521\
        );

    \I__8649\ : Span4Mux_v
    port map (
            O => \N__42531\,
            I => \N__42521\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__42526\,
            I => \pid_front.un1_pid_prereg_93\
        );

    \I__8647\ : Odrv4
    port map (
            O => \N__42521\,
            I => \pid_front.un1_pid_prereg_93\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__42516\,
            I => \N__42513\
        );

    \I__8645\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42510\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__42510\,
            I => \N__42507\
        );

    \I__8643\ : Odrv4
    port map (
            O => \N__42507\,
            I => \pid_front.error_p_reg_esr_RNIGKTC2Z0Z_20\
        );

    \I__8642\ : InMux
    port map (
            O => \N__42504\,
            I => \N__42501\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__42501\,
            I => \N__42498\
        );

    \I__8640\ : Odrv4
    port map (
            O => \N__42498\,
            I => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__42495\,
            I => \N__42492\
        );

    \I__8638\ : InMux
    port map (
            O => \N__42492\,
            I => \N__42488\
        );

    \I__8637\ : InMux
    port map (
            O => \N__42491\,
            I => \N__42485\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__42488\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__42485\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__8634\ : CascadeMux
    port map (
            O => \N__42480\,
            I => \N__42477\
        );

    \I__8633\ : InMux
    port map (
            O => \N__42477\,
            I => \N__42471\
        );

    \I__8632\ : InMux
    port map (
            O => \N__42476\,
            I => \N__42471\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__42471\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__8630\ : InMux
    port map (
            O => \N__42468\,
            I => \N__42465\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__42465\,
            I => \N__42462\
        );

    \I__8628\ : Odrv4
    port map (
            O => \N__42462\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\
        );

    \I__8627\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42454\
        );

    \I__8626\ : InMux
    port map (
            O => \N__42458\,
            I => \N__42451\
        );

    \I__8625\ : IoInMux
    port map (
            O => \N__42457\,
            I => \N__42443\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__42454\,
            I => \N__42436\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__42451\,
            I => \N__42433\
        );

    \I__8622\ : CascadeMux
    port map (
            O => \N__42450\,
            I => \N__42429\
        );

    \I__8621\ : CascadeMux
    port map (
            O => \N__42449\,
            I => \N__42426\
        );

    \I__8620\ : CascadeMux
    port map (
            O => \N__42448\,
            I => \N__42423\
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__42447\,
            I => \N__42420\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__42446\,
            I => \N__42417\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__42443\,
            I => \N__42414\
        );

    \I__8616\ : CascadeMux
    port map (
            O => \N__42442\,
            I => \N__42411\
        );

    \I__8615\ : CascadeMux
    port map (
            O => \N__42441\,
            I => \N__42408\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__42440\,
            I => \N__42405\
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__42439\,
            I => \N__42402\
        );

    \I__8612\ : Span4Mux_v
    port map (
            O => \N__42436\,
            I => \N__42399\
        );

    \I__8611\ : Span4Mux_v
    port map (
            O => \N__42433\,
            I => \N__42396\
        );

    \I__8610\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42393\
        );

    \I__8609\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42389\
        );

    \I__8608\ : InMux
    port map (
            O => \N__42426\,
            I => \N__42380\
        );

    \I__8607\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42380\
        );

    \I__8606\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42380\
        );

    \I__8605\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42380\
        );

    \I__8604\ : Span4Mux_s2_v
    port map (
            O => \N__42414\,
            I => \N__42377\
        );

    \I__8603\ : InMux
    port map (
            O => \N__42411\,
            I => \N__42374\
        );

    \I__8602\ : InMux
    port map (
            O => \N__42408\,
            I => \N__42367\
        );

    \I__8601\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42367\
        );

    \I__8600\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42367\
        );

    \I__8599\ : Span4Mux_v
    port map (
            O => \N__42399\,
            I => \N__42356\
        );

    \I__8598\ : Span4Mux_v
    port map (
            O => \N__42396\,
            I => \N__42356\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__42393\,
            I => \N__42356\
        );

    \I__8596\ : InMux
    port map (
            O => \N__42392\,
            I => \N__42353\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__42389\,
            I => \N__42347\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__42380\,
            I => \N__42347\
        );

    \I__8593\ : Span4Mux_v
    port map (
            O => \N__42377\,
            I => \N__42340\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__42374\,
            I => \N__42340\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__42367\,
            I => \N__42340\
        );

    \I__8590\ : CascadeMux
    port map (
            O => \N__42366\,
            I => \N__42337\
        );

    \I__8589\ : CascadeMux
    port map (
            O => \N__42365\,
            I => \N__42333\
        );

    \I__8588\ : CascadeMux
    port map (
            O => \N__42364\,
            I => \N__42330\
        );

    \I__8587\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42327\
        );

    \I__8586\ : Span4Mux_v
    port map (
            O => \N__42356\,
            I => \N__42321\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__42353\,
            I => \N__42321\
        );

    \I__8584\ : CascadeMux
    port map (
            O => \N__42352\,
            I => \N__42318\
        );

    \I__8583\ : Span4Mux_v
    port map (
            O => \N__42347\,
            I => \N__42310\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__42340\,
            I => \N__42310\
        );

    \I__8581\ : InMux
    port map (
            O => \N__42337\,
            I => \N__42307\
        );

    \I__8580\ : InMux
    port map (
            O => \N__42336\,
            I => \N__42300\
        );

    \I__8579\ : InMux
    port map (
            O => \N__42333\,
            I => \N__42300\
        );

    \I__8578\ : InMux
    port map (
            O => \N__42330\,
            I => \N__42300\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__42327\,
            I => \N__42292\
        );

    \I__8576\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42289\
        );

    \I__8575\ : Span4Mux_v
    port map (
            O => \N__42321\,
            I => \N__42282\
        );

    \I__8574\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42279\
        );

    \I__8573\ : CascadeMux
    port map (
            O => \N__42317\,
            I => \N__42275\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__42316\,
            I => \N__42272\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__42315\,
            I => \N__42269\
        );

    \I__8570\ : Span4Mux_h
    port map (
            O => \N__42310\,
            I => \N__42262\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__42307\,
            I => \N__42262\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__42300\,
            I => \N__42262\
        );

    \I__8567\ : InMux
    port map (
            O => \N__42299\,
            I => \N__42259\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__42298\,
            I => \N__42255\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__42297\,
            I => \N__42252\
        );

    \I__8564\ : CascadeMux
    port map (
            O => \N__42296\,
            I => \N__42249\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__42295\,
            I => \N__42246\
        );

    \I__8562\ : Span4Mux_v
    port map (
            O => \N__42292\,
            I => \N__42241\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__42289\,
            I => \N__42241\
        );

    \I__8560\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42238\
        );

    \I__8559\ : InMux
    port map (
            O => \N__42287\,
            I => \N__42234\
        );

    \I__8558\ : InMux
    port map (
            O => \N__42286\,
            I => \N__42231\
        );

    \I__8557\ : InMux
    port map (
            O => \N__42285\,
            I => \N__42225\
        );

    \I__8556\ : Span4Mux_h
    port map (
            O => \N__42282\,
            I => \N__42222\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__42279\,
            I => \N__42219\
        );

    \I__8554\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42212\
        );

    \I__8553\ : InMux
    port map (
            O => \N__42275\,
            I => \N__42212\
        );

    \I__8552\ : InMux
    port map (
            O => \N__42272\,
            I => \N__42212\
        );

    \I__8551\ : InMux
    port map (
            O => \N__42269\,
            I => \N__42209\
        );

    \I__8550\ : Span4Mux_v
    port map (
            O => \N__42262\,
            I => \N__42206\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__42259\,
            I => \N__42203\
        );

    \I__8548\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42200\
        );

    \I__8547\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42197\
        );

    \I__8546\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42194\
        );

    \I__8545\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42189\
        );

    \I__8544\ : InMux
    port map (
            O => \N__42246\,
            I => \N__42189\
        );

    \I__8543\ : Span4Mux_v
    port map (
            O => \N__42241\,
            I => \N__42184\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__42238\,
            I => \N__42184\
        );

    \I__8541\ : InMux
    port map (
            O => \N__42237\,
            I => \N__42181\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__42234\,
            I => \N__42176\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__42231\,
            I => \N__42176\
        );

    \I__8538\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42173\
        );

    \I__8537\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42170\
        );

    \I__8536\ : InMux
    port map (
            O => \N__42228\,
            I => \N__42167\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__42225\,
            I => \N__42164\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__42222\,
            I => \N__42161\
        );

    \I__8533\ : Span4Mux_v
    port map (
            O => \N__42219\,
            I => \N__42156\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__42212\,
            I => \N__42156\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42153\
        );

    \I__8530\ : Span4Mux_h
    port map (
            O => \N__42206\,
            I => \N__42148\
        );

    \I__8529\ : Span4Mux_v
    port map (
            O => \N__42203\,
            I => \N__42148\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__42200\,
            I => \N__42139\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__42197\,
            I => \N__42139\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__42194\,
            I => \N__42139\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__42189\,
            I => \N__42139\
        );

    \I__8524\ : Span4Mux_v
    port map (
            O => \N__42184\,
            I => \N__42134\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__42181\,
            I => \N__42134\
        );

    \I__8522\ : Span4Mux_v
    port map (
            O => \N__42176\,
            I => \N__42127\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__42173\,
            I => \N__42127\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__42170\,
            I => \N__42127\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__42167\,
            I => \N__42124\
        );

    \I__8518\ : Span12Mux_s8_h
    port map (
            O => \N__42164\,
            I => \N__42119\
        );

    \I__8517\ : Sp12to4
    port map (
            O => \N__42161\,
            I => \N__42119\
        );

    \I__8516\ : Span4Mux_v
    port map (
            O => \N__42156\,
            I => \N__42114\
        );

    \I__8515\ : Span4Mux_v
    port map (
            O => \N__42153\,
            I => \N__42114\
        );

    \I__8514\ : Span4Mux_v
    port map (
            O => \N__42148\,
            I => \N__42109\
        );

    \I__8513\ : Span4Mux_v
    port map (
            O => \N__42139\,
            I => \N__42109\
        );

    \I__8512\ : Span4Mux_v
    port map (
            O => \N__42134\,
            I => \N__42104\
        );

    \I__8511\ : Span4Mux_v
    port map (
            O => \N__42127\,
            I => \N__42104\
        );

    \I__8510\ : Span12Mux_s8_h
    port map (
            O => \N__42124\,
            I => \N__42095\
        );

    \I__8509\ : Span12Mux_v
    port map (
            O => \N__42119\,
            I => \N__42095\
        );

    \I__8508\ : Sp12to4
    port map (
            O => \N__42114\,
            I => \N__42095\
        );

    \I__8507\ : Sp12to4
    port map (
            O => \N__42109\,
            I => \N__42095\
        );

    \I__8506\ : Span4Mux_h
    port map (
            O => \N__42104\,
            I => \N__42092\
        );

    \I__8505\ : Odrv12
    port map (
            O => \N__42095\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8504\ : Odrv4
    port map (
            O => \N__42092\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8503\ : InMux
    port map (
            O => \N__42087\,
            I => \ppm_encoder_1.counter24_0_N_2\
        );

    \I__8502\ : InMux
    port map (
            O => \N__42084\,
            I => \N__42081\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__42081\,
            I => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\
        );

    \I__8500\ : InMux
    port map (
            O => \N__42078\,
            I => \N__42072\
        );

    \I__8499\ : InMux
    port map (
            O => \N__42077\,
            I => \N__42069\
        );

    \I__8498\ : InMux
    port map (
            O => \N__42076\,
            I => \N__42064\
        );

    \I__8497\ : InMux
    port map (
            O => \N__42075\,
            I => \N__42064\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__42072\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__42069\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__42064\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__42057\,
            I => \N__42053\
        );

    \I__8492\ : InMux
    port map (
            O => \N__42056\,
            I => \N__42048\
        );

    \I__8491\ : InMux
    port map (
            O => \N__42053\,
            I => \N__42045\
        );

    \I__8490\ : InMux
    port map (
            O => \N__42052\,
            I => \N__42040\
        );

    \I__8489\ : InMux
    port map (
            O => \N__42051\,
            I => \N__42040\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__42048\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__42045\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__42040\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__8485\ : InMux
    port map (
            O => \N__42033\,
            I => \N__42030\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__42030\,
            I => \ppm_encoder_1.pulses2countZ0Z_2\
        );

    \I__8483\ : CascadeMux
    port map (
            O => \N__42027\,
            I => \N__42022\
        );

    \I__8482\ : InMux
    port map (
            O => \N__42026\,
            I => \N__42018\
        );

    \I__8481\ : InMux
    port map (
            O => \N__42025\,
            I => \N__42015\
        );

    \I__8480\ : InMux
    port map (
            O => \N__42022\,
            I => \N__42010\
        );

    \I__8479\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42010\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__42018\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__42015\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__42010\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__8475\ : InMux
    port map (
            O => \N__42003\,
            I => \N__42000\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__42000\,
            I => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\
        );

    \I__8473\ : InMux
    port map (
            O => \N__41997\,
            I => \N__41994\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__41994\,
            I => \N__41991\
        );

    \I__8471\ : Odrv4
    port map (
            O => \N__41991\,
            I => \ppm_encoder_1.pulses2countZ0Z_4\
        );

    \I__8470\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41985\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__41985\,
            I => \N__41982\
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__41982\,
            I => \ppm_encoder_1.pulses2countZ0Z_5\
        );

    \I__8467\ : InMux
    port map (
            O => \N__41979\,
            I => \N__41976\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__41976\,
            I => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\
        );

    \I__8465\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41970\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__41970\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\
        );

    \I__8463\ : CascadeMux
    port map (
            O => \N__41967\,
            I => \ppm_encoder_1.N_232_cascade_\
        );

    \I__8462\ : IoInMux
    port map (
            O => \N__41964\,
            I => \N__41961\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__8460\ : Span4Mux_s1_v
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__41955\,
            I => \N__41952\
        );

    \I__8458\ : Span4Mux_v
    port map (
            O => \N__41952\,
            I => \N__41949\
        );

    \I__8457\ : Odrv4
    port map (
            O => \N__41949\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\
        );

    \I__8456\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41941\
        );

    \I__8455\ : InMux
    port map (
            O => \N__41945\,
            I => \N__41938\
        );

    \I__8454\ : InMux
    port map (
            O => \N__41944\,
            I => \N__41935\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__41941\,
            I => \N__41932\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__41938\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__41935\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__8450\ : Odrv4
    port map (
            O => \N__41932\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__8449\ : CascadeMux
    port map (
            O => \N__41925\,
            I => \N__41922\
        );

    \I__8448\ : InMux
    port map (
            O => \N__41922\,
            I => \N__41917\
        );

    \I__8447\ : InMux
    port map (
            O => \N__41921\,
            I => \N__41914\
        );

    \I__8446\ : InMux
    port map (
            O => \N__41920\,
            I => \N__41911\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__41917\,
            I => \N__41908\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__41914\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__41911\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__8442\ : Odrv4
    port map (
            O => \N__41908\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__8441\ : InMux
    port map (
            O => \N__41901\,
            I => \N__41898\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__41898\,
            I => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\
        );

    \I__8439\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41892\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__41892\,
            I => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\
        );

    \I__8437\ : InMux
    port map (
            O => \N__41889\,
            I => \N__41886\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__41886\,
            I => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\
        );

    \I__8435\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41880\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__41880\,
            I => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\
        );

    \I__8433\ : InMux
    port map (
            O => \N__41877\,
            I => \N__41874\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__41874\,
            I => \N__41869\
        );

    \I__8431\ : InMux
    port map (
            O => \N__41873\,
            I => \N__41866\
        );

    \I__8430\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41863\
        );

    \I__8429\ : Span4Mux_v
    port map (
            O => \N__41869\,
            I => \N__41858\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__41866\,
            I => \N__41858\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__41863\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__8426\ : Odrv4
    port map (
            O => \N__41858\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__8425\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41849\
        );

    \I__8424\ : InMux
    port map (
            O => \N__41852\,
            I => \N__41845\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__41849\,
            I => \N__41842\
        );

    \I__8422\ : InMux
    port map (
            O => \N__41848\,
            I => \N__41839\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__41845\,
            I => \N__41832\
        );

    \I__8420\ : Span4Mux_v
    port map (
            O => \N__41842\,
            I => \N__41832\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__41839\,
            I => \N__41832\
        );

    \I__8418\ : Odrv4
    port map (
            O => \N__41832\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__8417\ : InMux
    port map (
            O => \N__41829\,
            I => \N__41826\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__41826\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\
        );

    \I__8415\ : InMux
    port map (
            O => \N__41823\,
            I => \N__41820\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__41820\,
            I => \ppm_encoder_1.pulses2countZ0Z_10\
        );

    \I__8413\ : InMux
    port map (
            O => \N__41817\,
            I => \N__41814\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__41814\,
            I => \N__41811\
        );

    \I__8411\ : Span4Mux_v
    port map (
            O => \N__41811\,
            I => \N__41808\
        );

    \I__8410\ : Odrv4
    port map (
            O => \N__41808\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\
        );

    \I__8409\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41802\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__41802\,
            I => \N__41799\
        );

    \I__8407\ : Span12Mux_v
    port map (
            O => \N__41799\,
            I => \N__41796\
        );

    \I__8406\ : Odrv12
    port map (
            O => \N__41796\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__41793\,
            I => \N__41790\
        );

    \I__8404\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41787\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__41787\,
            I => \ppm_encoder_1.pulses2countZ0Z_11\
        );

    \I__8402\ : InMux
    port map (
            O => \N__41784\,
            I => \N__41781\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__41781\,
            I => \N__41778\
        );

    \I__8400\ : Span4Mux_v
    port map (
            O => \N__41778\,
            I => \N__41775\
        );

    \I__8399\ : Span4Mux_v
    port map (
            O => \N__41775\,
            I => \N__41772\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__41772\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\
        );

    \I__8397\ : InMux
    port map (
            O => \N__41769\,
            I => \N__41766\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__41766\,
            I => \ppm_encoder_1.pulses2countZ0Z_12\
        );

    \I__8395\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41760\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__41760\,
            I => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\
        );

    \I__8393\ : CascadeMux
    port map (
            O => \N__41757\,
            I => \N__41754\
        );

    \I__8392\ : InMux
    port map (
            O => \N__41754\,
            I => \N__41751\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__41751\,
            I => \N__41748\
        );

    \I__8390\ : Span4Mux_v
    port map (
            O => \N__41748\,
            I => \N__41745\
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__41745\,
            I => \ppm_encoder_1.elevator_RNIH72D6Z0Z_12\
        );

    \I__8388\ : InMux
    port map (
            O => \N__41742\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_11\
        );

    \I__8387\ : CascadeMux
    port map (
            O => \N__41739\,
            I => \N__41736\
        );

    \I__8386\ : InMux
    port map (
            O => \N__41736\,
            I => \N__41733\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__41733\,
            I => \N__41730\
        );

    \I__8384\ : Odrv4
    port map (
            O => \N__41730\,
            I => \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13\
        );

    \I__8383\ : InMux
    port map (
            O => \N__41727\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_12\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__41724\,
            I => \N__41721\
        );

    \I__8381\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41718\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__41718\,
            I => \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14\
        );

    \I__8379\ : InMux
    port map (
            O => \N__41715\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_13\
        );

    \I__8378\ : InMux
    port map (
            O => \N__41712\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_14\
        );

    \I__8377\ : InMux
    port map (
            O => \N__41709\,
            I => \bfn_15_19_0_\
        );

    \I__8376\ : InMux
    port map (
            O => \N__41706\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_16\
        );

    \I__8375\ : InMux
    port map (
            O => \N__41703\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_17\
        );

    \I__8374\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41697\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__41697\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_18\
        );

    \I__8372\ : InMux
    port map (
            O => \N__41694\,
            I => \N__41691\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__41691\,
            I => \N__41688\
        );

    \I__8370\ : Odrv12
    port map (
            O => \N__41688\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0\
        );

    \I__8369\ : InMux
    port map (
            O => \N__41685\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_2\
        );

    \I__8368\ : CascadeMux
    port map (
            O => \N__41682\,
            I => \N__41679\
        );

    \I__8367\ : InMux
    port map (
            O => \N__41679\,
            I => \N__41676\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__41676\,
            I => \N__41673\
        );

    \I__8365\ : Odrv4
    port map (
            O => \N__41673\,
            I => \ppm_encoder_1.elevator_RNIFISN6Z0Z_4\
        );

    \I__8364\ : InMux
    port map (
            O => \N__41670\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_3\
        );

    \I__8363\ : CascadeMux
    port map (
            O => \N__41667\,
            I => \N__41664\
        );

    \I__8362\ : InMux
    port map (
            O => \N__41664\,
            I => \N__41661\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__41661\,
            I => \N__41658\
        );

    \I__8360\ : Odrv4
    port map (
            O => \N__41658\,
            I => \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5\
        );

    \I__8359\ : InMux
    port map (
            O => \N__41655\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_4\
        );

    \I__8358\ : CascadeMux
    port map (
            O => \N__41652\,
            I => \N__41649\
        );

    \I__8357\ : InMux
    port map (
            O => \N__41649\,
            I => \N__41646\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__41646\,
            I => \N__41643\
        );

    \I__8355\ : Odrv4
    port map (
            O => \N__41643\,
            I => \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6\
        );

    \I__8354\ : InMux
    port map (
            O => \N__41640\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_5\
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__41637\,
            I => \N__41634\
        );

    \I__8352\ : InMux
    port map (
            O => \N__41634\,
            I => \N__41631\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__41631\,
            I => \ppm_encoder_1.throttle_RNILVOO6Z0Z_7\
        );

    \I__8350\ : InMux
    port map (
            O => \N__41628\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_6\
        );

    \I__8349\ : CascadeMux
    port map (
            O => \N__41625\,
            I => \N__41622\
        );

    \I__8348\ : InMux
    port map (
            O => \N__41622\,
            I => \N__41619\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__41619\,
            I => \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8\
        );

    \I__8346\ : InMux
    port map (
            O => \N__41616\,
            I => \bfn_15_18_0_\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__41613\,
            I => \N__41610\
        );

    \I__8344\ : InMux
    port map (
            O => \N__41610\,
            I => \N__41607\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__41607\,
            I => \N__41604\
        );

    \I__8342\ : Span4Mux_v
    port map (
            O => \N__41604\,
            I => \N__41601\
        );

    \I__8341\ : Odrv4
    port map (
            O => \N__41601\,
            I => \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9\
        );

    \I__8340\ : InMux
    port map (
            O => \N__41598\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_8\
        );

    \I__8339\ : CascadeMux
    port map (
            O => \N__41595\,
            I => \N__41592\
        );

    \I__8338\ : InMux
    port map (
            O => \N__41592\,
            I => \N__41589\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__41589\,
            I => \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10\
        );

    \I__8336\ : InMux
    port map (
            O => \N__41586\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_9\
        );

    \I__8335\ : CascadeMux
    port map (
            O => \N__41583\,
            I => \N__41580\
        );

    \I__8334\ : InMux
    port map (
            O => \N__41580\,
            I => \N__41577\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__41577\,
            I => \N__41574\
        );

    \I__8332\ : Span4Mux_v
    port map (
            O => \N__41574\,
            I => \N__41571\
        );

    \I__8331\ : Odrv4
    port map (
            O => \N__41571\,
            I => \ppm_encoder_1.elevator_RNIC22D6Z0Z_11\
        );

    \I__8330\ : InMux
    port map (
            O => \N__41568\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_10\
        );

    \I__8329\ : CascadeMux
    port map (
            O => \N__41565\,
            I => \ppm_encoder_1.N_287_cascade_\
        );

    \I__8328\ : CascadeMux
    port map (
            O => \N__41562\,
            I => \N__41559\
        );

    \I__8327\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41556\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__41556\,
            I => \N__41553\
        );

    \I__8325\ : Span4Mux_v
    port map (
            O => \N__41553\,
            I => \N__41550\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__41550\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\
        );

    \I__8323\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41543\
        );

    \I__8322\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41540\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__41543\,
            I => \N__41537\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__41540\,
            I => \N__41534\
        );

    \I__8319\ : Span12Mux_v
    port map (
            O => \N__41537\,
            I => \N__41531\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__41534\,
            I => side_order_1
        );

    \I__8317\ : Odrv12
    port map (
            O => \N__41531\,
            I => side_order_1
        );

    \I__8316\ : CascadeMux
    port map (
            O => \N__41526\,
            I => \N__41523\
        );

    \I__8315\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41520\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__41520\,
            I => \N__41517\
        );

    \I__8313\ : Span4Mux_v
    port map (
            O => \N__41517\,
            I => \N__41514\
        );

    \I__8312\ : Odrv4
    port map (
            O => \N__41514\,
            I => \ppm_encoder_1.un1_aileron_cry_0_THRU_CO\
        );

    \I__8311\ : InMux
    port map (
            O => \N__41511\,
            I => \N__41506\
        );

    \I__8310\ : InMux
    port map (
            O => \N__41510\,
            I => \N__41501\
        );

    \I__8309\ : InMux
    port map (
            O => \N__41509\,
            I => \N__41501\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__41506\,
            I => \ppm_encoder_1.aileronZ0Z_1\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__41501\,
            I => \ppm_encoder_1.aileronZ0Z_1\
        );

    \I__8306\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41493\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__41493\,
            I => \N__41490\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__41490\,
            I => \ppm_encoder_1.un1_elevator_cry_0_THRU_CO\
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__41487\,
            I => \N__41484\
        );

    \I__8302\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41481\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__41481\,
            I => \N__41477\
        );

    \I__8300\ : InMux
    port map (
            O => \N__41480\,
            I => \N__41474\
        );

    \I__8299\ : Span4Mux_h
    port map (
            O => \N__41477\,
            I => \N__41469\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__41474\,
            I => \N__41469\
        );

    \I__8297\ : Span4Mux_h
    port map (
            O => \N__41469\,
            I => \N__41466\
        );

    \I__8296\ : Odrv4
    port map (
            O => \N__41466\,
            I => front_order_1
        );

    \I__8295\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41454\
        );

    \I__8294\ : InMux
    port map (
            O => \N__41462\,
            I => \N__41454\
        );

    \I__8293\ : InMux
    port map (
            O => \N__41461\,
            I => \N__41454\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__41454\,
            I => \ppm_encoder_1.elevatorZ0Z_1\
        );

    \I__8291\ : InMux
    port map (
            O => \N__41451\,
            I => \N__41448\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41445\
        );

    \I__8289\ : Span4Mux_h
    port map (
            O => \N__41445\,
            I => \N__41442\
        );

    \I__8288\ : Odrv4
    port map (
            O => \N__41442\,
            I => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\
        );

    \I__8287\ : InMux
    port map (
            O => \N__41439\,
            I => \N__41436\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__41436\,
            I => \N__41432\
        );

    \I__8285\ : InMux
    port map (
            O => \N__41435\,
            I => \N__41429\
        );

    \I__8284\ : Span4Mux_v
    port map (
            O => \N__41432\,
            I => \N__41426\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__41429\,
            I => \N__41423\
        );

    \I__8282\ : Span4Mux_h
    port map (
            O => \N__41426\,
            I => \N__41418\
        );

    \I__8281\ : Span4Mux_v
    port map (
            O => \N__41423\,
            I => \N__41418\
        );

    \I__8280\ : Span4Mux_h
    port map (
            O => \N__41418\,
            I => \N__41415\
        );

    \I__8279\ : Odrv4
    port map (
            O => \N__41415\,
            I => throttle_order_1
        );

    \I__8278\ : InMux
    port map (
            O => \N__41412\,
            I => \N__41403\
        );

    \I__8277\ : InMux
    port map (
            O => \N__41411\,
            I => \N__41403\
        );

    \I__8276\ : InMux
    port map (
            O => \N__41410\,
            I => \N__41403\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__41403\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__8274\ : CascadeMux
    port map (
            O => \N__41400\,
            I => \N__41397\
        );

    \I__8273\ : InMux
    port map (
            O => \N__41397\,
            I => \N__41394\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__41394\,
            I => \ppm_encoder_1.throttle_RNIUINC6Z0Z_1\
        );

    \I__8271\ : InMux
    port map (
            O => \N__41391\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_0\
        );

    \I__8270\ : InMux
    port map (
            O => \N__41388\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_1\
        );

    \I__8269\ : CascadeMux
    port map (
            O => \N__41385\,
            I => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\
        );

    \I__8268\ : InMux
    port map (
            O => \N__41382\,
            I => \N__41379\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__41379\,
            I => \ppm_encoder_1.un2_throttle_iv_1_4\
        );

    \I__8266\ : CascadeMux
    port map (
            O => \N__41376\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__41373\,
            I => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\
        );

    \I__8264\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41367\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__41367\,
            I => \ppm_encoder_1.un2_throttle_iv_1_5\
        );

    \I__8262\ : CascadeMux
    port map (
            O => \N__41364\,
            I => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\
        );

    \I__8261\ : CascadeMux
    port map (
            O => \N__41361\,
            I => \N__41358\
        );

    \I__8260\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41349\
        );

    \I__8259\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41345\
        );

    \I__8258\ : CascadeMux
    port map (
            O => \N__41356\,
            I => \N__41342\
        );

    \I__8257\ : CascadeMux
    port map (
            O => \N__41355\,
            I => \N__41339\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__41354\,
            I => \N__41336\
        );

    \I__8255\ : CascadeMux
    port map (
            O => \N__41353\,
            I => \N__41333\
        );

    \I__8254\ : CascadeMux
    port map (
            O => \N__41352\,
            I => \N__41329\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__41349\,
            I => \N__41324\
        );

    \I__8252\ : InMux
    port map (
            O => \N__41348\,
            I => \N__41321\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__41345\,
            I => \N__41318\
        );

    \I__8250\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41313\
        );

    \I__8249\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41313\
        );

    \I__8248\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41310\
        );

    \I__8247\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41307\
        );

    \I__8246\ : InMux
    port map (
            O => \N__41332\,
            I => \N__41304\
        );

    \I__8245\ : InMux
    port map (
            O => \N__41329\,
            I => \N__41301\
        );

    \I__8244\ : InMux
    port map (
            O => \N__41328\,
            I => \N__41298\
        );

    \I__8243\ : InMux
    port map (
            O => \N__41327\,
            I => \N__41295\
        );

    \I__8242\ : Span4Mux_h
    port map (
            O => \N__41324\,
            I => \N__41286\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41286\
        );

    \I__8240\ : Span4Mux_v
    port map (
            O => \N__41318\,
            I => \N__41286\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__41313\,
            I => \N__41286\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__41310\,
            I => \N__41281\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__41307\,
            I => \N__41281\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__41304\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__41301\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__41298\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__41295\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__41286\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__41281\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__8230\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41265\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__41265\,
            I => \ppm_encoder_1.throttle_m_1\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__41262\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\
        );

    \I__8227\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41255\
        );

    \I__8226\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41252\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__41255\,
            I => \N__41249\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__41252\,
            I => \N__41246\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__41249\,
            I => \N__41242\
        );

    \I__8222\ : Span4Mux_v
    port map (
            O => \N__41246\,
            I => \N__41239\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__41245\,
            I => \N__41236\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__41242\,
            I => \N__41232\
        );

    \I__8219\ : Span4Mux_h
    port map (
            O => \N__41239\,
            I => \N__41229\
        );

    \I__8218\ : InMux
    port map (
            O => \N__41236\,
            I => \N__41224\
        );

    \I__8217\ : InMux
    port map (
            O => \N__41235\,
            I => \N__41224\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__41232\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__41229\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__41224\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__8213\ : InMux
    port map (
            O => \N__41217\,
            I => \N__41214\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__41214\,
            I => \N__41210\
        );

    \I__8211\ : InMux
    port map (
            O => \N__41213\,
            I => \N__41207\
        );

    \I__8210\ : Span4Mux_v
    port map (
            O => \N__41210\,
            I => \N__41201\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__41207\,
            I => \N__41201\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__41206\,
            I => \N__41198\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__41201\,
            I => \N__41194\
        );

    \I__8206\ : InMux
    port map (
            O => \N__41198\,
            I => \N__41191\
        );

    \I__8205\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41188\
        );

    \I__8204\ : Span4Mux_h
    port map (
            O => \N__41194\,
            I => \N__41185\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__41191\,
            I => \N__41182\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__41188\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__8201\ : Odrv4
    port map (
            O => \N__41185\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__8200\ : Odrv12
    port map (
            O => \N__41182\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__8199\ : InMux
    port map (
            O => \N__41175\,
            I => \N__41170\
        );

    \I__8198\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41167\
        );

    \I__8197\ : InMux
    port map (
            O => \N__41173\,
            I => \N__41164\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__41170\,
            I => \N__41161\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__41167\,
            I => \N__41157\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__41164\,
            I => \N__41154\
        );

    \I__8193\ : Span4Mux_h
    port map (
            O => \N__41161\,
            I => \N__41151\
        );

    \I__8192\ : InMux
    port map (
            O => \N__41160\,
            I => \N__41148\
        );

    \I__8191\ : Odrv12
    port map (
            O => \N__41157\,
            I => \frame_decoder_CH4data_0\
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__41154\,
            I => \frame_decoder_CH4data_0\
        );

    \I__8189\ : Odrv4
    port map (
            O => \N__41151\,
            I => \frame_decoder_CH4data_0\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__41148\,
            I => \frame_decoder_CH4data_0\
        );

    \I__8187\ : CascadeMux
    port map (
            O => \N__41139\,
            I => \N__41136\
        );

    \I__8186\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41133\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__41133\,
            I => \N__41130\
        );

    \I__8184\ : Span4Mux_h
    port map (
            O => \N__41130\,
            I => \N__41127\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__41127\,
            I => \scaler_4.un2_source_data_0_cry_1_c_RNOZ0\
        );

    \I__8182\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41120\
        );

    \I__8181\ : InMux
    port map (
            O => \N__41123\,
            I => \N__41117\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__41120\,
            I => \N__41114\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__41117\,
            I => \N__41109\
        );

    \I__8178\ : Span4Mux_v
    port map (
            O => \N__41114\,
            I => \N__41109\
        );

    \I__8177\ : Span4Mux_h
    port map (
            O => \N__41109\,
            I => \N__41106\
        );

    \I__8176\ : Odrv4
    port map (
            O => \N__41106\,
            I => side_order_2
        );

    \I__8175\ : InMux
    port map (
            O => \N__41103\,
            I => \N__41099\
        );

    \I__8174\ : InMux
    port map (
            O => \N__41102\,
            I => \N__41096\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__41099\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__41096\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__41091\,
            I => \ppm_encoder_1.N_221_cascade_\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__41088\,
            I => \ppm_encoder_1.N_313_cascade_\
        );

    \I__8169\ : InMux
    port map (
            O => \N__41085\,
            I => \N__41082\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__41082\,
            I => \ppm_encoder_1.un2_throttle_iv_0_12\
        );

    \I__8167\ : InMux
    port map (
            O => \N__41079\,
            I => \N__41076\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__41076\,
            I => \ppm_encoder_1.un2_throttle_iv_1_12\
        );

    \I__8165\ : CascadeMux
    port map (
            O => \N__41073\,
            I => \N__41069\
        );

    \I__8164\ : InMux
    port map (
            O => \N__41072\,
            I => \N__41066\
        );

    \I__8163\ : InMux
    port map (
            O => \N__41069\,
            I => \N__41063\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__41066\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__41063\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__8160\ : InMux
    port map (
            O => \N__41058\,
            I => \ppm_encoder_1.un1_counter_13_cry_14\
        );

    \I__8159\ : InMux
    port map (
            O => \N__41055\,
            I => \bfn_14_25_0_\
        );

    \I__8158\ : InMux
    port map (
            O => \N__41052\,
            I => \ppm_encoder_1.un1_counter_13_cry_16\
        );

    \I__8157\ : InMux
    port map (
            O => \N__41049\,
            I => \ppm_encoder_1.un1_counter_13_cry_17\
        );

    \I__8156\ : SRMux
    port map (
            O => \N__41046\,
            I => \N__41037\
        );

    \I__8155\ : SRMux
    port map (
            O => \N__41045\,
            I => \N__41037\
        );

    \I__8154\ : SRMux
    port map (
            O => \N__41044\,
            I => \N__41037\
        );

    \I__8153\ : GlobalMux
    port map (
            O => \N__41037\,
            I => \N__41034\
        );

    \I__8152\ : gio2CtrlBuf
    port map (
            O => \N__41034\,
            I => \ppm_encoder_1.N_419_g\
        );

    \I__8151\ : IoInMux
    port map (
            O => \N__41031\,
            I => \N__41028\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__8149\ : Span4Mux_s2_v
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__8148\ : Span4Mux_v
    port map (
            O => \N__41022\,
            I => \N__41018\
        );

    \I__8147\ : InMux
    port map (
            O => \N__41021\,
            I => \N__41015\
        );

    \I__8146\ : Span4Mux_v
    port map (
            O => \N__41018\,
            I => \N__41010\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41010\
        );

    \I__8144\ : Span4Mux_h
    port map (
            O => \N__41010\,
            I => \N__41005\
        );

    \I__8143\ : CascadeMux
    port map (
            O => \N__41009\,
            I => \N__41002\
        );

    \I__8142\ : InMux
    port map (
            O => \N__41008\,
            I => \N__40999\
        );

    \I__8141\ : Span4Mux_h
    port map (
            O => \N__41005\,
            I => \N__40996\
        );

    \I__8140\ : InMux
    port map (
            O => \N__41002\,
            I => \N__40993\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__40999\,
            I => \N__40990\
        );

    \I__8138\ : Odrv4
    port map (
            O => \N__40996\,
            I => \debug_CH3_20A_c\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__40993\,
            I => \debug_CH3_20A_c\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__40990\,
            I => \debug_CH3_20A_c\
        );

    \I__8135\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40976\
        );

    \I__8134\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40971\
        );

    \I__8133\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40965\
        );

    \I__8132\ : InMux
    port map (
            O => \N__40980\,
            I => \N__40961\
        );

    \I__8131\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40958\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__40976\,
            I => \N__40955\
        );

    \I__8129\ : InMux
    port map (
            O => \N__40975\,
            I => \N__40952\
        );

    \I__8128\ : InMux
    port map (
            O => \N__40974\,
            I => \N__40949\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__40971\,
            I => \N__40946\
        );

    \I__8126\ : InMux
    port map (
            O => \N__40970\,
            I => \N__40938\
        );

    \I__8125\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40938\
        );

    \I__8124\ : InMux
    port map (
            O => \N__40968\,
            I => \N__40935\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__40965\,
            I => \N__40932\
        );

    \I__8122\ : InMux
    port map (
            O => \N__40964\,
            I => \N__40929\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__40961\,
            I => \N__40924\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__40958\,
            I => \N__40924\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__40955\,
            I => \N__40919\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__40952\,
            I => \N__40919\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__40949\,
            I => \N__40914\
        );

    \I__8116\ : Span4Mux_h
    port map (
            O => \N__40946\,
            I => \N__40914\
        );

    \I__8115\ : InMux
    port map (
            O => \N__40945\,
            I => \N__40909\
        );

    \I__8114\ : InMux
    port map (
            O => \N__40944\,
            I => \N__40909\
        );

    \I__8113\ : InMux
    port map (
            O => \N__40943\,
            I => \N__40906\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__40938\,
            I => \N__40897\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__40935\,
            I => \N__40897\
        );

    \I__8110\ : Span4Mux_v
    port map (
            O => \N__40932\,
            I => \N__40897\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__40929\,
            I => \N__40897\
        );

    \I__8108\ : Span4Mux_v
    port map (
            O => \N__40924\,
            I => \N__40894\
        );

    \I__8107\ : Span4Mux_v
    port map (
            O => \N__40919\,
            I => \N__40891\
        );

    \I__8106\ : Span4Mux_h
    port map (
            O => \N__40914\,
            I => \N__40882\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__40909\,
            I => \N__40882\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__40906\,
            I => \N__40882\
        );

    \I__8103\ : Span4Mux_v
    port map (
            O => \N__40897\,
            I => \N__40882\
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__40894\,
            I => uart_drone_data_rdy
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__40891\,
            I => uart_drone_data_rdy
        );

    \I__8100\ : Odrv4
    port map (
            O => \N__40882\,
            I => uart_drone_data_rdy
        );

    \I__8099\ : SRMux
    port map (
            O => \N__40875\,
            I => \N__40872\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__40872\,
            I => \N__40868\
        );

    \I__8097\ : SRMux
    port map (
            O => \N__40871\,
            I => \N__40865\
        );

    \I__8096\ : Span4Mux_v
    port map (
            O => \N__40868\,
            I => \N__40860\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__40865\,
            I => \N__40860\
        );

    \I__8094\ : Span4Mux_v
    port map (
            O => \N__40860\,
            I => \N__40857\
        );

    \I__8093\ : Span4Mux_h
    port map (
            O => \N__40857\,
            I => \N__40854\
        );

    \I__8092\ : Odrv4
    port map (
            O => \N__40854\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__8091\ : InMux
    port map (
            O => \N__40851\,
            I => \N__40846\
        );

    \I__8090\ : InMux
    port map (
            O => \N__40850\,
            I => \N__40843\
        );

    \I__8089\ : InMux
    port map (
            O => \N__40849\,
            I => \N__40840\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__40846\,
            I => \N__40837\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__40843\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__40840\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__40837\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__8084\ : InMux
    port map (
            O => \N__40830\,
            I => \ppm_encoder_1.un1_counter_13_cry_4\
        );

    \I__8083\ : InMux
    port map (
            O => \N__40827\,
            I => \ppm_encoder_1.un1_counter_13_cry_5\
        );

    \I__8082\ : InMux
    port map (
            O => \N__40824\,
            I => \ppm_encoder_1.un1_counter_13_cry_6\
        );

    \I__8081\ : InMux
    port map (
            O => \N__40821\,
            I => \bfn_14_24_0_\
        );

    \I__8080\ : InMux
    port map (
            O => \N__40818\,
            I => \ppm_encoder_1.un1_counter_13_cry_8\
        );

    \I__8079\ : InMux
    port map (
            O => \N__40815\,
            I => \ppm_encoder_1.un1_counter_13_cry_9\
        );

    \I__8078\ : InMux
    port map (
            O => \N__40812\,
            I => \ppm_encoder_1.un1_counter_13_cry_10\
        );

    \I__8077\ : InMux
    port map (
            O => \N__40809\,
            I => \ppm_encoder_1.un1_counter_13_cry_11\
        );

    \I__8076\ : InMux
    port map (
            O => \N__40806\,
            I => \ppm_encoder_1.un1_counter_13_cry_12\
        );

    \I__8075\ : InMux
    port map (
            O => \N__40803\,
            I => \ppm_encoder_1.un1_counter_13_cry_13\
        );

    \I__8074\ : InMux
    port map (
            O => \N__40800\,
            I => \N__40797\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__40797\,
            I => \N__40794\
        );

    \I__8072\ : Odrv4
    port map (
            O => \N__40794\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\
        );

    \I__8071\ : InMux
    port map (
            O => \N__40791\,
            I => \N__40788\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__40788\,
            I => \N__40785\
        );

    \I__8069\ : Span12Mux_s9_v
    port map (
            O => \N__40785\,
            I => \N__40782\
        );

    \I__8068\ : Odrv12
    port map (
            O => \N__40782\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\
        );

    \I__8067\ : InMux
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__40776\,
            I => \ppm_encoder_1.pulses2countZ0Z_0\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__40773\,
            I => \N__40770\
        );

    \I__8064\ : InMux
    port map (
            O => \N__40770\,
            I => \N__40767\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__40767\,
            I => \ppm_encoder_1.pulses2countZ0Z_1\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__40764\,
            I => \N__40760\
        );

    \I__8061\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40757\
        );

    \I__8060\ : InMux
    port map (
            O => \N__40760\,
            I => \N__40754\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__40757\,
            I => \N__40749\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__40754\,
            I => \N__40749\
        );

    \I__8057\ : Span4Mux_v
    port map (
            O => \N__40749\,
            I => \N__40746\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__40746\,
            I => \ppm_encoder_1.N_2150_i\
        );

    \I__8055\ : InMux
    port map (
            O => \N__40743\,
            I => \ppm_encoder_1.un1_counter_13_cry_0\
        );

    \I__8054\ : InMux
    port map (
            O => \N__40740\,
            I => \ppm_encoder_1.un1_counter_13_cry_1\
        );

    \I__8053\ : InMux
    port map (
            O => \N__40737\,
            I => \ppm_encoder_1.un1_counter_13_cry_2\
        );

    \I__8052\ : InMux
    port map (
            O => \N__40734\,
            I => \ppm_encoder_1.un1_counter_13_cry_3\
        );

    \I__8051\ : CascadeMux
    port map (
            O => \N__40731\,
            I => \N__40728\
        );

    \I__8050\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40725\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__40725\,
            I => \N__40722\
        );

    \I__8048\ : Span4Mux_v
    port map (
            O => \N__40722\,
            I => \N__40718\
        );

    \I__8047\ : InMux
    port map (
            O => \N__40721\,
            I => \N__40715\
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__40718\,
            I => \drone_H_disp_front_13\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__40715\,
            I => \drone_H_disp_front_13\
        );

    \I__8044\ : InMux
    port map (
            O => \N__40710\,
            I => \N__40707\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__40707\,
            I => \N__40704\
        );

    \I__8042\ : Span4Mux_v
    port map (
            O => \N__40704\,
            I => \N__40701\
        );

    \I__8041\ : Odrv4
    port map (
            O => \N__40701\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\
        );

    \I__8040\ : InMux
    port map (
            O => \N__40698\,
            I => \N__40695\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__40695\,
            I => \N__40692\
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__40692\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\
        );

    \I__8037\ : InMux
    port map (
            O => \N__40689\,
            I => \N__40686\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__40686\,
            I => \ppm_encoder_1.pulses2countZ0Z_6\
        );

    \I__8035\ : InMux
    port map (
            O => \N__40683\,
            I => \N__40680\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__40680\,
            I => \N__40677\
        );

    \I__8033\ : Odrv4
    port map (
            O => \N__40677\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\
        );

    \I__8032\ : InMux
    port map (
            O => \N__40674\,
            I => \N__40671\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__40671\,
            I => \N__40668\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__40668\,
            I => \N__40665\
        );

    \I__8029\ : Odrv4
    port map (
            O => \N__40665\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__40662\,
            I => \N__40659\
        );

    \I__8027\ : InMux
    port map (
            O => \N__40659\,
            I => \N__40656\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__40656\,
            I => \ppm_encoder_1.pulses2countZ0Z_7\
        );

    \I__8025\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40650\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__40650\,
            I => \N__40647\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__40647\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\
        );

    \I__8022\ : InMux
    port map (
            O => \N__40644\,
            I => \N__40641\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__40641\,
            I => \ppm_encoder_1.pulses2countZ0Z_13\
        );

    \I__8020\ : InMux
    port map (
            O => \N__40638\,
            I => \N__40635\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__40635\,
            I => \N__40632\
        );

    \I__8018\ : Span4Mux_v
    port map (
            O => \N__40632\,
            I => \N__40629\
        );

    \I__8017\ : Odrv4
    port map (
            O => \N__40629\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\
        );

    \I__8016\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40623\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__40623\,
            I => \ppm_encoder_1.pulses2countZ0Z_8\
        );

    \I__8014\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40617\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__40617\,
            I => \N__40614\
        );

    \I__8012\ : Odrv12
    port map (
            O => \N__40614\,
            I => \ppm_encoder_1.pulses2countZ0Z_9\
        );

    \I__8011\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40607\
        );

    \I__8010\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40603\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__40607\,
            I => \N__40600\
        );

    \I__8008\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40597\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__40603\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__8006\ : Odrv4
    port map (
            O => \N__40600\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__40597\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__8004\ : CascadeMux
    port map (
            O => \N__40590\,
            I => \ppm_encoder_1.un2_throttle_iv_1_10_cascade_\
        );

    \I__8003\ : InMux
    port map (
            O => \N__40587\,
            I => \N__40584\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__40584\,
            I => \ppm_encoder_1.un2_throttle_iv_0_10\
        );

    \I__8001\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40578\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__40578\,
            I => \N__40573\
        );

    \I__7999\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40570\
        );

    \I__7998\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40567\
        );

    \I__7997\ : Span4Mux_v
    port map (
            O => \N__40573\,
            I => \N__40562\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__40570\,
            I => \N__40562\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__40567\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__7994\ : Odrv4
    port map (
            O => \N__40562\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__7993\ : InMux
    port map (
            O => \N__40557\,
            I => \N__40554\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__40554\,
            I => \N__40549\
        );

    \I__7991\ : InMux
    port map (
            O => \N__40553\,
            I => \N__40546\
        );

    \I__7990\ : CascadeMux
    port map (
            O => \N__40552\,
            I => \N__40543\
        );

    \I__7989\ : Span4Mux_v
    port map (
            O => \N__40549\,
            I => \N__40538\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__40546\,
            I => \N__40538\
        );

    \I__7987\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40535\
        );

    \I__7986\ : Span4Mux_h
    port map (
            O => \N__40538\,
            I => \N__40532\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__40535\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__40532\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__7983\ : InMux
    port map (
            O => \N__40527\,
            I => \N__40521\
        );

    \I__7982\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40521\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__40521\,
            I => \N__40517\
        );

    \I__7980\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40514\
        );

    \I__7979\ : Span4Mux_h
    port map (
            O => \N__40517\,
            I => \N__40511\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__40514\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__7977\ : Odrv4
    port map (
            O => \N__40511\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__40506\,
            I => \ppm_encoder_1.N_296_cascade_\
        );

    \I__7975\ : InMux
    port map (
            O => \N__40503\,
            I => \N__40497\
        );

    \I__7974\ : InMux
    port map (
            O => \N__40502\,
            I => \N__40497\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__40497\,
            I => \N__40493\
        );

    \I__7972\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40490\
        );

    \I__7971\ : Span4Mux_h
    port map (
            O => \N__40493\,
            I => \N__40487\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__40490\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__40487\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__7968\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40479\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__40479\,
            I => \ppm_encoder_1.un2_throttle_iv_1_8\
        );

    \I__7966\ : InMux
    port map (
            O => \N__40476\,
            I => \N__40470\
        );

    \I__7965\ : InMux
    port map (
            O => \N__40475\,
            I => \N__40470\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__40470\,
            I => \N__40466\
        );

    \I__7963\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40463\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__40466\,
            I => \N__40460\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__40463\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__7960\ : Odrv4
    port map (
            O => \N__40460\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__7959\ : InMux
    port map (
            O => \N__40455\,
            I => \N__40450\
        );

    \I__7958\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40445\
        );

    \I__7957\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40445\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__40450\,
            I => \N__40442\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__40445\,
            I => \N__40439\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__40442\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__40439\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__40434\,
            I => \ppm_encoder_1.N_294_cascade_\
        );

    \I__7951\ : InMux
    port map (
            O => \N__40431\,
            I => \N__40428\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__40428\,
            I => \N__40425\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__40425\,
            I => \N__40422\
        );

    \I__7948\ : Odrv4
    port map (
            O => \N__40422\,
            I => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\
        );

    \I__7947\ : InMux
    port map (
            O => \N__40419\,
            I => \N__40410\
        );

    \I__7946\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40410\
        );

    \I__7945\ : InMux
    port map (
            O => \N__40417\,
            I => \N__40410\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__40410\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__40407\,
            I => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\
        );

    \I__7942\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40401\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__40401\,
            I => \ppm_encoder_1.un2_throttle_iv_1_14\
        );

    \I__7940\ : InMux
    port map (
            O => \N__40398\,
            I => \N__40392\
        );

    \I__7939\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40392\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__40392\,
            I => \N__40389\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__40389\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__7936\ : InMux
    port map (
            O => \N__40386\,
            I => \N__40382\
        );

    \I__7935\ : InMux
    port map (
            O => \N__40385\,
            I => \N__40379\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__40382\,
            I => \N__40374\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__40379\,
            I => \N__40374\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__40374\,
            I => \N__40371\
        );

    \I__7931\ : Odrv4
    port map (
            O => \N__40371\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__7930\ : CascadeMux
    port map (
            O => \N__40368\,
            I => \ppm_encoder_1.N_300_cascade_\
        );

    \I__7929\ : InMux
    port map (
            O => \N__40365\,
            I => \N__40359\
        );

    \I__7928\ : InMux
    port map (
            O => \N__40364\,
            I => \N__40359\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__40359\,
            I => \N__40356\
        );

    \I__7926\ : Odrv12
    port map (
            O => \N__40356\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__7925\ : CascadeMux
    port map (
            O => \N__40353\,
            I => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\
        );

    \I__7924\ : InMux
    port map (
            O => \N__40350\,
            I => \N__40347\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__40347\,
            I => \ppm_encoder_1.un2_throttle_iv_1_7\
        );

    \I__7922\ : InMux
    port map (
            O => \N__40344\,
            I => \N__40337\
        );

    \I__7921\ : InMux
    port map (
            O => \N__40343\,
            I => \N__40337\
        );

    \I__7920\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40334\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40331\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__40334\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__7917\ : Odrv12
    port map (
            O => \N__40331\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__7916\ : CascadeMux
    port map (
            O => \N__40326\,
            I => \ppm_encoder_1.N_293_cascade_\
        );

    \I__7915\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40320\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__40320\,
            I => \N__40317\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__40317\,
            I => \N__40314\
        );

    \I__7912\ : Odrv4
    port map (
            O => \N__40314\,
            I => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\
        );

    \I__7911\ : InMux
    port map (
            O => \N__40311\,
            I => \N__40302\
        );

    \I__7910\ : InMux
    port map (
            O => \N__40310\,
            I => \N__40302\
        );

    \I__7909\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40302\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__40302\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__7907\ : InMux
    port map (
            O => \N__40299\,
            I => \N__40296\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__40296\,
            I => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\
        );

    \I__7905\ : InMux
    port map (
            O => \N__40293\,
            I => \N__40288\
        );

    \I__7904\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40285\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__40291\,
            I => \N__40282\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__40288\,
            I => \N__40277\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__40285\,
            I => \N__40277\
        );

    \I__7900\ : InMux
    port map (
            O => \N__40282\,
            I => \N__40274\
        );

    \I__7899\ : Span4Mux_v
    port map (
            O => \N__40277\,
            I => \N__40271\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__40274\,
            I => front_order_7
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__40271\,
            I => front_order_7
        );

    \I__7896\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40257\
        );

    \I__7895\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40257\
        );

    \I__7894\ : InMux
    port map (
            O => \N__40264\,
            I => \N__40257\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__40257\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__7892\ : CascadeMux
    port map (
            O => \N__40254\,
            I => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\
        );

    \I__7891\ : CascadeMux
    port map (
            O => \N__40251\,
            I => \N__40246\
        );

    \I__7890\ : InMux
    port map (
            O => \N__40250\,
            I => \N__40241\
        );

    \I__7889\ : InMux
    port map (
            O => \N__40249\,
            I => \N__40241\
        );

    \I__7888\ : InMux
    port map (
            O => \N__40246\,
            I => \N__40238\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__40241\,
            I => \N__40235\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__40238\,
            I => \N__40230\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__40235\,
            I => \N__40230\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__40230\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__7883\ : InMux
    port map (
            O => \N__40227\,
            I => \N__40222\
        );

    \I__7882\ : InMux
    port map (
            O => \N__40226\,
            I => \N__40217\
        );

    \I__7881\ : InMux
    port map (
            O => \N__40225\,
            I => \N__40217\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__40222\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__40217\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__7878\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__40209\,
            I => \ppm_encoder_1.N_295\
        );

    \I__7876\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40199\
        );

    \I__7875\ : InMux
    port map (
            O => \N__40205\,
            I => \N__40199\
        );

    \I__7874\ : InMux
    port map (
            O => \N__40204\,
            I => \N__40196\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__40199\,
            I => \N__40193\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__40196\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__7871\ : Odrv12
    port map (
            O => \N__40193\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__7870\ : InMux
    port map (
            O => \N__40188\,
            I => \N__40185\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__40185\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\
        );

    \I__7868\ : CascadeMux
    port map (
            O => \N__40182\,
            I => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\
        );

    \I__7867\ : InMux
    port map (
            O => \N__40179\,
            I => \N__40176\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__40176\,
            I => \ppm_encoder_1.un2_throttle_iv_1_6\
        );

    \I__7865\ : InMux
    port map (
            O => \N__40173\,
            I => \N__40166\
        );

    \I__7864\ : InMux
    port map (
            O => \N__40172\,
            I => \N__40166\
        );

    \I__7863\ : CascadeMux
    port map (
            O => \N__40171\,
            I => \N__40163\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__40166\,
            I => \N__40160\
        );

    \I__7861\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40157\
        );

    \I__7860\ : Span4Mux_h
    port map (
            O => \N__40160\,
            I => \N__40154\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__40157\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__7858\ : Odrv4
    port map (
            O => \N__40154\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__40149\,
            I => \N__40145\
        );

    \I__7856\ : CascadeMux
    port map (
            O => \N__40148\,
            I => \N__40141\
        );

    \I__7855\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40138\
        );

    \I__7854\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40133\
        );

    \I__7853\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40133\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__40138\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__40133\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__7850\ : CascadeMux
    port map (
            O => \N__40128\,
            I => \ppm_encoder_1.N_292_cascade_\
        );

    \I__7849\ : InMux
    port map (
            O => \N__40125\,
            I => \N__40122\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__40122\,
            I => \N__40119\
        );

    \I__7847\ : Span4Mux_h
    port map (
            O => \N__40119\,
            I => \N__40116\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__40116\,
            I => \ppm_encoder_1.un1_aileron_cry_5_THRU_CO\
        );

    \I__7845\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40104\
        );

    \I__7844\ : InMux
    port map (
            O => \N__40112\,
            I => \N__40104\
        );

    \I__7843\ : InMux
    port map (
            O => \N__40111\,
            I => \N__40104\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__40104\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__7841\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40094\
        );

    \I__7840\ : InMux
    port map (
            O => \N__40100\,
            I => \N__40094\
        );

    \I__7839\ : InMux
    port map (
            O => \N__40099\,
            I => \N__40091\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__40094\,
            I => \N__40088\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__40091\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__40088\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__40083\,
            I => \ppm_encoder_1.N_297_cascade_\
        );

    \I__7834\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40077\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__40077\,
            I => \N__40074\
        );

    \I__7832\ : Span4Mux_h
    port map (
            O => \N__40074\,
            I => \N__40071\
        );

    \I__7831\ : Span4Mux_v
    port map (
            O => \N__40071\,
            I => \N__40068\
        );

    \I__7830\ : Odrv4
    port map (
            O => \N__40068\,
            I => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\
        );

    \I__7829\ : InMux
    port map (
            O => \N__40065\,
            I => \N__40056\
        );

    \I__7828\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40056\
        );

    \I__7827\ : InMux
    port map (
            O => \N__40063\,
            I => \N__40056\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__40056\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__7825\ : InMux
    port map (
            O => \N__40053\,
            I => \N__40050\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__40050\,
            I => \N__40047\
        );

    \I__7823\ : Span4Mux_v
    port map (
            O => \N__40047\,
            I => \N__40042\
        );

    \I__7822\ : InMux
    port map (
            O => \N__40046\,
            I => \N__40039\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__40045\,
            I => \N__40036\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__40042\,
            I => \N__40033\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__40039\,
            I => \N__40030\
        );

    \I__7818\ : InMux
    port map (
            O => \N__40036\,
            I => \N__40027\
        );

    \I__7817\ : Sp12to4
    port map (
            O => \N__40033\,
            I => \N__40022\
        );

    \I__7816\ : Span12Mux_v
    port map (
            O => \N__40030\,
            I => \N__40022\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__40027\,
            I => throttle_order_11
        );

    \I__7814\ : Odrv12
    port map (
            O => \N__40022\,
            I => throttle_order_11
        );

    \I__7813\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40014\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__40014\,
            I => \N__40011\
        );

    \I__7811\ : Span4Mux_v
    port map (
            O => \N__40011\,
            I => \N__40008\
        );

    \I__7810\ : Odrv4
    port map (
            O => \N__40008\,
            I => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__40005\,
            I => \N__40002\
        );

    \I__7808\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39997\
        );

    \I__7807\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39992\
        );

    \I__7806\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39992\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__39997\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__39992\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__7803\ : CascadeMux
    port map (
            O => \N__39987\,
            I => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\
        );

    \I__7802\ : CascadeMux
    port map (
            O => \N__39984\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\
        );

    \I__7801\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39975\
        );

    \I__7800\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39975\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__39975\,
            I => \N__39971\
        );

    \I__7798\ : InMux
    port map (
            O => \N__39974\,
            I => \N__39968\
        );

    \I__7797\ : Span4Mux_h
    port map (
            O => \N__39971\,
            I => \N__39965\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__39968\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__7795\ : Odrv4
    port map (
            O => \N__39965\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__7794\ : InMux
    port map (
            O => \N__39960\,
            I => \N__39957\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__39957\,
            I => \ppm_encoder_1.un2_throttle_iv_1_9\
        );

    \I__7792\ : InMux
    port map (
            O => \N__39954\,
            I => \N__39947\
        );

    \I__7791\ : InMux
    port map (
            O => \N__39953\,
            I => \N__39947\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__39952\,
            I => \N__39944\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__39947\,
            I => \N__39941\
        );

    \I__7788\ : InMux
    port map (
            O => \N__39944\,
            I => \N__39938\
        );

    \I__7787\ : Span4Mux_h
    port map (
            O => \N__39941\,
            I => \N__39935\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__39938\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__39935\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__7784\ : CascadeMux
    port map (
            O => \N__39930\,
            I => \ppm_encoder_1.N_298_cascade_\
        );

    \I__7783\ : CascadeMux
    port map (
            O => \N__39927\,
            I => \N__39924\
        );

    \I__7782\ : InMux
    port map (
            O => \N__39924\,
            I => \N__39921\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__39921\,
            I => \N__39918\
        );

    \I__7780\ : Span4Mux_h
    port map (
            O => \N__39918\,
            I => \N__39915\
        );

    \I__7779\ : Span4Mux_v
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__7778\ : Odrv4
    port map (
            O => \N__39912\,
            I => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\
        );

    \I__7777\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39900\
        );

    \I__7776\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39900\
        );

    \I__7775\ : InMux
    port map (
            O => \N__39907\,
            I => \N__39900\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__39900\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__7773\ : InMux
    port map (
            O => \N__39897\,
            I => \N__39894\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__39894\,
            I => \N__39891\
        );

    \I__7771\ : Span4Mux_h
    port map (
            O => \N__39891\,
            I => \N__39887\
        );

    \I__7770\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39884\
        );

    \I__7769\ : Sp12to4
    port map (
            O => \N__39887\,
            I => \N__39879\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__39884\,
            I => \N__39879\
        );

    \I__7767\ : Span12Mux_v
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__7766\ : Odrv12
    port map (
            O => \N__39876\,
            I => front_order_12
        );

    \I__7765\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39870\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__39870\,
            I => \N__39867\
        );

    \I__7763\ : Span4Mux_v
    port map (
            O => \N__39867\,
            I => \N__39864\
        );

    \I__7762\ : Odrv4
    port map (
            O => \N__39864\,
            I => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\
        );

    \I__7761\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39852\
        );

    \I__7760\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39852\
        );

    \I__7759\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39852\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__39852\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__7757\ : CascadeMux
    port map (
            O => \N__39849\,
            I => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\
        );

    \I__7756\ : InMux
    port map (
            O => \N__39846\,
            I => \N__39843\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__39843\,
            I => \ppm_encoder_1.un2_throttle_iv_1_11\
        );

    \I__7754\ : CEMux
    port map (
            O => \N__39840\,
            I => \N__39837\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__39837\,
            I => \N__39834\
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__39834\,
            I => \pid_alt.state_1_0_0\
        );

    \I__7751\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39827\
        );

    \I__7750\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39824\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__39827\,
            I => \N__39821\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__39824\,
            I => \N__39818\
        );

    \I__7747\ : Odrv4
    port map (
            O => \N__39821\,
            I => scaler_4_data_9
        );

    \I__7746\ : Odrv4
    port map (
            O => \N__39818\,
            I => scaler_4_data_9
        );

    \I__7745\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39810\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__39810\,
            I => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\
        );

    \I__7743\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39804\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__39804\,
            I => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\
        );

    \I__7741\ : InMux
    port map (
            O => \N__39801\,
            I => \N__39797\
        );

    \I__7740\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39794\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__39797\,
            I => \N__39791\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__39794\,
            I => \N__39788\
        );

    \I__7737\ : Odrv4
    port map (
            O => \N__39791\,
            I => scaler_4_data_8
        );

    \I__7736\ : Odrv4
    port map (
            O => \N__39788\,
            I => scaler_4_data_8
        );

    \I__7735\ : InMux
    port map (
            O => \N__39783\,
            I => \N__39779\
        );

    \I__7734\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39776\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__39779\,
            I => \N__39771\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__39776\,
            I => \N__39771\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__39771\,
            I => scaler_4_data_10
        );

    \I__7730\ : InMux
    port map (
            O => \N__39768\,
            I => \N__39765\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__39765\,
            I => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\
        );

    \I__7728\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39758\
        );

    \I__7727\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39755\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__39758\,
            I => \N__39752\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__39755\,
            I => \N__39749\
        );

    \I__7724\ : Odrv4
    port map (
            O => \N__39752\,
            I => scaler_4_data_13
        );

    \I__7723\ : Odrv4
    port map (
            O => \N__39749\,
            I => scaler_4_data_13
        );

    \I__7722\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__39741\,
            I => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\
        );

    \I__7720\ : CascadeMux
    port map (
            O => \N__39738\,
            I => \N__39732\
        );

    \I__7719\ : InMux
    port map (
            O => \N__39737\,
            I => \N__39706\
        );

    \I__7718\ : InMux
    port map (
            O => \N__39736\,
            I => \N__39706\
        );

    \I__7717\ : InMux
    port map (
            O => \N__39735\,
            I => \N__39706\
        );

    \I__7716\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39706\
        );

    \I__7715\ : InMux
    port map (
            O => \N__39731\,
            I => \N__39706\
        );

    \I__7714\ : InMux
    port map (
            O => \N__39730\,
            I => \N__39701\
        );

    \I__7713\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39701\
        );

    \I__7712\ : InMux
    port map (
            O => \N__39728\,
            I => \N__39686\
        );

    \I__7711\ : InMux
    port map (
            O => \N__39727\,
            I => \N__39686\
        );

    \I__7710\ : InMux
    port map (
            O => \N__39726\,
            I => \N__39686\
        );

    \I__7709\ : InMux
    port map (
            O => \N__39725\,
            I => \N__39686\
        );

    \I__7708\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39686\
        );

    \I__7707\ : InMux
    port map (
            O => \N__39723\,
            I => \N__39686\
        );

    \I__7706\ : InMux
    port map (
            O => \N__39722\,
            I => \N__39686\
        );

    \I__7705\ : InMux
    port map (
            O => \N__39721\,
            I => \N__39679\
        );

    \I__7704\ : InMux
    port map (
            O => \N__39720\,
            I => \N__39679\
        );

    \I__7703\ : InMux
    port map (
            O => \N__39719\,
            I => \N__39679\
        );

    \I__7702\ : InMux
    port map (
            O => \N__39718\,
            I => \N__39672\
        );

    \I__7701\ : InMux
    port map (
            O => \N__39717\,
            I => \N__39669\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__39706\,
            I => \N__39666\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__39701\,
            I => \N__39659\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__39686\,
            I => \N__39659\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__39679\,
            I => \N__39659\
        );

    \I__7696\ : InMux
    port map (
            O => \N__39678\,
            I => \N__39656\
        );

    \I__7695\ : InMux
    port map (
            O => \N__39677\,
            I => \N__39653\
        );

    \I__7694\ : InMux
    port map (
            O => \N__39676\,
            I => \N__39650\
        );

    \I__7693\ : InMux
    port map (
            O => \N__39675\,
            I => \N__39647\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__39672\,
            I => \N__39642\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__39669\,
            I => \N__39642\
        );

    \I__7690\ : Span4Mux_v
    port map (
            O => \N__39666\,
            I => \N__39635\
        );

    \I__7689\ : Span4Mux_v
    port map (
            O => \N__39659\,
            I => \N__39635\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__39656\,
            I => \N__39635\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__39653\,
            I => \N__39632\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__39650\,
            I => \N__39629\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__39647\,
            I => \N__39626\
        );

    \I__7684\ : Span4Mux_v
    port map (
            O => \N__39642\,
            I => \N__39623\
        );

    \I__7683\ : Span4Mux_h
    port map (
            O => \N__39635\,
            I => \N__39618\
        );

    \I__7682\ : Span4Mux_h
    port map (
            O => \N__39632\,
            I => \N__39618\
        );

    \I__7681\ : Span4Mux_v
    port map (
            O => \N__39629\,
            I => \N__39615\
        );

    \I__7680\ : Span12Mux_h
    port map (
            O => \N__39626\,
            I => \N__39612\
        );

    \I__7679\ : Span4Mux_v
    port map (
            O => \N__39623\,
            I => \N__39607\
        );

    \I__7678\ : Span4Mux_h
    port map (
            O => \N__39618\,
            I => \N__39607\
        );

    \I__7677\ : Odrv4
    port map (
            O => \N__39615\,
            I => \pid_alt.N_72_i\
        );

    \I__7676\ : Odrv12
    port map (
            O => \N__39612\,
            I => \pid_alt.N_72_i\
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__39607\,
            I => \pid_alt.N_72_i\
        );

    \I__7674\ : InMux
    port map (
            O => \N__39600\,
            I => \N__39596\
        );

    \I__7673\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39592\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__39596\,
            I => \N__39589\
        );

    \I__7671\ : CascadeMux
    port map (
            O => \N__39595\,
            I => \N__39585\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__39592\,
            I => \N__39581\
        );

    \I__7669\ : Sp12to4
    port map (
            O => \N__39589\,
            I => \N__39578\
        );

    \I__7668\ : InMux
    port map (
            O => \N__39588\,
            I => \N__39575\
        );

    \I__7667\ : InMux
    port map (
            O => \N__39585\,
            I => \N__39572\
        );

    \I__7666\ : InMux
    port map (
            O => \N__39584\,
            I => \N__39569\
        );

    \I__7665\ : Sp12to4
    port map (
            O => \N__39581\,
            I => \N__39564\
        );

    \I__7664\ : Span12Mux_s9_v
    port map (
            O => \N__39578\,
            I => \N__39564\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__39575\,
            I => \N__39559\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__39572\,
            I => \N__39559\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__39569\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__7660\ : Odrv12
    port map (
            O => \N__39564\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__7659\ : Odrv4
    port map (
            O => \N__39559\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__39552\,
            I => \N__39548\
        );

    \I__7657\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39545\
        );

    \I__7656\ : InMux
    port map (
            O => \N__39548\,
            I => \N__39542\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__39545\,
            I => \N__39537\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__39542\,
            I => \N__39537\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__39537\,
            I => scaler_4_data_11
        );

    \I__7652\ : InMux
    port map (
            O => \N__39534\,
            I => \N__39531\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__39531\,
            I => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\
        );

    \I__7650\ : InMux
    port map (
            O => \N__39528\,
            I => \N__39524\
        );

    \I__7649\ : InMux
    port map (
            O => \N__39527\,
            I => \N__39521\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__39524\,
            I => \N__39518\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__39521\,
            I => scaler_4_data_12
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__39518\,
            I => scaler_4_data_12
        );

    \I__7645\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39510\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__39510\,
            I => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\
        );

    \I__7643\ : InMux
    port map (
            O => \N__39507\,
            I => \N__39504\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__39504\,
            I => \N__39501\
        );

    \I__7641\ : Odrv12
    port map (
            O => \N__39501\,
            I => \drone_H_disp_front_i_13\
        );

    \I__7640\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39495\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__39495\,
            I => \N__39491\
        );

    \I__7638\ : InMux
    port map (
            O => \N__39494\,
            I => \N__39488\
        );

    \I__7637\ : Span4Mux_s2_h
    port map (
            O => \N__39491\,
            I => \N__39485\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__39488\,
            I => \N__39482\
        );

    \I__7635\ : Span4Mux_v
    port map (
            O => \N__39485\,
            I => \N__39479\
        );

    \I__7634\ : Span4Mux_s3_h
    port map (
            O => \N__39482\,
            I => \N__39476\
        );

    \I__7633\ : Span4Mux_h
    port map (
            O => \N__39479\,
            I => \N__39473\
        );

    \I__7632\ : Span4Mux_h
    port map (
            O => \N__39476\,
            I => \N__39470\
        );

    \I__7631\ : Span4Mux_h
    port map (
            O => \N__39473\,
            I => \N__39467\
        );

    \I__7630\ : Span4Mux_h
    port map (
            O => \N__39470\,
            I => \N__39462\
        );

    \I__7629\ : Span4Mux_h
    port map (
            O => \N__39467\,
            I => \N__39462\
        );

    \I__7628\ : Odrv4
    port map (
            O => \N__39462\,
            I => \pid_front.error_14\
        );

    \I__7627\ : InMux
    port map (
            O => \N__39459\,
            I => \pid_front.error_cry_9\
        );

    \I__7626\ : InMux
    port map (
            O => \N__39456\,
            I => \pid_front.error_cry_10\
        );

    \I__7625\ : InMux
    port map (
            O => \N__39453\,
            I => \N__39449\
        );

    \I__7624\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39446\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39443\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__39446\,
            I => \N__39440\
        );

    \I__7621\ : Span4Mux_s2_h
    port map (
            O => \N__39443\,
            I => \N__39437\
        );

    \I__7620\ : Span4Mux_s3_h
    port map (
            O => \N__39440\,
            I => \N__39434\
        );

    \I__7619\ : Sp12to4
    port map (
            O => \N__39437\,
            I => \N__39431\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__39434\,
            I => \N__39428\
        );

    \I__7617\ : Span12Mux_v
    port map (
            O => \N__39431\,
            I => \N__39425\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__39428\,
            I => \N__39422\
        );

    \I__7615\ : Odrv12
    port map (
            O => \N__39425\,
            I => \pid_front.error_15\
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__39422\,
            I => \pid_front.error_15\
        );

    \I__7613\ : InMux
    port map (
            O => \N__39417\,
            I => \N__39414\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__39414\,
            I => \dron_frame_decoder_1.drone_H_disp_front_10\
        );

    \I__7611\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39405\
        );

    \I__7610\ : InMux
    port map (
            O => \N__39410\,
            I => \N__39405\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__39405\,
            I => \drone_H_disp_front_11\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__39402\,
            I => \N__39399\
        );

    \I__7607\ : InMux
    port map (
            O => \N__39399\,
            I => \N__39394\
        );

    \I__7606\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39389\
        );

    \I__7605\ : InMux
    port map (
            O => \N__39397\,
            I => \N__39389\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__39394\,
            I => \drone_H_disp_front_12\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__39389\,
            I => \drone_H_disp_front_12\
        );

    \I__7602\ : CascadeMux
    port map (
            O => \N__39384\,
            I => \N__39380\
        );

    \I__7601\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39375\
        );

    \I__7600\ : InMux
    port map (
            O => \N__39380\,
            I => \N__39375\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__39375\,
            I => \N__39372\
        );

    \I__7598\ : Odrv4
    port map (
            O => \N__39372\,
            I => \drone_H_disp_front_14\
        );

    \I__7597\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39366\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__39366\,
            I => \N__39363\
        );

    \I__7595\ : Odrv4
    port map (
            O => \N__39363\,
            I => \drone_H_disp_front_15\
        );

    \I__7594\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39357\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__39357\,
            I => \N__39354\
        );

    \I__7592\ : Odrv12
    port map (
            O => \N__39354\,
            I => \dron_frame_decoder_1.drone_H_disp_front_8\
        );

    \I__7591\ : IoInMux
    port map (
            O => \N__39351\,
            I => \N__39348\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__39348\,
            I => \N__39345\
        );

    \I__7589\ : Odrv4
    port map (
            O => \N__39345\,
            I => \pid_alt.state_0_0\
        );

    \I__7588\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39339\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__39339\,
            I => \drone_H_disp_front_i_6\
        );

    \I__7586\ : CascadeMux
    port map (
            O => \N__39336\,
            I => \N__39333\
        );

    \I__7585\ : InMux
    port map (
            O => \N__39333\,
            I => \N__39330\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__39330\,
            I => front_command_2
        );

    \I__7583\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39323\
        );

    \I__7582\ : InMux
    port map (
            O => \N__39326\,
            I => \N__39320\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__39323\,
            I => \N__39317\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__39320\,
            I => \N__39314\
        );

    \I__7579\ : Span4Mux_s3_h
    port map (
            O => \N__39317\,
            I => \N__39311\
        );

    \I__7578\ : Span12Mux_s1_h
    port map (
            O => \N__39314\,
            I => \N__39308\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__39311\,
            I => \N__39305\
        );

    \I__7576\ : Span12Mux_h
    port map (
            O => \N__39308\,
            I => \N__39302\
        );

    \I__7575\ : Span4Mux_h
    port map (
            O => \N__39305\,
            I => \N__39299\
        );

    \I__7574\ : Odrv12
    port map (
            O => \N__39302\,
            I => \pid_front.error_6\
        );

    \I__7573\ : Odrv4
    port map (
            O => \N__39299\,
            I => \pid_front.error_6\
        );

    \I__7572\ : InMux
    port map (
            O => \N__39294\,
            I => \pid_front.error_cry_1_0\
        );

    \I__7571\ : InMux
    port map (
            O => \N__39291\,
            I => \N__39288\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__39288\,
            I => \N__39285\
        );

    \I__7569\ : Span4Mux_v
    port map (
            O => \N__39285\,
            I => \N__39282\
        );

    \I__7568\ : Odrv4
    port map (
            O => \N__39282\,
            I => \drone_H_disp_front_i_7\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__39279\,
            I => \N__39276\
        );

    \I__7566\ : InMux
    port map (
            O => \N__39276\,
            I => \N__39273\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__39273\,
            I => front_command_3
        );

    \I__7564\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39267\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__39267\,
            I => \N__39263\
        );

    \I__7562\ : InMux
    port map (
            O => \N__39266\,
            I => \N__39260\
        );

    \I__7561\ : Span4Mux_v
    port map (
            O => \N__39263\,
            I => \N__39257\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__39260\,
            I => \N__39254\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__39257\,
            I => \N__39251\
        );

    \I__7558\ : Span4Mux_s3_h
    port map (
            O => \N__39254\,
            I => \N__39248\
        );

    \I__7557\ : Span4Mux_h
    port map (
            O => \N__39251\,
            I => \N__39245\
        );

    \I__7556\ : Span4Mux_h
    port map (
            O => \N__39248\,
            I => \N__39242\
        );

    \I__7555\ : Span4Mux_h
    port map (
            O => \N__39245\,
            I => \N__39239\
        );

    \I__7554\ : Span4Mux_h
    port map (
            O => \N__39242\,
            I => \N__39236\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__39239\,
            I => \pid_front.error_7\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__39236\,
            I => \pid_front.error_7\
        );

    \I__7551\ : InMux
    port map (
            O => \N__39231\,
            I => \pid_front.error_cry_2_0\
        );

    \I__7550\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39225\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__39225\,
            I => \N__39222\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__39222\,
            I => \drone_H_disp_front_i_8\
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__7546\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39213\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__39213\,
            I => front_command_4
        );

    \I__7544\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39207\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__39207\,
            I => \N__39203\
        );

    \I__7542\ : InMux
    port map (
            O => \N__39206\,
            I => \N__39200\
        );

    \I__7541\ : Span4Mux_v
    port map (
            O => \N__39203\,
            I => \N__39197\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__39200\,
            I => \N__39194\
        );

    \I__7539\ : Span4Mux_h
    port map (
            O => \N__39197\,
            I => \N__39191\
        );

    \I__7538\ : Span4Mux_s3_h
    port map (
            O => \N__39194\,
            I => \N__39188\
        );

    \I__7537\ : Span4Mux_h
    port map (
            O => \N__39191\,
            I => \N__39185\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__39188\,
            I => \N__39182\
        );

    \I__7535\ : Span4Mux_h
    port map (
            O => \N__39185\,
            I => \N__39179\
        );

    \I__7534\ : Span4Mux_h
    port map (
            O => \N__39182\,
            I => \N__39176\
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__39179\,
            I => \pid_front.error_8\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__39176\,
            I => \pid_front.error_8\
        );

    \I__7531\ : InMux
    port map (
            O => \N__39171\,
            I => \bfn_13_24_0_\
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__39168\,
            I => \N__39165\
        );

    \I__7529\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39162\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__39162\,
            I => front_command_5
        );

    \I__7527\ : InMux
    port map (
            O => \N__39159\,
            I => \N__39156\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__39156\,
            I => \N__39152\
        );

    \I__7525\ : InMux
    port map (
            O => \N__39155\,
            I => \N__39149\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__39152\,
            I => \N__39146\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__39149\,
            I => \N__39143\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__39146\,
            I => \N__39140\
        );

    \I__7521\ : Span4Mux_s3_h
    port map (
            O => \N__39143\,
            I => \N__39137\
        );

    \I__7520\ : Span4Mux_h
    port map (
            O => \N__39140\,
            I => \N__39134\
        );

    \I__7519\ : Span4Mux_h
    port map (
            O => \N__39137\,
            I => \N__39131\
        );

    \I__7518\ : Span4Mux_h
    port map (
            O => \N__39134\,
            I => \N__39128\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__39131\,
            I => \N__39125\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__39128\,
            I => \pid_front.error_9\
        );

    \I__7515\ : Odrv4
    port map (
            O => \N__39125\,
            I => \pid_front.error_9\
        );

    \I__7514\ : InMux
    port map (
            O => \N__39120\,
            I => \pid_front.error_cry_4\
        );

    \I__7513\ : InMux
    port map (
            O => \N__39117\,
            I => \N__39114\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__39114\,
            I => \drone_H_disp_front_i_10\
        );

    \I__7511\ : CascadeMux
    port map (
            O => \N__39111\,
            I => \N__39108\
        );

    \I__7510\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39105\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__39105\,
            I => \N__39102\
        );

    \I__7508\ : Odrv4
    port map (
            O => \N__39102\,
            I => front_command_6
        );

    \I__7507\ : InMux
    port map (
            O => \N__39099\,
            I => \N__39096\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__39096\,
            I => \N__39092\
        );

    \I__7505\ : InMux
    port map (
            O => \N__39095\,
            I => \N__39089\
        );

    \I__7504\ : Span4Mux_v
    port map (
            O => \N__39092\,
            I => \N__39086\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__39089\,
            I => \N__39083\
        );

    \I__7502\ : Span4Mux_h
    port map (
            O => \N__39086\,
            I => \N__39080\
        );

    \I__7501\ : Span4Mux_s3_h
    port map (
            O => \N__39083\,
            I => \N__39077\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__39080\,
            I => \N__39074\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__39077\,
            I => \N__39071\
        );

    \I__7498\ : Span4Mux_h
    port map (
            O => \N__39074\,
            I => \N__39068\
        );

    \I__7497\ : Span4Mux_h
    port map (
            O => \N__39071\,
            I => \N__39065\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__39068\,
            I => \pid_front.error_10\
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__39065\,
            I => \pid_front.error_10\
        );

    \I__7494\ : InMux
    port map (
            O => \N__39060\,
            I => \pid_front.error_cry_5\
        );

    \I__7493\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39054\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__39054\,
            I => \pid_front.error_axbZ0Z_7\
        );

    \I__7491\ : InMux
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__39048\,
            I => \N__39044\
        );

    \I__7489\ : InMux
    port map (
            O => \N__39047\,
            I => \N__39041\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__39044\,
            I => \N__39038\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__39041\,
            I => \N__39035\
        );

    \I__7486\ : Span4Mux_h
    port map (
            O => \N__39038\,
            I => \N__39032\
        );

    \I__7485\ : Span4Mux_s3_h
    port map (
            O => \N__39035\,
            I => \N__39029\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__39032\,
            I => \N__39026\
        );

    \I__7483\ : Span4Mux_h
    port map (
            O => \N__39029\,
            I => \N__39023\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__39026\,
            I => \N__39020\
        );

    \I__7481\ : Span4Mux_h
    port map (
            O => \N__39023\,
            I => \N__39017\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__39020\,
            I => \pid_front.error_11\
        );

    \I__7479\ : Odrv4
    port map (
            O => \N__39017\,
            I => \pid_front.error_11\
        );

    \I__7478\ : InMux
    port map (
            O => \N__39012\,
            I => \pid_front.error_cry_6\
        );

    \I__7477\ : InMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__39006\,
            I => \pid_front.error_axb_8_l_ofx_0\
        );

    \I__7475\ : InMux
    port map (
            O => \N__39003\,
            I => \N__39000\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__39000\,
            I => \N__38997\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__38997\,
            I => \N__38994\
        );

    \I__7472\ : Span4Mux_h
    port map (
            O => \N__38994\,
            I => \N__38990\
        );

    \I__7471\ : InMux
    port map (
            O => \N__38993\,
            I => \N__38987\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__38990\,
            I => \N__38984\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__38987\,
            I => \N__38981\
        );

    \I__7468\ : Span4Mux_h
    port map (
            O => \N__38984\,
            I => \N__38978\
        );

    \I__7467\ : Span12Mux_s6_v
    port map (
            O => \N__38981\,
            I => \N__38975\
        );

    \I__7466\ : Odrv4
    port map (
            O => \N__38978\,
            I => \pid_front.error_12\
        );

    \I__7465\ : Odrv12
    port map (
            O => \N__38975\,
            I => \pid_front.error_12\
        );

    \I__7464\ : InMux
    port map (
            O => \N__38970\,
            I => \pid_front.error_cry_7\
        );

    \I__7463\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38964\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__38964\,
            I => \drone_H_disp_front_i_12\
        );

    \I__7461\ : InMux
    port map (
            O => \N__38961\,
            I => \N__38957\
        );

    \I__7460\ : InMux
    port map (
            O => \N__38960\,
            I => \N__38954\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__38957\,
            I => \N__38951\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__38954\,
            I => \N__38948\
        );

    \I__7457\ : Span4Mux_v
    port map (
            O => \N__38951\,
            I => \N__38945\
        );

    \I__7456\ : Span12Mux_s1_h
    port map (
            O => \N__38948\,
            I => \N__38942\
        );

    \I__7455\ : Span4Mux_h
    port map (
            O => \N__38945\,
            I => \N__38939\
        );

    \I__7454\ : Span12Mux_h
    port map (
            O => \N__38942\,
            I => \N__38936\
        );

    \I__7453\ : Span4Mux_h
    port map (
            O => \N__38939\,
            I => \N__38933\
        );

    \I__7452\ : Odrv12
    port map (
            O => \N__38936\,
            I => \pid_front.error_13\
        );

    \I__7451\ : Odrv4
    port map (
            O => \N__38933\,
            I => \pid_front.error_13\
        );

    \I__7450\ : InMux
    port map (
            O => \N__38928\,
            I => \pid_front.error_cry_8\
        );

    \I__7449\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38922\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__38922\,
            I => \N__38919\
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__38919\,
            I => \drone_H_disp_front_2\
        );

    \I__7446\ : InMux
    port map (
            O => \N__38916\,
            I => \N__38913\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__38913\,
            I => \N__38909\
        );

    \I__7444\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38906\
        );

    \I__7443\ : Span4Mux_v
    port map (
            O => \N__38909\,
            I => \N__38903\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__38906\,
            I => \N__38899\
        );

    \I__7441\ : Span4Mux_h
    port map (
            O => \N__38903\,
            I => \N__38896\
        );

    \I__7440\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38893\
        );

    \I__7439\ : Span12Mux_v
    port map (
            O => \N__38899\,
            I => \N__38890\
        );

    \I__7438\ : Span4Mux_h
    port map (
            O => \N__38896\,
            I => \N__38887\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__38893\,
            I => \N__38884\
        );

    \I__7436\ : Span12Mux_h
    port map (
            O => \N__38890\,
            I => \N__38881\
        );

    \I__7435\ : Span4Mux_h
    port map (
            O => \N__38887\,
            I => \N__38876\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__38884\,
            I => \N__38876\
        );

    \I__7433\ : Odrv12
    port map (
            O => \N__38881\,
            I => \drone_H_disp_front_0\
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__38876\,
            I => \drone_H_disp_front_0\
        );

    \I__7431\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38868\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__38868\,
            I => \pid_front.error_axb_0\
        );

    \I__7429\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38862\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__38862\,
            I => \N__38859\
        );

    \I__7427\ : Span4Mux_v
    port map (
            O => \N__38859\,
            I => \N__38856\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__38856\,
            I => \pid_front.error_axbZ0Z_1\
        );

    \I__7425\ : InMux
    port map (
            O => \N__38853\,
            I => \N__38850\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__38850\,
            I => \N__38846\
        );

    \I__7423\ : InMux
    port map (
            O => \N__38849\,
            I => \N__38843\
        );

    \I__7422\ : Span4Mux_s1_h
    port map (
            O => \N__38846\,
            I => \N__38840\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__38843\,
            I => \N__38837\
        );

    \I__7420\ : Span4Mux_v
    port map (
            O => \N__38840\,
            I => \N__38834\
        );

    \I__7419\ : Span4Mux_s0_h
    port map (
            O => \N__38837\,
            I => \N__38831\
        );

    \I__7418\ : Span4Mux_h
    port map (
            O => \N__38834\,
            I => \N__38828\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__38831\,
            I => \N__38825\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__38828\,
            I => \N__38822\
        );

    \I__7415\ : Span4Mux_h
    port map (
            O => \N__38825\,
            I => \N__38819\
        );

    \I__7414\ : Span4Mux_h
    port map (
            O => \N__38822\,
            I => \N__38814\
        );

    \I__7413\ : Span4Mux_h
    port map (
            O => \N__38819\,
            I => \N__38814\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__38814\,
            I => \pid_front.error_1\
        );

    \I__7411\ : InMux
    port map (
            O => \N__38811\,
            I => \pid_front.error_cry_0\
        );

    \I__7410\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38805\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__38805\,
            I => \pid_front.error_axbZ0Z_2\
        );

    \I__7408\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38799\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38796\
        );

    \I__7406\ : Span4Mux_v
    port map (
            O => \N__38796\,
            I => \N__38792\
        );

    \I__7405\ : InMux
    port map (
            O => \N__38795\,
            I => \N__38789\
        );

    \I__7404\ : Span4Mux_v
    port map (
            O => \N__38792\,
            I => \N__38786\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__38789\,
            I => \N__38783\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__38786\,
            I => \N__38780\
        );

    \I__7401\ : Span4Mux_v
    port map (
            O => \N__38783\,
            I => \N__38777\
        );

    \I__7400\ : Span4Mux_h
    port map (
            O => \N__38780\,
            I => \N__38774\
        );

    \I__7399\ : Span4Mux_h
    port map (
            O => \N__38777\,
            I => \N__38771\
        );

    \I__7398\ : Span4Mux_h
    port map (
            O => \N__38774\,
            I => \N__38766\
        );

    \I__7397\ : Span4Mux_h
    port map (
            O => \N__38771\,
            I => \N__38766\
        );

    \I__7396\ : Odrv4
    port map (
            O => \N__38766\,
            I => \pid_front.error_2\
        );

    \I__7395\ : InMux
    port map (
            O => \N__38763\,
            I => \pid_front.error_cry_1\
        );

    \I__7394\ : InMux
    port map (
            O => \N__38760\,
            I => \N__38757\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__38757\,
            I => \N__38754\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__38754\,
            I => \pid_front.error_axbZ0Z_3\
        );

    \I__7391\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38748\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__38748\,
            I => \N__38744\
        );

    \I__7389\ : InMux
    port map (
            O => \N__38747\,
            I => \N__38741\
        );

    \I__7388\ : Span4Mux_v
    port map (
            O => \N__38744\,
            I => \N__38738\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__38741\,
            I => \N__38735\
        );

    \I__7386\ : Span4Mux_h
    port map (
            O => \N__38738\,
            I => \N__38732\
        );

    \I__7385\ : Span4Mux_v
    port map (
            O => \N__38735\,
            I => \N__38729\
        );

    \I__7384\ : Span4Mux_h
    port map (
            O => \N__38732\,
            I => \N__38726\
        );

    \I__7383\ : Span4Mux_h
    port map (
            O => \N__38729\,
            I => \N__38723\
        );

    \I__7382\ : Span4Mux_h
    port map (
            O => \N__38726\,
            I => \N__38720\
        );

    \I__7381\ : Span4Mux_h
    port map (
            O => \N__38723\,
            I => \N__38717\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__38720\,
            I => \pid_front.error_3\
        );

    \I__7379\ : Odrv4
    port map (
            O => \N__38717\,
            I => \pid_front.error_3\
        );

    \I__7378\ : InMux
    port map (
            O => \N__38712\,
            I => \pid_front.error_cry_2\
        );

    \I__7377\ : InMux
    port map (
            O => \N__38709\,
            I => \N__38706\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__38706\,
            I => \drone_H_disp_front_i_4\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__38703\,
            I => \N__38700\
        );

    \I__7374\ : InMux
    port map (
            O => \N__38700\,
            I => \N__38697\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__7372\ : Odrv4
    port map (
            O => \N__38694\,
            I => front_command_0
        );

    \I__7371\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38688\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__38688\,
            I => \N__38685\
        );

    \I__7369\ : Span4Mux_s2_h
    port map (
            O => \N__38685\,
            I => \N__38681\
        );

    \I__7368\ : InMux
    port map (
            O => \N__38684\,
            I => \N__38678\
        );

    \I__7367\ : Span4Mux_v
    port map (
            O => \N__38681\,
            I => \N__38675\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__38678\,
            I => \N__38672\
        );

    \I__7365\ : Span4Mux_h
    port map (
            O => \N__38675\,
            I => \N__38669\
        );

    \I__7364\ : Span4Mux_s3_h
    port map (
            O => \N__38672\,
            I => \N__38666\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__38669\,
            I => \N__38663\
        );

    \I__7362\ : Span4Mux_h
    port map (
            O => \N__38666\,
            I => \N__38660\
        );

    \I__7361\ : Span4Mux_h
    port map (
            O => \N__38663\,
            I => \N__38655\
        );

    \I__7360\ : Span4Mux_h
    port map (
            O => \N__38660\,
            I => \N__38655\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__38655\,
            I => \pid_front.error_4\
        );

    \I__7358\ : InMux
    port map (
            O => \N__38652\,
            I => \pid_front.error_cry_3\
        );

    \I__7357\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38646\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__38646\,
            I => \drone_H_disp_front_i_5\
        );

    \I__7355\ : CascadeMux
    port map (
            O => \N__38643\,
            I => \N__38640\
        );

    \I__7354\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38637\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__38637\,
            I => front_command_1
        );

    \I__7352\ : InMux
    port map (
            O => \N__38634\,
            I => \N__38631\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__38631\,
            I => \N__38627\
        );

    \I__7350\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38624\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__38627\,
            I => \N__38621\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__38624\,
            I => \N__38618\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__38621\,
            I => \N__38615\
        );

    \I__7346\ : Span4Mux_v
    port map (
            O => \N__38618\,
            I => \N__38612\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__38615\,
            I => \N__38609\
        );

    \I__7344\ : Span4Mux_h
    port map (
            O => \N__38612\,
            I => \N__38606\
        );

    \I__7343\ : Span4Mux_h
    port map (
            O => \N__38609\,
            I => \N__38603\
        );

    \I__7342\ : Span4Mux_h
    port map (
            O => \N__38606\,
            I => \N__38600\
        );

    \I__7341\ : Odrv4
    port map (
            O => \N__38603\,
            I => \pid_front.error_5\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__38600\,
            I => \pid_front.error_5\
        );

    \I__7339\ : InMux
    port map (
            O => \N__38595\,
            I => \pid_front.error_cry_0_0\
        );

    \I__7338\ : CascadeMux
    port map (
            O => \N__38592\,
            I => \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1_cascade_\
        );

    \I__7337\ : CascadeMux
    port map (
            O => \N__38589\,
            I => \N__38585\
        );

    \I__7336\ : InMux
    port map (
            O => \N__38588\,
            I => \N__38582\
        );

    \I__7335\ : InMux
    port map (
            O => \N__38585\,
            I => \N__38579\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__38582\,
            I => \pid_front.un1_pid_prereg\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__38579\,
            I => \pid_front.un1_pid_prereg\
        );

    \I__7332\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38571\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__38571\,
            I => \drone_H_disp_front_3\
        );

    \I__7330\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38565\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__38565\,
            I => \N__38561\
        );

    \I__7328\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38558\
        );

    \I__7327\ : Odrv4
    port map (
            O => \N__38561\,
            I => \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__38558\,
            I => \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1\
        );

    \I__7325\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38546\
        );

    \I__7324\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38546\
        );

    \I__7323\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38543\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__38546\,
            I => \N__38540\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__38543\,
            I => \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__38540\,
            I => \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2\
        );

    \I__7319\ : InMux
    port map (
            O => \N__38535\,
            I => \N__38532\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__38532\,
            I => \pid_front.error_p_reg_esr_RNIUQTFZ0Z_1\
        );

    \I__7317\ : InMux
    port map (
            O => \N__38529\,
            I => \N__38524\
        );

    \I__7316\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38521\
        );

    \I__7315\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38518\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__38524\,
            I => \N__38515\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__38521\,
            I => \N__38512\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__38518\,
            I => \N__38507\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__38515\,
            I => \N__38507\
        );

    \I__7310\ : Span12Mux_v
    port map (
            O => \N__38512\,
            I => \N__38504\
        );

    \I__7309\ : Span4Mux_v
    port map (
            O => \N__38507\,
            I => \N__38501\
        );

    \I__7308\ : Span12Mux_h
    port map (
            O => \N__38504\,
            I => \N__38498\
        );

    \I__7307\ : Span4Mux_v
    port map (
            O => \N__38501\,
            I => \N__38495\
        );

    \I__7306\ : Odrv12
    port map (
            O => \N__38498\,
            I => \pid_alt.error_d_regZ0Z_15\
        );

    \I__7305\ : Odrv4
    port map (
            O => \N__38495\,
            I => \pid_alt.error_d_regZ0Z_15\
        );

    \I__7304\ : InMux
    port map (
            O => \N__38490\,
            I => \N__38487\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__38487\,
            I => \N__38483\
        );

    \I__7302\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38480\
        );

    \I__7301\ : Span4Mux_v
    port map (
            O => \N__38483\,
            I => \N__38477\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__38480\,
            I => \N__38474\
        );

    \I__7299\ : Span4Mux_h
    port map (
            O => \N__38477\,
            I => \N__38471\
        );

    \I__7298\ : Span4Mux_v
    port map (
            O => \N__38474\,
            I => \N__38468\
        );

    \I__7297\ : Span4Mux_h
    port map (
            O => \N__38471\,
            I => \N__38465\
        );

    \I__7296\ : Span4Mux_v
    port map (
            O => \N__38468\,
            I => \N__38462\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__38465\,
            I => \pid_alt.error_p_regZ0Z_15\
        );

    \I__7294\ : Odrv4
    port map (
            O => \N__38462\,
            I => \pid_alt.error_p_regZ0Z_15\
        );

    \I__7293\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38454\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__38454\,
            I => \N__38450\
        );

    \I__7291\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38447\
        );

    \I__7290\ : Span12Mux_h
    port map (
            O => \N__38450\,
            I => \N__38444\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__38447\,
            I => \N__38441\
        );

    \I__7288\ : Span12Mux_v
    port map (
            O => \N__38444\,
            I => \N__38438\
        );

    \I__7287\ : Span4Mux_v
    port map (
            O => \N__38441\,
            I => \N__38435\
        );

    \I__7286\ : Odrv12
    port map (
            O => \N__38438\,
            I => \pid_alt.error_d_reg_prevZ0Z_15\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__38435\,
            I => \pid_alt.error_d_reg_prevZ0Z_15\
        );

    \I__7284\ : InMux
    port map (
            O => \N__38430\,
            I => \N__38424\
        );

    \I__7283\ : InMux
    port map (
            O => \N__38429\,
            I => \N__38424\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__7281\ : Span12Mux_h
    port map (
            O => \N__38421\,
            I => \N__38418\
        );

    \I__7280\ : Odrv12
    port map (
            O => \N__38418\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\
        );

    \I__7279\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38412\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__38412\,
            I => \N__38409\
        );

    \I__7277\ : Odrv4
    port map (
            O => \N__38409\,
            I => \dron_frame_decoder_1.drone_H_disp_front_5\
        );

    \I__7276\ : InMux
    port map (
            O => \N__38406\,
            I => \N__38403\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__38403\,
            I => \N__38400\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__38400\,
            I => \dron_frame_decoder_1.drone_H_disp_front_4\
        );

    \I__7273\ : InMux
    port map (
            O => \N__38397\,
            I => \N__38393\
        );

    \I__7272\ : InMux
    port map (
            O => \N__38396\,
            I => \N__38390\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__38393\,
            I => \N__38387\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__38390\,
            I => \N__38383\
        );

    \I__7269\ : Span4Mux_h
    port map (
            O => \N__38387\,
            I => \N__38380\
        );

    \I__7268\ : InMux
    port map (
            O => \N__38386\,
            I => \N__38377\
        );

    \I__7267\ : Span4Mux_h
    port map (
            O => \N__38383\,
            I => \N__38374\
        );

    \I__7266\ : Span4Mux_h
    port map (
            O => \N__38380\,
            I => \N__38371\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__38377\,
            I => \N__38368\
        );

    \I__7264\ : Span4Mux_h
    port map (
            O => \N__38374\,
            I => \N__38365\
        );

    \I__7263\ : Span4Mux_v
    port map (
            O => \N__38371\,
            I => \N__38362\
        );

    \I__7262\ : Span4Mux_h
    port map (
            O => \N__38368\,
            I => \N__38357\
        );

    \I__7261\ : Span4Mux_v
    port map (
            O => \N__38365\,
            I => \N__38357\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__38362\,
            I => \pid_front.error_p_regZ0Z_0\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__38357\,
            I => \pid_front.error_p_regZ0Z_0\
        );

    \I__7258\ : InMux
    port map (
            O => \N__38352\,
            I => \N__38349\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__38349\,
            I => \N__38344\
        );

    \I__7256\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38341\
        );

    \I__7255\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38338\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__38344\,
            I => \N__38335\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__38341\,
            I => \N__38332\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__38338\,
            I => \pid_front.error_d_reg_prevZ0Z_0\
        );

    \I__7251\ : Odrv4
    port map (
            O => \N__38335\,
            I => \pid_front.error_d_reg_prevZ0Z_0\
        );

    \I__7250\ : Odrv4
    port map (
            O => \N__38332\,
            I => \pid_front.error_d_reg_prevZ0Z_0\
        );

    \I__7249\ : InMux
    port map (
            O => \N__38325\,
            I => \N__38321\
        );

    \I__7248\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38318\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__38321\,
            I => \pid_front.N_1427_i\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__38318\,
            I => \pid_front.N_1427_i\
        );

    \I__7245\ : InMux
    port map (
            O => \N__38313\,
            I => \N__38310\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__38310\,
            I => \N__38307\
        );

    \I__7243\ : Odrv4
    port map (
            O => \N__38307\,
            I => \dron_frame_decoder_1.drone_H_disp_front_6\
        );

    \I__7242\ : InMux
    port map (
            O => \N__38304\,
            I => \N__38298\
        );

    \I__7241\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38298\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__38298\,
            I => \N__38295\
        );

    \I__7239\ : Span4Mux_v
    port map (
            O => \N__38295\,
            I => \N__38290\
        );

    \I__7238\ : InMux
    port map (
            O => \N__38294\,
            I => \N__38285\
        );

    \I__7237\ : InMux
    port map (
            O => \N__38293\,
            I => \N__38285\
        );

    \I__7236\ : Odrv4
    port map (
            O => \N__38290\,
            I => \pid_front.error_d_reg_prevZ0Z_5\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__38285\,
            I => \pid_front.error_d_reg_prevZ0Z_5\
        );

    \I__7234\ : InMux
    port map (
            O => \N__38280\,
            I => \N__38274\
        );

    \I__7233\ : InMux
    port map (
            O => \N__38279\,
            I => \N__38274\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__38274\,
            I => \N__38271\
        );

    \I__7231\ : Span4Mux_h
    port map (
            O => \N__38271\,
            I => \N__38268\
        );

    \I__7230\ : Span4Mux_h
    port map (
            O => \N__38268\,
            I => \N__38265\
        );

    \I__7229\ : Span4Mux_h
    port map (
            O => \N__38265\,
            I => \N__38262\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__38262\,
            I => \pid_front.error_p_regZ0Z_4\
        );

    \I__7227\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38253\
        );

    \I__7226\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38253\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__38253\,
            I => \pid_front.error_d_reg_prevZ0Z_4\
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__38250\,
            I => \N__38247\
        );

    \I__7223\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38243\
        );

    \I__7222\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38240\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__38243\,
            I => \pid_front.un1_pid_prereg_17\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__38240\,
            I => \pid_front.un1_pid_prereg_17\
        );

    \I__7219\ : CascadeMux
    port map (
            O => \N__38235\,
            I => \pid_front.un1_pid_prereg_17_cascade_\
        );

    \I__7218\ : InMux
    port map (
            O => \N__38232\,
            I => \N__38225\
        );

    \I__7217\ : InMux
    port map (
            O => \N__38231\,
            I => \N__38225\
        );

    \I__7216\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38222\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__38225\,
            I => \pid_front.un1_pid_prereg_3\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__38222\,
            I => \pid_front.un1_pid_prereg_3\
        );

    \I__7213\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38214\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__38214\,
            I => \pid_front.error_p_reg_esr_RNIPISGZ0Z_3\
        );

    \I__7211\ : CascadeMux
    port map (
            O => \N__38211\,
            I => \pid_front.error_p_reg_esr_RNI4KF7Z0Z_0_cascade_\
        );

    \I__7210\ : InMux
    port map (
            O => \N__38208\,
            I => \N__38205\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__38205\,
            I => \pid_front.error_d_reg_esr_RNINGRVZ0Z_1\
        );

    \I__7208\ : InMux
    port map (
            O => \N__38202\,
            I => \N__38196\
        );

    \I__7207\ : InMux
    port map (
            O => \N__38201\,
            I => \N__38196\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__38196\,
            I => \N__38193\
        );

    \I__7205\ : Span12Mux_v
    port map (
            O => \N__38193\,
            I => \N__38190\
        );

    \I__7204\ : Odrv12
    port map (
            O => \N__38190\,
            I => \pid_front.error_p_regZ0Z_1\
        );

    \I__7203\ : InMux
    port map (
            O => \N__38187\,
            I => \N__38184\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__38184\,
            I => \ppm_encoder_1.un2_throttle_iv_1_13\
        );

    \I__7201\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38178\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__38178\,
            I => \ppm_encoder_1.N_299\
        );

    \I__7199\ : CascadeMux
    port map (
            O => \N__38175\,
            I => \N__38172\
        );

    \I__7198\ : InMux
    port map (
            O => \N__38172\,
            I => \N__38167\
        );

    \I__7197\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38162\
        );

    \I__7196\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38162\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__38167\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__38162\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__7193\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38154\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__38154\,
            I => \N__38150\
        );

    \I__7191\ : InMux
    port map (
            O => \N__38153\,
            I => \N__38147\
        );

    \I__7190\ : Span4Mux_h
    port map (
            O => \N__38150\,
            I => \N__38144\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__38147\,
            I => \N__38141\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__38144\,
            I => \N__38138\
        );

    \I__7187\ : Span12Mux_h
    port map (
            O => \N__38141\,
            I => \N__38135\
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__38138\,
            I => front_order_13
        );

    \I__7185\ : Odrv12
    port map (
            O => \N__38135\,
            I => front_order_13
        );

    \I__7184\ : InMux
    port map (
            O => \N__38130\,
            I => \N__38127\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__38127\,
            I => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\
        );

    \I__7182\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38119\
        );

    \I__7181\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38114\
        );

    \I__7180\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38114\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__38119\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__38114\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__7177\ : InMux
    port map (
            O => \N__38109\,
            I => \N__38106\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__38106\,
            I => \dron_frame_decoder_1.drone_H_disp_front_7\
        );

    \I__7175\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38099\
        );

    \I__7174\ : InMux
    port map (
            O => \N__38102\,
            I => \N__38096\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__38099\,
            I => \N__38091\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__38096\,
            I => \N__38091\
        );

    \I__7171\ : Span4Mux_h
    port map (
            O => \N__38091\,
            I => \N__38088\
        );

    \I__7170\ : Span4Mux_v
    port map (
            O => \N__38088\,
            I => \N__38085\
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__38085\,
            I => \pid_front.error_p_regZ0Z_2\
        );

    \I__7168\ : InMux
    port map (
            O => \N__38082\,
            I => \N__38078\
        );

    \I__7167\ : InMux
    port map (
            O => \N__38081\,
            I => \N__38075\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__38078\,
            I => \pid_front.error_d_reg_prevZ0Z_2\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__38075\,
            I => \pid_front.error_d_reg_prevZ0Z_2\
        );

    \I__7164\ : CascadeMux
    port map (
            O => \N__38070\,
            I => \N__38067\
        );

    \I__7163\ : InMux
    port map (
            O => \N__38067\,
            I => \N__38064\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__38064\,
            I => \pid_front.error_d_reg_esr_RNIOBP11Z0Z_5\
        );

    \I__7161\ : InMux
    port map (
            O => \N__38061\,
            I => \N__38058\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__38058\,
            I => \pid_front.un1_pid_prereg_40_0\
        );

    \I__7159\ : InMux
    port map (
            O => \N__38055\,
            I => \N__38052\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__38052\,
            I => \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4\
        );

    \I__7157\ : InMux
    port map (
            O => \N__38049\,
            I => \N__38041\
        );

    \I__7156\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38041\
        );

    \I__7155\ : InMux
    port map (
            O => \N__38047\,
            I => \N__38036\
        );

    \I__7154\ : InMux
    port map (
            O => \N__38046\,
            I => \N__38036\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__38041\,
            I => \N__38033\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__38036\,
            I => \N__38030\
        );

    \I__7151\ : Span4Mux_v
    port map (
            O => \N__38033\,
            I => \N__38025\
        );

    \I__7150\ : Span4Mux_h
    port map (
            O => \N__38030\,
            I => \N__38025\
        );

    \I__7149\ : Span4Mux_h
    port map (
            O => \N__38025\,
            I => \N__38022\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__38022\,
            I => \N__38019\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__38019\,
            I => \pid_front.error_p_regZ0Z_5\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__38016\,
            I => \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_\
        );

    \I__7145\ : InMux
    port map (
            O => \N__38013\,
            I => \N__38010\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__38010\,
            I => \N__38007\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__38007\,
            I => \N__38003\
        );

    \I__7142\ : InMux
    port map (
            O => \N__38006\,
            I => \N__38000\
        );

    \I__7141\ : Odrv4
    port map (
            O => \N__38003\,
            I => \pid_front.error_d_reg_esr_RNIVOSGZ0Z_5\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__38000\,
            I => \pid_front.error_d_reg_esr_RNIVOSGZ0Z_5\
        );

    \I__7139\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37990\
        );

    \I__7138\ : InMux
    port map (
            O => \N__37994\,
            I => \N__37987\
        );

    \I__7137\ : CascadeMux
    port map (
            O => \N__37993\,
            I => \N__37984\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__37990\,
            I => \N__37979\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__37987\,
            I => \N__37979\
        );

    \I__7134\ : InMux
    port map (
            O => \N__37984\,
            I => \N__37976\
        );

    \I__7133\ : Span4Mux_h
    port map (
            O => \N__37979\,
            I => \N__37973\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__37976\,
            I => front_order_8
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__37973\,
            I => front_order_8
        );

    \I__7130\ : InMux
    port map (
            O => \N__37968\,
            I => \N__37965\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__37965\,
            I => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\
        );

    \I__7128\ : InMux
    port map (
            O => \N__37962\,
            I => \bfn_13_17_0_\
        );

    \I__7127\ : InMux
    port map (
            O => \N__37959\,
            I => \N__37956\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__37956\,
            I => \N__37951\
        );

    \I__7125\ : InMux
    port map (
            O => \N__37955\,
            I => \N__37948\
        );

    \I__7124\ : CascadeMux
    port map (
            O => \N__37954\,
            I => \N__37945\
        );

    \I__7123\ : Span4Mux_v
    port map (
            O => \N__37951\,
            I => \N__37940\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__37948\,
            I => \N__37940\
        );

    \I__7121\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37937\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__37940\,
            I => \N__37934\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__37937\,
            I => front_order_9
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__37934\,
            I => front_order_9
        );

    \I__7117\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37926\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__37926\,
            I => \N__37923\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__37923\,
            I => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\
        );

    \I__7114\ : InMux
    port map (
            O => \N__37920\,
            I => \ppm_encoder_1.un1_elevator_cry_8\
        );

    \I__7113\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37912\
        );

    \I__7112\ : InMux
    port map (
            O => \N__37916\,
            I => \N__37909\
        );

    \I__7111\ : CascadeMux
    port map (
            O => \N__37915\,
            I => \N__37906\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__37912\,
            I => \N__37903\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__37909\,
            I => \N__37900\
        );

    \I__7108\ : InMux
    port map (
            O => \N__37906\,
            I => \N__37897\
        );

    \I__7107\ : Span4Mux_v
    port map (
            O => \N__37903\,
            I => \N__37894\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__37900\,
            I => \N__37891\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__37897\,
            I => front_order_10
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__37894\,
            I => front_order_10
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__37891\,
            I => front_order_10
        );

    \I__7102\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37881\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__37881\,
            I => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\
        );

    \I__7100\ : InMux
    port map (
            O => \N__37878\,
            I => \ppm_encoder_1.un1_elevator_cry_9\
        );

    \I__7099\ : InMux
    port map (
            O => \N__37875\,
            I => \N__37870\
        );

    \I__7098\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37867\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__37873\,
            I => \N__37864\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__37870\,
            I => \N__37861\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__37867\,
            I => \N__37858\
        );

    \I__7094\ : InMux
    port map (
            O => \N__37864\,
            I => \N__37855\
        );

    \I__7093\ : Span4Mux_h
    port map (
            O => \N__37861\,
            I => \N__37852\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__37858\,
            I => \N__37849\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__37855\,
            I => front_order_11
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__37852\,
            I => front_order_11
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__37849\,
            I => front_order_11
        );

    \I__7088\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37839\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__37839\,
            I => \N__37836\
        );

    \I__7086\ : Odrv4
    port map (
            O => \N__37836\,
            I => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\
        );

    \I__7085\ : InMux
    port map (
            O => \N__37833\,
            I => \ppm_encoder_1.un1_elevator_cry_10\
        );

    \I__7084\ : InMux
    port map (
            O => \N__37830\,
            I => \ppm_encoder_1.un1_elevator_cry_11\
        );

    \I__7083\ : InMux
    port map (
            O => \N__37827\,
            I => \ppm_encoder_1.un1_elevator_cry_12\
        );

    \I__7082\ : InMux
    port map (
            O => \N__37824\,
            I => \ppm_encoder_1.un1_elevator_cry_13\
        );

    \I__7081\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37817\
        );

    \I__7080\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37814\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__37817\,
            I => \N__37808\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37808\
        );

    \I__7077\ : InMux
    port map (
            O => \N__37813\,
            I => \N__37805\
        );

    \I__7076\ : Span4Mux_h
    port map (
            O => \N__37808\,
            I => \N__37802\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__37805\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__37802\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__37797\,
            I => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\
        );

    \I__7072\ : InMux
    port map (
            O => \N__37794\,
            I => \ppm_encoder_1.un1_elevator_cry_0\
        );

    \I__7071\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37787\
        );

    \I__7070\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37784\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__37787\,
            I => \N__37779\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__37784\,
            I => \N__37779\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__37779\,
            I => \N__37776\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__37776\,
            I => front_order_2
        );

    \I__7065\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37770\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__37770\,
            I => \ppm_encoder_1.un1_elevator_cry_1_THRU_CO\
        );

    \I__7063\ : InMux
    port map (
            O => \N__37767\,
            I => \ppm_encoder_1.un1_elevator_cry_1\
        );

    \I__7062\ : InMux
    port map (
            O => \N__37764\,
            I => \ppm_encoder_1.un1_elevator_cry_2\
        );

    \I__7061\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37757\
        );

    \I__7060\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37754\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37751\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__37754\,
            I => \N__37748\
        );

    \I__7057\ : Span4Mux_v
    port map (
            O => \N__37751\,
            I => \N__37743\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__37748\,
            I => \N__37743\
        );

    \I__7055\ : Span4Mux_v
    port map (
            O => \N__37743\,
            I => \N__37740\
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__37740\,
            I => front_order_4
        );

    \I__7053\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37734\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__37734\,
            I => \ppm_encoder_1.un1_elevator_cry_3_THRU_CO\
        );

    \I__7051\ : InMux
    port map (
            O => \N__37731\,
            I => \ppm_encoder_1.un1_elevator_cry_3\
        );

    \I__7050\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37724\
        );

    \I__7049\ : InMux
    port map (
            O => \N__37727\,
            I => \N__37721\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__37724\,
            I => \N__37718\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__37721\,
            I => \N__37715\
        );

    \I__7046\ : Span4Mux_h
    port map (
            O => \N__37718\,
            I => \N__37712\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__37715\,
            I => \N__37709\
        );

    \I__7044\ : Span4Mux_v
    port map (
            O => \N__37712\,
            I => \N__37706\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__37709\,
            I => \N__37703\
        );

    \I__7042\ : Odrv4
    port map (
            O => \N__37706\,
            I => front_order_5
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__37703\,
            I => front_order_5
        );

    \I__7040\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37695\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__37695\,
            I => \ppm_encoder_1.un1_elevator_cry_4_THRU_CO\
        );

    \I__7038\ : InMux
    port map (
            O => \N__37692\,
            I => \ppm_encoder_1.un1_elevator_cry_4\
        );

    \I__7037\ : InMux
    port map (
            O => \N__37689\,
            I => \N__37685\
        );

    \I__7036\ : CascadeMux
    port map (
            O => \N__37688\,
            I => \N__37682\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__37685\,
            I => \N__37678\
        );

    \I__7034\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37675\
        );

    \I__7033\ : CascadeMux
    port map (
            O => \N__37681\,
            I => \N__37672\
        );

    \I__7032\ : Span4Mux_v
    port map (
            O => \N__37678\,
            I => \N__37667\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__37675\,
            I => \N__37667\
        );

    \I__7030\ : InMux
    port map (
            O => \N__37672\,
            I => \N__37664\
        );

    \I__7029\ : Span4Mux_h
    port map (
            O => \N__37667\,
            I => \N__37661\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__37664\,
            I => front_order_6
        );

    \I__7027\ : Odrv4
    port map (
            O => \N__37661\,
            I => front_order_6
        );

    \I__7026\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37653\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__37653\,
            I => \ppm_encoder_1.un1_elevator_cry_5_THRU_CO\
        );

    \I__7024\ : InMux
    port map (
            O => \N__37650\,
            I => \ppm_encoder_1.un1_elevator_cry_5\
        );

    \I__7023\ : InMux
    port map (
            O => \N__37647\,
            I => \ppm_encoder_1.un1_elevator_cry_6\
        );

    \I__7022\ : CascadeMux
    port map (
            O => \N__37644\,
            I => \ppm_encoder_1.N_134_0_cascade_\
        );

    \I__7021\ : IoInMux
    port map (
            O => \N__37641\,
            I => \N__37638\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__37638\,
            I => \N__37635\
        );

    \I__7019\ : Span12Mux_s11_v
    port map (
            O => \N__37635\,
            I => \N__37631\
        );

    \I__7018\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37628\
        );

    \I__7017\ : Odrv12
    port map (
            O => \N__37631\,
            I => ppm_output_c
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__37628\,
            I => ppm_output_c
        );

    \I__7015\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37617\
        );

    \I__7013\ : Odrv12
    port map (
            O => \N__37617\,
            I => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\
        );

    \I__7012\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37610\
        );

    \I__7011\ : InMux
    port map (
            O => \N__37613\,
            I => \N__37607\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__37610\,
            I => \N__37602\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__37607\,
            I => \N__37602\
        );

    \I__7008\ : Span12Mux_h
    port map (
            O => \N__37602\,
            I => \N__37599\
        );

    \I__7007\ : Odrv12
    port map (
            O => \N__37599\,
            I => throttle_order_2
        );

    \I__7006\ : InMux
    port map (
            O => \N__37596\,
            I => \N__37592\
        );

    \I__7005\ : InMux
    port map (
            O => \N__37595\,
            I => \N__37589\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__37592\,
            I => \N__37586\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__37589\,
            I => \N__37583\
        );

    \I__7002\ : Odrv12
    port map (
            O => \N__37586\,
            I => scaler_4_data_6
        );

    \I__7001\ : Odrv4
    port map (
            O => \N__37583\,
            I => scaler_4_data_6
        );

    \I__7000\ : InMux
    port map (
            O => \N__37578\,
            I => \N__37575\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__37575\,
            I => \N__37572\
        );

    \I__6998\ : Span4Mux_h
    port map (
            O => \N__37572\,
            I => \N__37569\
        );

    \I__6997\ : Span4Mux_h
    port map (
            O => \N__37569\,
            I => \N__37566\
        );

    \I__6996\ : Odrv4
    port map (
            O => \N__37566\,
            I => \ppm_encoder_1.un1_aileron_cry_4_THRU_CO\
        );

    \I__6995\ : CascadeMux
    port map (
            O => \N__37563\,
            I => \N__37560\
        );

    \I__6994\ : InMux
    port map (
            O => \N__37560\,
            I => \N__37554\
        );

    \I__6993\ : InMux
    port map (
            O => \N__37559\,
            I => \N__37554\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__37554\,
            I => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\
        );

    \I__6991\ : InMux
    port map (
            O => \N__37551\,
            I => \scaler_4.un2_source_data_0_cry_4\
        );

    \I__6990\ : CascadeMux
    port map (
            O => \N__37548\,
            I => \N__37545\
        );

    \I__6989\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37539\
        );

    \I__6988\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37539\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__37539\,
            I => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\
        );

    \I__6986\ : InMux
    port map (
            O => \N__37536\,
            I => \scaler_4.un2_source_data_0_cry_5\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__37533\,
            I => \N__37530\
        );

    \I__6984\ : InMux
    port map (
            O => \N__37530\,
            I => \N__37524\
        );

    \I__6983\ : InMux
    port map (
            O => \N__37529\,
            I => \N__37524\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__37524\,
            I => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\
        );

    \I__6981\ : InMux
    port map (
            O => \N__37521\,
            I => \scaler_4.un2_source_data_0_cry_6\
        );

    \I__6980\ : CascadeMux
    port map (
            O => \N__37518\,
            I => \N__37515\
        );

    \I__6979\ : InMux
    port map (
            O => \N__37515\,
            I => \N__37509\
        );

    \I__6978\ : InMux
    port map (
            O => \N__37514\,
            I => \N__37509\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__37509\,
            I => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\
        );

    \I__6976\ : InMux
    port map (
            O => \N__37506\,
            I => \scaler_4.un2_source_data_0_cry_7\
        );

    \I__6975\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37499\
        );

    \I__6974\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37496\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__37499\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__37496\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__6971\ : CascadeMux
    port map (
            O => \N__37491\,
            I => \N__37488\
        );

    \I__6970\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37485\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__37485\,
            I => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\
        );

    \I__6968\ : InMux
    port map (
            O => \N__37482\,
            I => \bfn_13_13_0_\
        );

    \I__6967\ : InMux
    port map (
            O => \N__37479\,
            I => \scaler_4.un2_source_data_0_cry_9\
        );

    \I__6966\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37473\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37470\
        );

    \I__6964\ : Odrv4
    port map (
            O => \N__37470\,
            I => scaler_4_data_14
        );

    \I__6963\ : CEMux
    port map (
            O => \N__37467\,
            I => \N__37463\
        );

    \I__6962\ : CEMux
    port map (
            O => \N__37466\,
            I => \N__37460\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__37463\,
            I => \N__37457\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__37460\,
            I => \N__37454\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__37457\,
            I => \N__37448\
        );

    \I__6958\ : Span4Mux_v
    port map (
            O => \N__37454\,
            I => \N__37448\
        );

    \I__6957\ : CEMux
    port map (
            O => \N__37453\,
            I => \N__37445\
        );

    \I__6956\ : Sp12to4
    port map (
            O => \N__37448\,
            I => \N__37440\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__37445\,
            I => \N__37440\
        );

    \I__6954\ : Odrv12
    port map (
            O => \N__37440\,
            I => \scaler_4.debug_CH3_20A_c_0\
        );

    \I__6953\ : InMux
    port map (
            O => \N__37437\,
            I => \N__37434\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37431\
        );

    \I__6951\ : Odrv12
    port map (
            O => \N__37431\,
            I => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\
        );

    \I__6950\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37424\
        );

    \I__6949\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37421\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37418\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__37421\,
            I => \N__37415\
        );

    \I__6946\ : Odrv4
    port map (
            O => \N__37418\,
            I => scaler_4_data_7
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__37415\,
            I => scaler_4_data_7
        );

    \I__6944\ : InMux
    port map (
            O => \N__37410\,
            I => \ppm_encoder_1.un1_rudder_cry_9\
        );

    \I__6943\ : InMux
    port map (
            O => \N__37407\,
            I => \ppm_encoder_1.un1_rudder_cry_10\
        );

    \I__6942\ : InMux
    port map (
            O => \N__37404\,
            I => \ppm_encoder_1.un1_rudder_cry_11\
        );

    \I__6941\ : InMux
    port map (
            O => \N__37401\,
            I => \ppm_encoder_1.un1_rudder_cry_12\
        );

    \I__6940\ : InMux
    port map (
            O => \N__37398\,
            I => \bfn_13_11_0_\
        );

    \I__6939\ : InMux
    port map (
            O => \N__37395\,
            I => \scaler_4.un2_source_data_0_cry_1\
        );

    \I__6938\ : CascadeMux
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__6937\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37383\
        );

    \I__6936\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37383\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__37383\,
            I => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\
        );

    \I__6934\ : InMux
    port map (
            O => \N__37380\,
            I => \scaler_4.un2_source_data_0_cry_2\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__6932\ : InMux
    port map (
            O => \N__37374\,
            I => \N__37368\
        );

    \I__6931\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37368\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__37368\,
            I => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\
        );

    \I__6929\ : InMux
    port map (
            O => \N__37365\,
            I => \scaler_4.un2_source_data_0_cry_3\
        );

    \I__6928\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37356\
        );

    \I__6927\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37356\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__37356\,
            I => \N__37353\
        );

    \I__6925\ : Span12Mux_h
    port map (
            O => \N__37353\,
            I => \N__37350\
        );

    \I__6924\ : Odrv12
    port map (
            O => \N__37350\,
            I => \pid_front.error_p_regZ0Z_20\
        );

    \I__6923\ : InMux
    port map (
            O => \N__37347\,
            I => \ppm_encoder_1.un1_rudder_cry_6\
        );

    \I__6922\ : InMux
    port map (
            O => \N__37344\,
            I => \ppm_encoder_1.un1_rudder_cry_7\
        );

    \I__6921\ : InMux
    port map (
            O => \N__37341\,
            I => \ppm_encoder_1.un1_rudder_cry_8\
        );

    \I__6920\ : CEMux
    port map (
            O => \N__37338\,
            I => \N__37335\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__37335\,
            I => \N__37332\
        );

    \I__6918\ : Span4Mux_h
    port map (
            O => \N__37332\,
            I => \N__37329\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__37329\,
            I => \N__37326\
        );

    \I__6916\ : Sp12to4
    port map (
            O => \N__37326\,
            I => \N__37323\
        );

    \I__6915\ : Odrv12
    port map (
            O => \N__37323\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6914\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37317\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37314\
        );

    \I__6912\ : Odrv4
    port map (
            O => \N__37314\,
            I => \pid_front.un1_pid_prereg_axb_21\
        );

    \I__6911\ : CascadeMux
    port map (
            O => \N__37311\,
            I => \N__37308\
        );

    \I__6910\ : InMux
    port map (
            O => \N__37308\,
            I => \N__37302\
        );

    \I__6909\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37302\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__37302\,
            I => front_command_7
        );

    \I__6907\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37296\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__37296\,
            I => \N__37293\
        );

    \I__6905\ : Odrv4
    port map (
            O => \N__37293\,
            I => \pid_front.error_p_reg_esr_RNIHGOC2Z0Z_16\
        );

    \I__6904\ : CascadeMux
    port map (
            O => \N__37290\,
            I => \N__37287\
        );

    \I__6903\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37284\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__37284\,
            I => \N__37281\
        );

    \I__6901\ : Odrv4
    port map (
            O => \N__37281\,
            I => \pid_front.error_p_reg_esr_RNI87HP4Z0Z_16\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__37278\,
            I => \N__37275\
        );

    \I__6899\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37272\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__37272\,
            I => \pid_front.pid_preregZ0Z_18\
        );

    \I__6897\ : InMux
    port map (
            O => \N__37269\,
            I => \pid_front.un1_pid_prereg_cry_15\
        );

    \I__6896\ : InMux
    port map (
            O => \N__37266\,
            I => \N__37263\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__37263\,
            I => \N__37260\
        );

    \I__6894\ : Odrv4
    port map (
            O => \N__37260\,
            I => \pid_front.error_p_reg_esr_RNINMOC2Z0Z_17\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__37257\,
            I => \N__37254\
        );

    \I__6892\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37251\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__37251\,
            I => \N__37248\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__37248\,
            I => \pid_front.error_p_reg_esr_RNIKJHP4Z0Z_17\
        );

    \I__6889\ : InMux
    port map (
            O => \N__37245\,
            I => \N__37242\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__37242\,
            I => \pid_front.pid_preregZ0Z_19\
        );

    \I__6887\ : InMux
    port map (
            O => \N__37239\,
            I => \pid_front.un1_pid_prereg_cry_16\
        );

    \I__6886\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37233\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__37233\,
            I => \N__37230\
        );

    \I__6884\ : Odrv12
    port map (
            O => \N__37230\,
            I => \pid_front.error_p_reg_esr_RNITSOC2Z0Z_18\
        );

    \I__6883\ : CascadeMux
    port map (
            O => \N__37227\,
            I => \N__37224\
        );

    \I__6882\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37221\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__37221\,
            I => \N__37218\
        );

    \I__6880\ : Span4Mux_h
    port map (
            O => \N__37218\,
            I => \N__37215\
        );

    \I__6879\ : Odrv4
    port map (
            O => \N__37215\,
            I => \pid_front.error_p_reg_esr_RNI57KP4Z0Z_18\
        );

    \I__6878\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37209\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__37209\,
            I => \pid_front.pid_preregZ0Z_20\
        );

    \I__6876\ : InMux
    port map (
            O => \N__37206\,
            I => \pid_front.un1_pid_prereg_cry_17\
        );

    \I__6875\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37200\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N__37197\
        );

    \I__6873\ : Odrv12
    port map (
            O => \N__37197\,
            I => \pid_front.error_p_reg_esr_RNI8ARC2Z0Z_19\
        );

    \I__6872\ : CascadeMux
    port map (
            O => \N__37194\,
            I => \N__37191\
        );

    \I__6871\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37188\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__37188\,
            I => \N__37185\
        );

    \I__6869\ : Span4Mux_v
    port map (
            O => \N__37185\,
            I => \N__37182\
        );

    \I__6868\ : Odrv4
    port map (
            O => \N__37182\,
            I => \pid_front.error_p_reg_esr_RNIOUOP4Z0Z_19\
        );

    \I__6867\ : InMux
    port map (
            O => \N__37179\,
            I => \N__37176\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__37176\,
            I => \pid_front.pid_preregZ0Z_21\
        );

    \I__6865\ : InMux
    port map (
            O => \N__37173\,
            I => \pid_front.un1_pid_prereg_cry_18\
        );

    \I__6864\ : InMux
    port map (
            O => \N__37170\,
            I => \N__37167\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__37167\,
            I => \N__37164\
        );

    \I__6862\ : Span4Mux_h
    port map (
            O => \N__37164\,
            I => \N__37161\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__37161\,
            I => \pid_front.error_p_reg_esr_RNI09RP4Z0Z_20\
        );

    \I__6860\ : InMux
    port map (
            O => \N__37158\,
            I => \N__37155\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__37155\,
            I => \pid_front.pid_preregZ0Z_22\
        );

    \I__6858\ : InMux
    port map (
            O => \N__37152\,
            I => \pid_front.un1_pid_prereg_cry_19\
        );

    \I__6857\ : InMux
    port map (
            O => \N__37149\,
            I => \pid_front.un1_pid_prereg_cry_20\
        );

    \I__6856\ : CascadeMux
    port map (
            O => \N__37146\,
            I => \N__37143\
        );

    \I__6855\ : InMux
    port map (
            O => \N__37143\,
            I => \N__37136\
        );

    \I__6854\ : InMux
    port map (
            O => \N__37142\,
            I => \N__37131\
        );

    \I__6853\ : InMux
    port map (
            O => \N__37141\,
            I => \N__37131\
        );

    \I__6852\ : InMux
    port map (
            O => \N__37140\,
            I => \N__37128\
        );

    \I__6851\ : CascadeMux
    port map (
            O => \N__37139\,
            I => \N__37125\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__37136\,
            I => \N__37121\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__37131\,
            I => \N__37118\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__37128\,
            I => \N__37115\
        );

    \I__6847\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37110\
        );

    \I__6846\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37110\
        );

    \I__6845\ : Span4Mux_v
    port map (
            O => \N__37121\,
            I => \N__37105\
        );

    \I__6844\ : Span4Mux_v
    port map (
            O => \N__37118\,
            I => \N__37105\
        );

    \I__6843\ : Span4Mux_h
    port map (
            O => \N__37115\,
            I => \N__37102\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__37110\,
            I => \pid_front.pid_preregZ0Z_23\
        );

    \I__6841\ : Odrv4
    port map (
            O => \N__37105\,
            I => \pid_front.pid_preregZ0Z_23\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__37102\,
            I => \pid_front.pid_preregZ0Z_23\
        );

    \I__6839\ : InMux
    port map (
            O => \N__37095\,
            I => \pid_front.un1_pid_prereg_cry_7\
        );

    \I__6838\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37089\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__37089\,
            I => \N__37086\
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__37086\,
            I => \pid_front.error_d_reg_esr_RNI9NAB3Z0Z_10\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__37083\,
            I => \N__37079\
        );

    \I__6834\ : CascadeMux
    port map (
            O => \N__37082\,
            I => \N__37076\
        );

    \I__6833\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37073\
        );

    \I__6832\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37070\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__37073\,
            I => \N__37067\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__37070\,
            I => \pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__37067\,
            I => \pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10\
        );

    \I__6828\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37059\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__37059\,
            I => \N__37056\
        );

    \I__6826\ : Span4Mux_h
    port map (
            O => \N__37056\,
            I => \N__37050\
        );

    \I__6825\ : InMux
    port map (
            O => \N__37055\,
            I => \N__37043\
        );

    \I__6824\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37043\
        );

    \I__6823\ : InMux
    port map (
            O => \N__37053\,
            I => \N__37043\
        );

    \I__6822\ : Odrv4
    port map (
            O => \N__37050\,
            I => \pid_front.pid_preregZ0Z_11\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__37043\,
            I => \pid_front.pid_preregZ0Z_11\
        );

    \I__6820\ : InMux
    port map (
            O => \N__37038\,
            I => \pid_front.un1_pid_prereg_cry_8\
        );

    \I__6819\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37032\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__37032\,
            I => \N__37029\
        );

    \I__6817\ : Span4Mux_h
    port map (
            O => \N__37029\,
            I => \N__37026\
        );

    \I__6816\ : Odrv4
    port map (
            O => \N__37026\,
            I => \pid_front.error_p_reg_esr_RNIESET1Z0Z_10\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__37023\,
            I => \N__37020\
        );

    \I__6814\ : InMux
    port map (
            O => \N__37020\,
            I => \N__37017\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__37017\,
            I => \N__37014\
        );

    \I__6812\ : Span4Mux_h
    port map (
            O => \N__37014\,
            I => \N__37011\
        );

    \I__6811\ : Odrv4
    port map (
            O => \N__37011\,
            I => \pid_front.error_p_reg_esr_RNI1E6A4Z0Z_12\
        );

    \I__6810\ : InMux
    port map (
            O => \N__37008\,
            I => \N__37005\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__37005\,
            I => \N__36999\
        );

    \I__6808\ : InMux
    port map (
            O => \N__37004\,
            I => \N__36992\
        );

    \I__6807\ : InMux
    port map (
            O => \N__37003\,
            I => \N__36992\
        );

    \I__6806\ : InMux
    port map (
            O => \N__37002\,
            I => \N__36992\
        );

    \I__6805\ : Odrv4
    port map (
            O => \N__36999\,
            I => \pid_front.pid_preregZ0Z_12\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__36992\,
            I => \pid_front.pid_preregZ0Z_12\
        );

    \I__6803\ : InMux
    port map (
            O => \N__36987\,
            I => \pid_front.un1_pid_prereg_cry_9\
        );

    \I__6802\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36980\
        );

    \I__6801\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__36980\,
            I => \N__36974\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__36977\,
            I => \pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__36974\,
            I => \pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12\
        );

    \I__6797\ : CascadeMux
    port map (
            O => \N__36969\,
            I => \N__36966\
        );

    \I__6796\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36963\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__36963\,
            I => \N__36960\
        );

    \I__6794\ : Odrv12
    port map (
            O => \N__36960\,
            I => \pid_front.error_d_reg_esr_RNIBO6A4Z0Z_12\
        );

    \I__6793\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36953\
        );

    \I__6792\ : InMux
    port map (
            O => \N__36956\,
            I => \N__36950\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__36953\,
            I => \N__36943\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__36950\,
            I => \N__36943\
        );

    \I__6789\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36937\
        );

    \I__6788\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36937\
        );

    \I__6787\ : Span4Mux_h
    port map (
            O => \N__36943\,
            I => \N__36934\
        );

    \I__6786\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36931\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__36937\,
            I => \pid_front.pid_preregZ0Z_13\
        );

    \I__6784\ : Odrv4
    port map (
            O => \N__36934\,
            I => \pid_front.pid_preregZ0Z_13\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__36931\,
            I => \pid_front.pid_preregZ0Z_13\
        );

    \I__6782\ : InMux
    port map (
            O => \N__36924\,
            I => \pid_front.un1_pid_prereg_cry_10\
        );

    \I__6781\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36918\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__36918\,
            I => \N__36915\
        );

    \I__6779\ : Odrv12
    port map (
            O => \N__36915\,
            I => \pid_front.error_p_reg_esr_RNIO6FT1Z0Z_12\
        );

    \I__6778\ : CascadeMux
    port map (
            O => \N__36912\,
            I => \N__36909\
        );

    \I__6777\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36906\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__36906\,
            I => \N__36903\
        );

    \I__6775\ : Odrv12
    port map (
            O => \N__36903\,
            I => \pid_front.error_p_reg_esr_RNIN47A4Z0Z_12\
        );

    \I__6774\ : InMux
    port map (
            O => \N__36900\,
            I => \N__36897\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__36897\,
            I => \pid_front.pid_preregZ0Z_14\
        );

    \I__6772\ : InMux
    port map (
            O => \N__36894\,
            I => \pid_front.un1_pid_prereg_cry_11\
        );

    \I__6771\ : InMux
    port map (
            O => \N__36891\,
            I => \N__36888\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__36888\,
            I => \N__36885\
        );

    \I__6769\ : Span4Mux_h
    port map (
            O => \N__36885\,
            I => \N__36882\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__36882\,
            I => \pid_front.error_p_reg_esr_RNI42GP4Z0Z_13\
        );

    \I__6767\ : CascadeMux
    port map (
            O => \N__36879\,
            I => \N__36876\
        );

    \I__6766\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36873\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__36873\,
            I => \N__36870\
        );

    \I__6764\ : Span4Mux_h
    port map (
            O => \N__36870\,
            I => \N__36867\
        );

    \I__6763\ : Odrv4
    port map (
            O => \N__36867\,
            I => \pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13\
        );

    \I__6762\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36861\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__36861\,
            I => \pid_front.pid_preregZ0Z_15\
        );

    \I__6760\ : InMux
    port map (
            O => \N__36858\,
            I => \pid_front.un1_pid_prereg_cry_12\
        );

    \I__6759\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36852\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__36852\,
            I => \N__36849\
        );

    \I__6757\ : Odrv12
    port map (
            O => \N__36849\,
            I => \pid_front.error_p_reg_esr_RNI54OC2Z0Z_14\
        );

    \I__6756\ : CascadeMux
    port map (
            O => \N__36846\,
            I => \N__36843\
        );

    \I__6755\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36840\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__36840\,
            I => \N__36837\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__36837\,
            I => \N__36834\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__36834\,
            I => \pid_front.error_p_reg_esr_RNIGEGP4Z0Z_14\
        );

    \I__6751\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36828\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__36828\,
            I => \pid_front.pid_preregZ0Z_16\
        );

    \I__6749\ : InMux
    port map (
            O => \N__36825\,
            I => \bfn_12_23_0_\
        );

    \I__6748\ : InMux
    port map (
            O => \N__36822\,
            I => \N__36819\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__36819\,
            I => \N__36816\
        );

    \I__6746\ : Odrv12
    port map (
            O => \N__36816\,
            I => \pid_front.error_p_reg_esr_RNIBAOC2Z0Z_15\
        );

    \I__6745\ : CascadeMux
    port map (
            O => \N__36813\,
            I => \N__36810\
        );

    \I__6744\ : InMux
    port map (
            O => \N__36810\,
            I => \N__36807\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__36807\,
            I => \N__36804\
        );

    \I__6742\ : Odrv12
    port map (
            O => \N__36804\,
            I => \pid_front.error_p_reg_esr_RNISQGP4Z0Z_15\
        );

    \I__6741\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36798\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__36798\,
            I => \pid_front.pid_preregZ0Z_17\
        );

    \I__6739\ : InMux
    port map (
            O => \N__36795\,
            I => \pid_front.un1_pid_prereg_cry_14\
        );

    \I__6738\ : CascadeMux
    port map (
            O => \N__36792\,
            I => \N__36789\
        );

    \I__6737\ : InMux
    port map (
            O => \N__36789\,
            I => \N__36786\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__36786\,
            I => \N__36783\
        );

    \I__6735\ : Odrv4
    port map (
            O => \N__36783\,
            I => \pid_front.error_p_reg_esr_RNIH7Q01Z0Z_1\
        );

    \I__6734\ : CascadeMux
    port map (
            O => \N__36780\,
            I => \N__36777\
        );

    \I__6733\ : InMux
    port map (
            O => \N__36777\,
            I => \N__36773\
        );

    \I__6732\ : CascadeMux
    port map (
            O => \N__36776\,
            I => \N__36770\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__36773\,
            I => \N__36767\
        );

    \I__6730\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36764\
        );

    \I__6729\ : Span4Mux_h
    port map (
            O => \N__36767\,
            I => \N__36761\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__36764\,
            I => \pid_front.pid_preregZ0Z_3\
        );

    \I__6727\ : Odrv4
    port map (
            O => \N__36761\,
            I => \pid_front.pid_preregZ0Z_3\
        );

    \I__6726\ : InMux
    port map (
            O => \N__36756\,
            I => \pid_front.un1_pid_prereg_cry_0_0\
        );

    \I__6725\ : InMux
    port map (
            O => \N__36753\,
            I => \N__36750\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__36747\,
            I => \pid_front.error_p_reg_esr_RNIJCSGZ0Z_2\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__36744\,
            I => \N__36741\
        );

    \I__6721\ : InMux
    port map (
            O => \N__36741\,
            I => \N__36738\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__36738\,
            I => \N__36735\
        );

    \I__6719\ : Odrv4
    port map (
            O => \N__36735\,
            I => \pid_front.error_p_reg_esr_RNICVO11Z0Z_2\
        );

    \I__6718\ : InMux
    port map (
            O => \N__36732\,
            I => \N__36728\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__36731\,
            I => \N__36720\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__36728\,
            I => \N__36717\
        );

    \I__6715\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36712\
        );

    \I__6714\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36712\
        );

    \I__6713\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36705\
        );

    \I__6712\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36705\
        );

    \I__6711\ : InMux
    port map (
            O => \N__36723\,
            I => \N__36705\
        );

    \I__6710\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36702\
        );

    \I__6709\ : Span4Mux_v
    port map (
            O => \N__36717\,
            I => \N__36699\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__36712\,
            I => \pid_front.pid_preregZ0Z_4\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__36705\,
            I => \pid_front.pid_preregZ0Z_4\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__36702\,
            I => \pid_front.pid_preregZ0Z_4\
        );

    \I__6705\ : Odrv4
    port map (
            O => \N__36699\,
            I => \pid_front.pid_preregZ0Z_4\
        );

    \I__6704\ : InMux
    port map (
            O => \N__36690\,
            I => \pid_front.un1_pid_prereg_cry_1_0\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__36687\,
            I => \N__36682\
        );

    \I__6702\ : CascadeMux
    port map (
            O => \N__36686\,
            I => \N__36679\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__36685\,
            I => \N__36675\
        );

    \I__6700\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36670\
        );

    \I__6699\ : InMux
    port map (
            O => \N__36679\,
            I => \N__36670\
        );

    \I__6698\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36667\
        );

    \I__6697\ : InMux
    port map (
            O => \N__36675\,
            I => \N__36664\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__36670\,
            I => \N__36661\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__36667\,
            I => \N__36658\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__36664\,
            I => \N__36655\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__36661\,
            I => \N__36650\
        );

    \I__6692\ : Span4Mux_h
    port map (
            O => \N__36658\,
            I => \N__36650\
        );

    \I__6691\ : Odrv4
    port map (
            O => \N__36655\,
            I => \pid_front.pid_preregZ0Z_5\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__36650\,
            I => \pid_front.pid_preregZ0Z_5\
        );

    \I__6689\ : InMux
    port map (
            O => \N__36645\,
            I => \pid_front.un1_pid_prereg_cry_2\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__36642\,
            I => \N__36639\
        );

    \I__6687\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36636\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__36636\,
            I => \pid_front.error_p_reg_esr_RNIH8R01Z0Z_5\
        );

    \I__6685\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36630\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__36630\,
            I => \N__36627\
        );

    \I__6683\ : Span4Mux_h
    port map (
            O => \N__36627\,
            I => \N__36622\
        );

    \I__6682\ : InMux
    port map (
            O => \N__36626\,
            I => \N__36619\
        );

    \I__6681\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36616\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__36622\,
            I => \pid_front.pid_preregZ0Z_6\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__36619\,
            I => \pid_front.pid_preregZ0Z_6\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__36616\,
            I => \pid_front.pid_preregZ0Z_6\
        );

    \I__6677\ : InMux
    port map (
            O => \N__36609\,
            I => \pid_front.un1_pid_prereg_cry_3\
        );

    \I__6676\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36602\
        );

    \I__6675\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36599\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__36602\,
            I => \pid_front.error_d_reg_esr_RNIIFUFZ0Z_6\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__36599\,
            I => \pid_front.error_d_reg_esr_RNIIFUFZ0Z_6\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__36594\,
            I => \N__36591\
        );

    \I__6671\ : InMux
    port map (
            O => \N__36591\,
            I => \N__36588\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__36588\,
            I => \pid_front.error_p_reg_esr_RNI94TVZ0Z_6\
        );

    \I__6669\ : InMux
    port map (
            O => \N__36585\,
            I => \N__36582\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__36582\,
            I => \N__36577\
        );

    \I__6667\ : CascadeMux
    port map (
            O => \N__36581\,
            I => \N__36574\
        );

    \I__6666\ : CascadeMux
    port map (
            O => \N__36580\,
            I => \N__36571\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__36577\,
            I => \N__36568\
        );

    \I__6664\ : InMux
    port map (
            O => \N__36574\,
            I => \N__36565\
        );

    \I__6663\ : InMux
    port map (
            O => \N__36571\,
            I => \N__36562\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__36568\,
            I => \pid_front.pid_preregZ0Z_7\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__36565\,
            I => \pid_front.pid_preregZ0Z_7\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__36562\,
            I => \pid_front.pid_preregZ0Z_7\
        );

    \I__6659\ : InMux
    port map (
            O => \N__36555\,
            I => \pid_front.un1_pid_prereg_cry_4\
        );

    \I__6658\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36549\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__36549\,
            I => \N__36546\
        );

    \I__6656\ : Span4Mux_h
    port map (
            O => \N__36546\,
            I => \N__36543\
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__36543\,
            I => \pid_front.error_p_reg_esr_RNIJETVZ0Z_7\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__36540\,
            I => \N__36537\
        );

    \I__6653\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36534\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__36534\,
            I => \N__36531\
        );

    \I__6651\ : Span4Mux_h
    port map (
            O => \N__36531\,
            I => \N__36528\
        );

    \I__6650\ : Odrv4
    port map (
            O => \N__36528\,
            I => \pid_front.error_d_reg_esr_RNINKUFZ0Z_7\
        );

    \I__6649\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36521\
        );

    \I__6648\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36518\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__36521\,
            I => \N__36515\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36511\
        );

    \I__6645\ : Span4Mux_h
    port map (
            O => \N__36515\,
            I => \N__36508\
        );

    \I__6644\ : InMux
    port map (
            O => \N__36514\,
            I => \N__36505\
        );

    \I__6643\ : Span4Mux_h
    port map (
            O => \N__36511\,
            I => \N__36502\
        );

    \I__6642\ : Odrv4
    port map (
            O => \N__36508\,
            I => \pid_front.pid_preregZ0Z_8\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__36505\,
            I => \pid_front.pid_preregZ0Z_8\
        );

    \I__6640\ : Odrv4
    port map (
            O => \N__36502\,
            I => \pid_front.pid_preregZ0Z_8\
        );

    \I__6639\ : InMux
    port map (
            O => \N__36495\,
            I => \bfn_12_22_0_\
        );

    \I__6638\ : InMux
    port map (
            O => \N__36492\,
            I => \N__36489\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__36489\,
            I => \N__36485\
        );

    \I__6636\ : InMux
    port map (
            O => \N__36488\,
            I => \N__36482\
        );

    \I__6635\ : Span4Mux_v
    port map (
            O => \N__36485\,
            I => \N__36479\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__36482\,
            I => \pid_front.error_d_reg_esr_RNISPUFZ0Z_8\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__36479\,
            I => \pid_front.error_d_reg_esr_RNISPUFZ0Z_8\
        );

    \I__6632\ : CascadeMux
    port map (
            O => \N__36474\,
            I => \N__36471\
        );

    \I__6631\ : InMux
    port map (
            O => \N__36471\,
            I => \N__36468\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__36468\,
            I => \N__36465\
        );

    \I__6629\ : Span4Mux_h
    port map (
            O => \N__36465\,
            I => \N__36462\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__36462\,
            I => \pid_front.error_p_reg_esr_RNITOTVZ0Z_8\
        );

    \I__6627\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36456\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__36456\,
            I => \N__36453\
        );

    \I__6625\ : Span4Mux_h
    port map (
            O => \N__36453\,
            I => \N__36448\
        );

    \I__6624\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36445\
        );

    \I__6623\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36442\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__36448\,
            I => \pid_front.pid_preregZ0Z_9\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__36445\,
            I => \pid_front.pid_preregZ0Z_9\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__36442\,
            I => \pid_front.pid_preregZ0Z_9\
        );

    \I__6619\ : InMux
    port map (
            O => \N__36435\,
            I => \pid_front.un1_pid_prereg_cry_6\
        );

    \I__6618\ : InMux
    port map (
            O => \N__36432\,
            I => \N__36429\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__36429\,
            I => \N__36426\
        );

    \I__6616\ : Span4Mux_h
    port map (
            O => \N__36426\,
            I => \N__36423\
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__36423\,
            I => \pid_front.error_d_reg_esr_RNISPQT1Z0Z_10\
        );

    \I__6614\ : CascadeMux
    port map (
            O => \N__36420\,
            I => \N__36416\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__36419\,
            I => \N__36413\
        );

    \I__6612\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36410\
        );

    \I__6611\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36407\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__36410\,
            I => \N__36404\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__36407\,
            I => \N__36401\
        );

    \I__6608\ : Span4Mux_h
    port map (
            O => \N__36404\,
            I => \N__36398\
        );

    \I__6607\ : Span4Mux_v
    port map (
            O => \N__36401\,
            I => \N__36395\
        );

    \I__6606\ : Span4Mux_v
    port map (
            O => \N__36398\,
            I => \N__36392\
        );

    \I__6605\ : Span4Mux_h
    port map (
            O => \N__36395\,
            I => \N__36389\
        );

    \I__6604\ : Span4Mux_v
    port map (
            O => \N__36392\,
            I => \N__36386\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__36389\,
            I => \N__36383\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__36386\,
            I => \pid_front.error_d_reg_esr_RNI1VUFZ0Z_9\
        );

    \I__6601\ : Odrv4
    port map (
            O => \N__36383\,
            I => \pid_front.error_d_reg_esr_RNI1VUFZ0Z_9\
        );

    \I__6600\ : InMux
    port map (
            O => \N__36378\,
            I => \N__36375\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__36375\,
            I => \N__36372\
        );

    \I__6598\ : Span4Mux_h
    port map (
            O => \N__36372\,
            I => \N__36366\
        );

    \I__6597\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36359\
        );

    \I__6596\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36359\
        );

    \I__6595\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36359\
        );

    \I__6594\ : Odrv4
    port map (
            O => \N__36366\,
            I => \pid_front.pid_preregZ0Z_10\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__36359\,
            I => \pid_front.pid_preregZ0Z_10\
        );

    \I__6592\ : CEMux
    port map (
            O => \N__36354\,
            I => \N__36351\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__36351\,
            I => \N__36348\
        );

    \I__6590\ : Span4Mux_v
    port map (
            O => \N__36348\,
            I => \N__36345\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__36345\,
            I => \N__36342\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__36342\,
            I => \dron_frame_decoder_1.N_489_0\
        );

    \I__6587\ : InMux
    port map (
            O => \N__36339\,
            I => \pid_front.un1_pid_prereg_cry_0\
        );

    \I__6586\ : InMux
    port map (
            O => \N__36336\,
            I => \N__36332\
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__36335\,
            I => \N__36329\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__36332\,
            I => \N__36326\
        );

    \I__6583\ : InMux
    port map (
            O => \N__36329\,
            I => \N__36323\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__36326\,
            I => \N__36320\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__36323\,
            I => \pid_front.pid_preregZ0Z_2\
        );

    \I__6580\ : Odrv4
    port map (
            O => \N__36320\,
            I => \pid_front.pid_preregZ0Z_2\
        );

    \I__6579\ : InMux
    port map (
            O => \N__36315\,
            I => \pid_front.un1_pid_prereg_cry_1\
        );

    \I__6578\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36306\
        );

    \I__6577\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36306\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__36306\,
            I => \N__36303\
        );

    \I__6575\ : Span4Mux_v
    port map (
            O => \N__36303\,
            I => \N__36300\
        );

    \I__6574\ : Sp12to4
    port map (
            O => \N__36300\,
            I => \N__36297\
        );

    \I__6573\ : Odrv12
    port map (
            O => \N__36297\,
            I => \pid_front.error_p_regZ0Z_3\
        );

    \I__6572\ : CascadeMux
    port map (
            O => \N__36294\,
            I => \pid_front.un1_pid_prereg_2_cascade_\
        );

    \I__6571\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36285\
        );

    \I__6570\ : InMux
    port map (
            O => \N__36290\,
            I => \N__36285\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__36285\,
            I => \pid_front.un1_pid_prereg_0\
        );

    \I__6568\ : CascadeMux
    port map (
            O => \N__36282\,
            I => \N__36279\
        );

    \I__6567\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36273\
        );

    \I__6566\ : InMux
    port map (
            O => \N__36278\,
            I => \N__36273\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__36273\,
            I => \pid_front.un1_pid_prereg_2\
        );

    \I__6564\ : CascadeMux
    port map (
            O => \N__36270\,
            I => \pid_front.un1_pid_prereg_0_cascade_\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__36267\,
            I => \N__36264\
        );

    \I__6562\ : InMux
    port map (
            O => \N__36264\,
            I => \N__36258\
        );

    \I__6561\ : InMux
    port map (
            O => \N__36263\,
            I => \N__36258\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__36258\,
            I => \pid_front.error_d_reg_prevZ0Z_3\
        );

    \I__6559\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36252\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__36252\,
            I => \drone_H_disp_front_1\
        );

    \I__6557\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36245\
        );

    \I__6556\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36242\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__36245\,
            I => \N__36237\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__36242\,
            I => \N__36237\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__36237\,
            I => \N__36234\
        );

    \I__6552\ : Span4Mux_h
    port map (
            O => \N__36234\,
            I => \N__36231\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__36231\,
            I => throttle_order_0
        );

    \I__6550\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36225\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__36225\,
            I => \N__36222\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__36222\,
            I => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\
        );

    \I__6547\ : InMux
    port map (
            O => \N__36219\,
            I => \N__36216\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__36216\,
            I => \N__36211\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__36215\,
            I => \N__36208\
        );

    \I__6544\ : InMux
    port map (
            O => \N__36214\,
            I => \N__36205\
        );

    \I__6543\ : Span4Mux_h
    port map (
            O => \N__36211\,
            I => \N__36202\
        );

    \I__6542\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36199\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__36205\,
            I => \N__36196\
        );

    \I__6540\ : Span4Mux_h
    port map (
            O => \N__36202\,
            I => \N__36193\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__36199\,
            I => throttle_order_7
        );

    \I__6538\ : Odrv12
    port map (
            O => \N__36196\,
            I => throttle_order_7
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__36193\,
            I => throttle_order_7
        );

    \I__6536\ : InMux
    port map (
            O => \N__36186\,
            I => \N__36183\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__36183\,
            I => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\
        );

    \I__6534\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36177\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__36177\,
            I => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\
        );

    \I__6532\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36171\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__36171\,
            I => \N__36167\
        );

    \I__6530\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36164\
        );

    \I__6529\ : Span4Mux_h
    port map (
            O => \N__36167\,
            I => \N__36161\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__36164\,
            I => \N__36158\
        );

    \I__6527\ : Odrv4
    port map (
            O => \N__36161\,
            I => \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\
        );

    \I__6526\ : Odrv12
    port map (
            O => \N__36158\,
            I => \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\
        );

    \I__6525\ : InMux
    port map (
            O => \N__36153\,
            I => \N__36149\
        );

    \I__6524\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36145\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__36149\,
            I => \N__36142\
        );

    \I__6522\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36139\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__36145\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__36142\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__36139\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__6518\ : InMux
    port map (
            O => \N__36132\,
            I => \N__36129\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__36129\,
            I => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\
        );

    \I__6516\ : InMux
    port map (
            O => \N__36126\,
            I => \N__36121\
        );

    \I__6515\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36118\
        );

    \I__6514\ : CascadeMux
    port map (
            O => \N__36124\,
            I => \N__36115\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__36121\,
            I => \N__36110\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__36118\,
            I => \N__36110\
        );

    \I__6511\ : InMux
    port map (
            O => \N__36115\,
            I => \N__36107\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__36110\,
            I => \N__36104\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__36107\,
            I => \N__36099\
        );

    \I__6508\ : Span4Mux_h
    port map (
            O => \N__36104\,
            I => \N__36099\
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__36099\,
            I => throttle_order_6
        );

    \I__6506\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36093\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__36093\,
            I => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\
        );

    \I__6504\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36087\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__36087\,
            I => \N__36083\
        );

    \I__6502\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36080\
        );

    \I__6501\ : Span4Mux_v
    port map (
            O => \N__36083\,
            I => \N__36077\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__36080\,
            I => \N__36074\
        );

    \I__6499\ : Sp12to4
    port map (
            O => \N__36077\,
            I => \N__36069\
        );

    \I__6498\ : Span12Mux_v
    port map (
            O => \N__36074\,
            I => \N__36069\
        );

    \I__6497\ : Odrv12
    port map (
            O => \N__36069\,
            I => throttle_order_3
        );

    \I__6496\ : InMux
    port map (
            O => \N__36066\,
            I => \N__36062\
        );

    \I__6495\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36059\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__36062\,
            I => \N__36053\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__36059\,
            I => \N__36053\
        );

    \I__6492\ : CascadeMux
    port map (
            O => \N__36058\,
            I => \N__36050\
        );

    \I__6491\ : Span4Mux_h
    port map (
            O => \N__36053\,
            I => \N__36047\
        );

    \I__6490\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36044\
        );

    \I__6489\ : Span4Mux_h
    port map (
            O => \N__36047\,
            I => \N__36041\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__36044\,
            I => throttle_order_9
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__36041\,
            I => throttle_order_9
        );

    \I__6486\ : InMux
    port map (
            O => \N__36036\,
            I => \N__36033\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__36033\,
            I => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\
        );

    \I__6484\ : InMux
    port map (
            O => \N__36030\,
            I => \N__36027\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__36027\,
            I => \N__36024\
        );

    \I__6482\ : Odrv4
    port map (
            O => \N__36024\,
            I => \ppm_encoder_1.un1_aileron_cry_3_THRU_CO\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__36021\,
            I => \N__36017\
        );

    \I__6480\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36014\
        );

    \I__6479\ : InMux
    port map (
            O => \N__36017\,
            I => \N__36011\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__36014\,
            I => \N__36008\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__36011\,
            I => \N__36005\
        );

    \I__6476\ : Span4Mux_h
    port map (
            O => \N__36008\,
            I => \N__36002\
        );

    \I__6475\ : Span4Mux_h
    port map (
            O => \N__36005\,
            I => \N__35999\
        );

    \I__6474\ : Span4Mux_v
    port map (
            O => \N__36002\,
            I => \N__35996\
        );

    \I__6473\ : Span4Mux_h
    port map (
            O => \N__35999\,
            I => \N__35993\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__35996\,
            I => \N__35990\
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__35993\,
            I => throttle_order_4
        );

    \I__6470\ : Odrv4
    port map (
            O => \N__35990\,
            I => throttle_order_4
        );

    \I__6469\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35982\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__35982\,
            I => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\
        );

    \I__6467\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35975\
        );

    \I__6466\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35972\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__35975\,
            I => \N__35966\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__35972\,
            I => \N__35966\
        );

    \I__6463\ : CascadeMux
    port map (
            O => \N__35971\,
            I => \N__35963\
        );

    \I__6462\ : Span4Mux_h
    port map (
            O => \N__35966\,
            I => \N__35960\
        );

    \I__6461\ : InMux
    port map (
            O => \N__35963\,
            I => \N__35957\
        );

    \I__6460\ : Span4Mux_h
    port map (
            O => \N__35960\,
            I => \N__35954\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__35957\,
            I => throttle_order_8
        );

    \I__6458\ : Odrv4
    port map (
            O => \N__35954\,
            I => throttle_order_8
        );

    \I__6457\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35946\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__35946\,
            I => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\
        );

    \I__6455\ : InMux
    port map (
            O => \N__35943\,
            I => \N__35940\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__35940\,
            I => \N__35936\
        );

    \I__6453\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35933\
        );

    \I__6452\ : Span4Mux_h
    port map (
            O => \N__35936\,
            I => \N__35928\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__35933\,
            I => \N__35928\
        );

    \I__6450\ : Span4Mux_h
    port map (
            O => \N__35928\,
            I => \N__35925\
        );

    \I__6449\ : Span4Mux_v
    port map (
            O => \N__35925\,
            I => \N__35922\
        );

    \I__6448\ : Sp12to4
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__6447\ : Odrv12
    port map (
            O => \N__35919\,
            I => throttle_order_12
        );

    \I__6446\ : InMux
    port map (
            O => \N__35916\,
            I => \N__35913\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__35913\,
            I => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\
        );

    \I__6444\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35907\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__35907\,
            I => \N__35904\
        );

    \I__6442\ : Odrv4
    port map (
            O => \N__35904\,
            I => \ppm_encoder_1.un1_aileron_cry_1_THRU_CO\
        );

    \I__6441\ : InMux
    port map (
            O => \N__35901\,
            I => \N__35898\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__35898\,
            I => \frame_decoder_CH4data_4\
        );

    \I__6439\ : CascadeMux
    port map (
            O => \N__35895\,
            I => \N__35892\
        );

    \I__6438\ : InMux
    port map (
            O => \N__35892\,
            I => \N__35889\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__35889\,
            I => \N__35886\
        );

    \I__6436\ : Span4Mux_h
    port map (
            O => \N__35886\,
            I => \N__35883\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__35883\,
            I => \frame_decoder_OFF4data_4\
        );

    \I__6434\ : InMux
    port map (
            O => \N__35880\,
            I => \scaler_4.un3_source_data_0_cry_3\
        );

    \I__6433\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35874\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__35874\,
            I => \frame_decoder_CH4data_5\
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__35871\,
            I => \N__35868\
        );

    \I__6430\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35865\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__35865\,
            I => \N__35862\
        );

    \I__6428\ : Odrv12
    port map (
            O => \N__35862\,
            I => \frame_decoder_OFF4data_5\
        );

    \I__6427\ : InMux
    port map (
            O => \N__35859\,
            I => \scaler_4.un3_source_data_0_cry_4\
        );

    \I__6426\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35853\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__35853\,
            I => \N__35850\
        );

    \I__6424\ : Odrv4
    port map (
            O => \N__35850\,
            I => \frame_decoder_OFF4data_6\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__35847\,
            I => \N__35844\
        );

    \I__6422\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35841\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__35841\,
            I => \frame_decoder_CH4data_6\
        );

    \I__6420\ : InMux
    port map (
            O => \N__35838\,
            I => \scaler_4.un3_source_data_0_cry_5\
        );

    \I__6419\ : InMux
    port map (
            O => \N__35835\,
            I => \N__35832\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__35832\,
            I => \N__35829\
        );

    \I__6417\ : Span4Mux_v
    port map (
            O => \N__35829\,
            I => \N__35826\
        );

    \I__6416\ : Span4Mux_h
    port map (
            O => \N__35826\,
            I => \N__35823\
        );

    \I__6415\ : Odrv4
    port map (
            O => \N__35823\,
            I => \scaler_4.un3_source_data_0_axb_7\
        );

    \I__6414\ : InMux
    port map (
            O => \N__35820\,
            I => \scaler_4.un3_source_data_0_cry_6\
        );

    \I__6413\ : InMux
    port map (
            O => \N__35817\,
            I => \bfn_12_13_0_\
        );

    \I__6412\ : InMux
    port map (
            O => \N__35814\,
            I => \scaler_4.un3_source_data_0_cry_8\
        );

    \I__6411\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35807\
        );

    \I__6410\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35804\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__35807\,
            I => \N__35801\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__35804\,
            I => \N__35798\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__35801\,
            I => \N__35795\
        );

    \I__6406\ : Span12Mux_v
    port map (
            O => \N__35798\,
            I => \N__35792\
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__35795\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__6404\ : Odrv12
    port map (
            O => \N__35792\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__6403\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35784\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__35784\,
            I => \N__35780\
        );

    \I__6401\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35777\
        );

    \I__6400\ : Span4Mux_v
    port map (
            O => \N__35780\,
            I => \N__35774\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__35777\,
            I => \N__35769\
        );

    \I__6398\ : Span4Mux_h
    port map (
            O => \N__35774\,
            I => \N__35769\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__35769\,
            I => \frame_decoder_CH4data_7\
        );

    \I__6396\ : InMux
    port map (
            O => \N__35766\,
            I => \N__35763\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__35763\,
            I => \scaler_4.N_1849_i_l_ofxZ0\
        );

    \I__6394\ : CEMux
    port map (
            O => \N__35760\,
            I => \N__35757\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__35757\,
            I => \N__35754\
        );

    \I__6392\ : Span4Mux_h
    port map (
            O => \N__35754\,
            I => \N__35751\
        );

    \I__6391\ : Odrv4
    port map (
            O => \N__35751\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__6390\ : InMux
    port map (
            O => \N__35748\,
            I => \N__35745\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__35745\,
            I => \frame_decoder_CH4data_1\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__35742\,
            I => \N__35739\
        );

    \I__6387\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35736\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__35736\,
            I => \N__35733\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__35733\,
            I => \frame_decoder_OFF4data_1\
        );

    \I__6384\ : InMux
    port map (
            O => \N__35730\,
            I => \scaler_4.un3_source_data_0_cry_0\
        );

    \I__6383\ : InMux
    port map (
            O => \N__35727\,
            I => \N__35724\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__35724\,
            I => \frame_decoder_CH4data_2\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__35721\,
            I => \N__35718\
        );

    \I__6380\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35715\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__35715\,
            I => \N__35712\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__35712\,
            I => \frame_decoder_OFF4data_2\
        );

    \I__6377\ : InMux
    port map (
            O => \N__35709\,
            I => \scaler_4.un3_source_data_0_cry_1\
        );

    \I__6376\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35703\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__35703\,
            I => \frame_decoder_CH4data_3\
        );

    \I__6374\ : CascadeMux
    port map (
            O => \N__35700\,
            I => \N__35697\
        );

    \I__6373\ : InMux
    port map (
            O => \N__35697\,
            I => \N__35694\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__35694\,
            I => \N__35691\
        );

    \I__6371\ : Odrv4
    port map (
            O => \N__35691\,
            I => \frame_decoder_OFF4data_3\
        );

    \I__6370\ : InMux
    port map (
            O => \N__35688\,
            I => \scaler_4.un3_source_data_0_cry_2\
        );

    \I__6369\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35679\
        );

    \I__6368\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35679\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__35679\,
            I => \pid_front.error_d_reg_prevZ0Z_10\
        );

    \I__6366\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35671\
        );

    \I__6365\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35666\
        );

    \I__6364\ : InMux
    port map (
            O => \N__35674\,
            I => \N__35666\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__35671\,
            I => \pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__35666\,
            I => \pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11\
        );

    \I__6361\ : InMux
    port map (
            O => \N__35661\,
            I => \N__35658\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__35658\,
            I => \N__35654\
        );

    \I__6359\ : InMux
    port map (
            O => \N__35657\,
            I => \N__35651\
        );

    \I__6358\ : Odrv4
    port map (
            O => \N__35654\,
            I => \pid_front.error_p_reg_esr_RNI653NZ0Z_10\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__35651\,
            I => \pid_front.error_p_reg_esr_RNI653NZ0Z_10\
        );

    \I__6356\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35642\
        );

    \I__6355\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35639\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__35642\,
            I => \pid_front.N_1463_i\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__35639\,
            I => \pid_front.N_1463_i\
        );

    \I__6352\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35630\
        );

    \I__6351\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35627\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__35630\,
            I => \N__35622\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__35627\,
            I => \N__35622\
        );

    \I__6348\ : Span4Mux_v
    port map (
            O => \N__35622\,
            I => \N__35619\
        );

    \I__6347\ : Odrv4
    port map (
            O => \N__35619\,
            I => \pid_front.error_p_reg_esr_RNIM6G7Z0Z_9\
        );

    \I__6346\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35612\
        );

    \I__6345\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35609\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__35612\,
            I => \N__35604\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__35609\,
            I => \N__35601\
        );

    \I__6342\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35596\
        );

    \I__6341\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35596\
        );

    \I__6340\ : Span4Mux_h
    port map (
            O => \N__35604\,
            I => \N__35591\
        );

    \I__6339\ : Span4Mux_h
    port map (
            O => \N__35601\,
            I => \N__35591\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__35596\,
            I => \uart_drone.N_152\
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__35591\,
            I => \uart_drone.N_152\
        );

    \I__6336\ : IoInMux
    port map (
            O => \N__35586\,
            I => \N__35583\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__35583\,
            I => \N__35580\
        );

    \I__6334\ : Odrv12
    port map (
            O => \N__35580\,
            I => \pid_side.state_0_0\
        );

    \I__6333\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35573\
        );

    \I__6332\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35568\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__35573\,
            I => \N__35565\
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__35572\,
            I => \N__35561\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__35571\,
            I => \N__35556\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35553\
        );

    \I__6327\ : Span4Mux_v
    port map (
            O => \N__35565\,
            I => \N__35550\
        );

    \I__6326\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35547\
        );

    \I__6325\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35542\
        );

    \I__6324\ : InMux
    port map (
            O => \N__35560\,
            I => \N__35542\
        );

    \I__6323\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35539\
        );

    \I__6322\ : InMux
    port map (
            O => \N__35556\,
            I => \N__35534\
        );

    \I__6321\ : Span4Mux_v
    port map (
            O => \N__35553\,
            I => \N__35531\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__35550\,
            I => \N__35526\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35526\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__35542\,
            I => \N__35521\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__35539\,
            I => \N__35521\
        );

    \I__6316\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35518\
        );

    \I__6315\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35515\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__35534\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6313\ : Odrv4
    port map (
            O => \N__35531\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6312\ : Odrv4
    port map (
            O => \N__35526\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__35521\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__35518\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__35515\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6308\ : InMux
    port map (
            O => \N__35502\,
            I => \N__35499\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__35499\,
            I => \N__35494\
        );

    \I__6306\ : InMux
    port map (
            O => \N__35498\,
            I => \N__35491\
        );

    \I__6305\ : InMux
    port map (
            O => \N__35497\,
            I => \N__35488\
        );

    \I__6304\ : Span4Mux_h
    port map (
            O => \N__35494\,
            I => \N__35480\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__35491\,
            I => \N__35477\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__35488\,
            I => \N__35474\
        );

    \I__6301\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35469\
        );

    \I__6300\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35469\
        );

    \I__6299\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35466\
        );

    \I__6298\ : InMux
    port map (
            O => \N__35484\,
            I => \N__35459\
        );

    \I__6297\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35459\
        );

    \I__6296\ : Span4Mux_v
    port map (
            O => \N__35480\,
            I => \N__35456\
        );

    \I__6295\ : Span4Mux_v
    port map (
            O => \N__35477\,
            I => \N__35447\
        );

    \I__6294\ : Span4Mux_h
    port map (
            O => \N__35474\,
            I => \N__35447\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__35469\,
            I => \N__35447\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__35466\,
            I => \N__35447\
        );

    \I__6291\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35444\
        );

    \I__6290\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35441\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__35459\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__6288\ : Odrv4
    port map (
            O => \N__35456\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__6287\ : Odrv4
    port map (
            O => \N__35447\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__35444\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__35441\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__6284\ : CascadeMux
    port map (
            O => \N__35430\,
            I => \N__35427\
        );

    \I__6283\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35423\
        );

    \I__6282\ : CascadeMux
    port map (
            O => \N__35426\,
            I => \N__35416\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__35423\,
            I => \N__35413\
        );

    \I__6280\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35410\
        );

    \I__6279\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35401\
        );

    \I__6278\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35401\
        );

    \I__6277\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35398\
        );

    \I__6276\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35395\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__35413\,
            I => \N__35390\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__35410\,
            I => \N__35390\
        );

    \I__6273\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35384\
        );

    \I__6272\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35384\
        );

    \I__6271\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35381\
        );

    \I__6270\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35378\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__35401\,
            I => \N__35375\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__35398\,
            I => \N__35370\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__35395\,
            I => \N__35370\
        );

    \I__6266\ : Span4Mux_v
    port map (
            O => \N__35390\,
            I => \N__35367\
        );

    \I__6265\ : InMux
    port map (
            O => \N__35389\,
            I => \N__35364\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__35384\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__35381\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__35378\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6261\ : Odrv4
    port map (
            O => \N__35375\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__35370\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__35367\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__35364\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6257\ : InMux
    port map (
            O => \N__35349\,
            I => \N__35346\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__35346\,
            I => \N__35343\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__35343\,
            I => \uart_drone.data_Auxce_0_3\
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__35340\,
            I => \pid_front.m9_e_4_cascade_\
        );

    \I__6253\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35334\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__35334\,
            I => \pid_front.m9_e_5\
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__35331\,
            I => \N__35327\
        );

    \I__6250\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35322\
        );

    \I__6249\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35319\
        );

    \I__6248\ : InMux
    port map (
            O => \N__35326\,
            I => \N__35313\
        );

    \I__6247\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35313\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__35322\,
            I => \N__35308\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__35319\,
            I => \N__35308\
        );

    \I__6244\ : InMux
    port map (
            O => \N__35318\,
            I => \N__35305\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__35313\,
            I => \pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20\
        );

    \I__6242\ : Odrv4
    port map (
            O => \N__35308\,
            I => \pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__35305\,
            I => \pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20\
        );

    \I__6240\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35291\
        );

    \I__6239\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35291\
        );

    \I__6238\ : InMux
    port map (
            O => \N__35296\,
            I => \N__35288\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__35291\,
            I => \N__35285\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__35288\,
            I => \pid_front.pid_prereg_esr_RNIVDO51Z0Z_10\
        );

    \I__6235\ : Odrv12
    port map (
            O => \N__35285\,
            I => \pid_front.pid_prereg_esr_RNIVDO51Z0Z_10\
        );

    \I__6234\ : InMux
    port map (
            O => \N__35280\,
            I => \N__35277\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__35277\,
            I => \N__35266\
        );

    \I__6232\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35253\
        );

    \I__6231\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35253\
        );

    \I__6230\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35253\
        );

    \I__6229\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35253\
        );

    \I__6228\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35253\
        );

    \I__6227\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35253\
        );

    \I__6226\ : InMux
    port map (
            O => \N__35270\,
            I => \N__35248\
        );

    \I__6225\ : InMux
    port map (
            O => \N__35269\,
            I => \N__35248\
        );

    \I__6224\ : Odrv12
    port map (
            O => \N__35266\,
            I => \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__35253\,
            I => \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__35248\,
            I => \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12\
        );

    \I__6221\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35238\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__35238\,
            I => \N__35235\
        );

    \I__6219\ : Span4Mux_v
    port map (
            O => \N__35235\,
            I => \N__35230\
        );

    \I__6218\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35225\
        );

    \I__6217\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35225\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__35230\,
            I => \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__35225\,
            I => \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13\
        );

    \I__6214\ : CEMux
    port map (
            O => \N__35220\,
            I => \N__35216\
        );

    \I__6213\ : CEMux
    port map (
            O => \N__35219\,
            I => \N__35213\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__35216\,
            I => \N__35210\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__35213\,
            I => \N__35206\
        );

    \I__6210\ : Span4Mux_v
    port map (
            O => \N__35210\,
            I => \N__35203\
        );

    \I__6209\ : CEMux
    port map (
            O => \N__35209\,
            I => \N__35200\
        );

    \I__6208\ : Odrv4
    port map (
            O => \N__35206\,
            I => \pid_front.state_0_1\
        );

    \I__6207\ : Odrv4
    port map (
            O => \N__35203\,
            I => \pid_front.state_0_1\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__35200\,
            I => \pid_front.state_0_1\
        );

    \I__6205\ : SRMux
    port map (
            O => \N__35193\,
            I => \N__35190\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__35190\,
            I => \N__35184\
        );

    \I__6203\ : SRMux
    port map (
            O => \N__35189\,
            I => \N__35181\
        );

    \I__6202\ : SRMux
    port map (
            O => \N__35188\,
            I => \N__35178\
        );

    \I__6201\ : SRMux
    port map (
            O => \N__35187\,
            I => \N__35175\
        );

    \I__6200\ : Span4Mux_v
    port map (
            O => \N__35184\,
            I => \N__35170\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__35181\,
            I => \N__35170\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__35178\,
            I => \N__35163\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__35175\,
            I => \N__35163\
        );

    \I__6196\ : Span4Mux_h
    port map (
            O => \N__35170\,
            I => \N__35163\
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__35163\,
            I => \pid_front.un1_reset_0_i\
        );

    \I__6194\ : CascadeMux
    port map (
            O => \N__35160\,
            I => \pid_front.state_RNIVIRQZ0Z_0_cascade_\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__35157\,
            I => \N__35154\
        );

    \I__6192\ : InMux
    port map (
            O => \N__35154\,
            I => \N__35148\
        );

    \I__6191\ : InMux
    port map (
            O => \N__35153\,
            I => \N__35148\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__35148\,
            I => \N__35145\
        );

    \I__6189\ : Span4Mux_v
    port map (
            O => \N__35145\,
            I => \N__35142\
        );

    \I__6188\ : Span4Mux_v
    port map (
            O => \N__35142\,
            I => \N__35139\
        );

    \I__6187\ : Sp12to4
    port map (
            O => \N__35139\,
            I => \N__35136\
        );

    \I__6186\ : Odrv12
    port map (
            O => \N__35136\,
            I => \pid_front.error_p_regZ0Z_10\
        );

    \I__6185\ : CascadeMux
    port map (
            O => \N__35133\,
            I => \pid_front.error_p_reg_esr_RNI653NZ0Z_10_cascade_\
        );

    \I__6184\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35125\
        );

    \I__6183\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35120\
        );

    \I__6182\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35120\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__35125\,
            I => \N__35114\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__35120\,
            I => \N__35114\
        );

    \I__6179\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35111\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__35114\,
            I => \pid_front.error_d_reg_prevZ0Z_7\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__35111\,
            I => \pid_front.error_d_reg_prevZ0Z_7\
        );

    \I__6176\ : CascadeMux
    port map (
            O => \N__35106\,
            I => \pid_front.m26_e_5_cascade_\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__35103\,
            I => \pid_front.m26_e_1_cascade_\
        );

    \I__6174\ : InMux
    port map (
            O => \N__35100\,
            I => \N__35097\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__35097\,
            I => \pid_front.m26_e_5\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__35094\,
            I => \N__35091\
        );

    \I__6171\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35088\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__35088\,
            I => \pid_front.pid_prereg_esr_RNIGSMQ1Z0Z_10\
        );

    \I__6169\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35082\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__35082\,
            I => \N__35079\
        );

    \I__6167\ : Odrv4
    port map (
            O => \N__35079\,
            I => \pid_front.m18_s_5\
        );

    \I__6166\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35073\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__35073\,
            I => \N__35070\
        );

    \I__6164\ : Odrv4
    port map (
            O => \N__35070\,
            I => \pid_front.m18_s_4\
        );

    \I__6163\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35058\
        );

    \I__6162\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35058\
        );

    \I__6161\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35058\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__35058\,
            I => \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5\
        );

    \I__6159\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35043\
        );

    \I__6158\ : InMux
    port map (
            O => \N__35054\,
            I => \N__35043\
        );

    \I__6157\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35043\
        );

    \I__6156\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35043\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__35043\,
            I => \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10\
        );

    \I__6154\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35034\
        );

    \I__6153\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35031\
        );

    \I__6152\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35026\
        );

    \I__6151\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35026\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__35034\,
            I => \N__35023\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__35031\,
            I => \pid_front.error_p_regZ0Z_7\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__35026\,
            I => \pid_front.error_p_regZ0Z_7\
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__35023\,
            I => \pid_front.error_p_regZ0Z_7\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__35016\,
            I => \pid_front.un1_pid_prereg_60_0_cascade_\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__35013\,
            I => \pid_front.N_1447_i_cascade_\
        );

    \I__6144\ : InMux
    port map (
            O => \N__35010\,
            I => \N__35004\
        );

    \I__6143\ : InMux
    port map (
            O => \N__35009\,
            I => \N__35001\
        );

    \I__6142\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34996\
        );

    \I__6141\ : InMux
    port map (
            O => \N__35007\,
            I => \N__34996\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__35004\,
            I => \N__34989\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__35001\,
            I => \N__34989\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__34996\,
            I => \N__34989\
        );

    \I__6137\ : Span12Mux_h
    port map (
            O => \N__34989\,
            I => \N__34986\
        );

    \I__6136\ : Odrv12
    port map (
            O => \N__34986\,
            I => \pid_front.error_p_regZ0Z_6\
        );

    \I__6135\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34980\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__34980\,
            I => \N__34974\
        );

    \I__6133\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34967\
        );

    \I__6132\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34967\
        );

    \I__6131\ : InMux
    port map (
            O => \N__34977\,
            I => \N__34967\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__34974\,
            I => \pid_front.error_d_reg_prevZ0Z_6\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__34967\,
            I => \pid_front.error_d_reg_prevZ0Z_6\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__34962\,
            I => \pid_front.un1_pid_prereg_50_0_cascade_\
        );

    \I__6127\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34956\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__34956\,
            I => drone_altitude_3
        );

    \I__6125\ : CEMux
    port map (
            O => \N__34953\,
            I => \N__34950\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__34950\,
            I => \N__34947\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__34947\,
            I => \N__34943\
        );

    \I__6122\ : CEMux
    port map (
            O => \N__34946\,
            I => \N__34940\
        );

    \I__6121\ : Sp12to4
    port map (
            O => \N__34943\,
            I => \N__34937\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__34940\,
            I => \N__34934\
        );

    \I__6119\ : Span12Mux_s9_h
    port map (
            O => \N__34937\,
            I => \N__34931\
        );

    \I__6118\ : Span4Mux_v
    port map (
            O => \N__34934\,
            I => \N__34928\
        );

    \I__6117\ : Odrv12
    port map (
            O => \N__34931\,
            I => \dron_frame_decoder_1.N_521_0\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__34928\,
            I => \dron_frame_decoder_1.N_521_0\
        );

    \I__6115\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__34920\,
            I => \N__34917\
        );

    \I__6113\ : Span12Mux_v
    port map (
            O => \N__34917\,
            I => \N__34914\
        );

    \I__6112\ : Odrv12
    port map (
            O => \N__34914\,
            I => \pid_alt.error_d_reg_prevZ0Z_0\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__34911\,
            I => \N__34908\
        );

    \I__6110\ : InMux
    port map (
            O => \N__34908\,
            I => \N__34905\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__34905\,
            I => \N__34901\
        );

    \I__6108\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34898\
        );

    \I__6107\ : Span4Mux_v
    port map (
            O => \N__34901\,
            I => \N__34895\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__34898\,
            I => \N__34892\
        );

    \I__6105\ : Sp12to4
    port map (
            O => \N__34895\,
            I => \N__34887\
        );

    \I__6104\ : Span12Mux_v
    port map (
            O => \N__34892\,
            I => \N__34887\
        );

    \I__6103\ : Odrv12
    port map (
            O => \N__34887\,
            I => \pid_alt.error_d_reg_prev_i_0\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__34884\,
            I => \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12_cascade_\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__34881\,
            I => \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10_cascade_\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__34878\,
            I => \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5_cascade_\
        );

    \I__6099\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34872\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__34872\,
            I => \N__34869\
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__34869\,
            I => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\
        );

    \I__6096\ : InMux
    port map (
            O => \N__34866\,
            I => \ppm_encoder_1.un1_aileron_cry_8\
        );

    \I__6095\ : InMux
    port map (
            O => \N__34863\,
            I => \ppm_encoder_1.un1_aileron_cry_9\
        );

    \I__6094\ : InMux
    port map (
            O => \N__34860\,
            I => \ppm_encoder_1.un1_aileron_cry_10\
        );

    \I__6093\ : InMux
    port map (
            O => \N__34857\,
            I => \ppm_encoder_1.un1_aileron_cry_11\
        );

    \I__6092\ : InMux
    port map (
            O => \N__34854\,
            I => \ppm_encoder_1.un1_aileron_cry_12\
        );

    \I__6091\ : InMux
    port map (
            O => \N__34851\,
            I => \ppm_encoder_1.un1_aileron_cry_13\
        );

    \I__6090\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34845\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__34845\,
            I => \N__34842\
        );

    \I__6088\ : Span12Mux_s7_h
    port map (
            O => \N__34842\,
            I => \N__34839\
        );

    \I__6087\ : Odrv12
    port map (
            O => \N__34839\,
            I => \pid_alt.error_axbZ0Z_2\
        );

    \I__6086\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34833\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__34833\,
            I => drone_altitude_2
        );

    \I__6084\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34827\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__6082\ : Span4Mux_h
    port map (
            O => \N__34824\,
            I => \N__34821\
        );

    \I__6081\ : Span4Mux_h
    port map (
            O => \N__34821\,
            I => \N__34818\
        );

    \I__6080\ : Odrv4
    port map (
            O => \N__34818\,
            I => \pid_alt.error_axbZ0Z_3\
        );

    \I__6079\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34812\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__34812\,
            I => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\
        );

    \I__6077\ : InMux
    port map (
            O => \N__34809\,
            I => \ppm_encoder_1.un1_aileron_cry_0\
        );

    \I__6076\ : InMux
    port map (
            O => \N__34806\,
            I => \ppm_encoder_1.un1_aileron_cry_1\
        );

    \I__6075\ : InMux
    port map (
            O => \N__34803\,
            I => \ppm_encoder_1.un1_aileron_cry_2\
        );

    \I__6074\ : InMux
    port map (
            O => \N__34800\,
            I => \ppm_encoder_1.un1_aileron_cry_3\
        );

    \I__6073\ : InMux
    port map (
            O => \N__34797\,
            I => \ppm_encoder_1.un1_aileron_cry_4\
        );

    \I__6072\ : InMux
    port map (
            O => \N__34794\,
            I => \ppm_encoder_1.un1_aileron_cry_5\
        );

    \I__6071\ : InMux
    port map (
            O => \N__34791\,
            I => \ppm_encoder_1.un1_aileron_cry_6\
        );

    \I__6070\ : InMux
    port map (
            O => \N__34788\,
            I => \bfn_11_18_0_\
        );

    \I__6069\ : InMux
    port map (
            O => \N__34785\,
            I => \bfn_11_15_0_\
        );

    \I__6068\ : InMux
    port map (
            O => \N__34782\,
            I => \ppm_encoder_1.un1_throttle_cry_8\
        );

    \I__6067\ : InMux
    port map (
            O => \N__34779\,
            I => \ppm_encoder_1.un1_throttle_cry_9\
        );

    \I__6066\ : InMux
    port map (
            O => \N__34776\,
            I => \ppm_encoder_1.un1_throttle_cry_10\
        );

    \I__6065\ : InMux
    port map (
            O => \N__34773\,
            I => \ppm_encoder_1.un1_throttle_cry_11\
        );

    \I__6064\ : InMux
    port map (
            O => \N__34770\,
            I => \ppm_encoder_1.un1_throttle_cry_12\
        );

    \I__6063\ : InMux
    port map (
            O => \N__34767\,
            I => \ppm_encoder_1.un1_throttle_cry_13\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__34764\,
            I => \N__34761\
        );

    \I__6061\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34757\
        );

    \I__6060\ : InMux
    port map (
            O => \N__34760\,
            I => \N__34754\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__34757\,
            I => \N__34751\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34748\
        );

    \I__6057\ : Span4Mux_h
    port map (
            O => \N__34751\,
            I => \N__34745\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__34748\,
            I => \N__34742\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__34745\,
            I => \N__34737\
        );

    \I__6054\ : Span4Mux_h
    port map (
            O => \N__34742\,
            I => \N__34737\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__34737\,
            I => throttle_order_13
        );

    \I__6052\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__34731\,
            I => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\
        );

    \I__6050\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34724\
        );

    \I__6049\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34721\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__34724\,
            I => \N__34718\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34714\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__34718\,
            I => \N__34711\
        );

    \I__6045\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34708\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__34714\,
            I => \N__34703\
        );

    \I__6043\ : Span4Mux_h
    port map (
            O => \N__34711\,
            I => \N__34703\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__34708\,
            I => throttle_order_10
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__34703\,
            I => throttle_order_10
        );

    \I__6040\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34695\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__34695\,
            I => \N__34688\
        );

    \I__6038\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34685\
        );

    \I__6037\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34680\
        );

    \I__6036\ : InMux
    port map (
            O => \N__34692\,
            I => \N__34680\
        );

    \I__6035\ : InMux
    port map (
            O => \N__34691\,
            I => \N__34674\
        );

    \I__6034\ : Span4Mux_h
    port map (
            O => \N__34688\,
            I => \N__34667\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__34685\,
            I => \N__34667\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__34680\,
            I => \N__34667\
        );

    \I__6031\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34662\
        );

    \I__6030\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34662\
        );

    \I__6029\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34659\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__34674\,
            I => \N__34656\
        );

    \I__6027\ : Span4Mux_v
    port map (
            O => \N__34667\,
            I => \N__34649\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__34662\,
            I => \N__34649\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__34659\,
            I => \N__34649\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__34656\,
            I => \dron_frame_decoder_1.N_218\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__34649\,
            I => \dron_frame_decoder_1.N_218\
        );

    \I__6022\ : InMux
    port map (
            O => \N__34644\,
            I => \ppm_encoder_1.un1_throttle_cry_0\
        );

    \I__6021\ : InMux
    port map (
            O => \N__34641\,
            I => \ppm_encoder_1.un1_throttle_cry_1\
        );

    \I__6020\ : InMux
    port map (
            O => \N__34638\,
            I => \ppm_encoder_1.un1_throttle_cry_2\
        );

    \I__6019\ : InMux
    port map (
            O => \N__34635\,
            I => \ppm_encoder_1.un1_throttle_cry_3\
        );

    \I__6018\ : InMux
    port map (
            O => \N__34632\,
            I => \N__34628\
        );

    \I__6017\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34625\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__34628\,
            I => \N__34622\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__34625\,
            I => \N__34619\
        );

    \I__6014\ : Span4Mux_h
    port map (
            O => \N__34622\,
            I => \N__34616\
        );

    \I__6013\ : Span4Mux_h
    port map (
            O => \N__34619\,
            I => \N__34613\
        );

    \I__6012\ : Span4Mux_v
    port map (
            O => \N__34616\,
            I => \N__34610\
        );

    \I__6011\ : Span4Mux_v
    port map (
            O => \N__34613\,
            I => \N__34607\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__34610\,
            I => \N__34604\
        );

    \I__6009\ : Span4Mux_h
    port map (
            O => \N__34607\,
            I => \N__34601\
        );

    \I__6008\ : Odrv4
    port map (
            O => \N__34604\,
            I => throttle_order_5
        );

    \I__6007\ : Odrv4
    port map (
            O => \N__34601\,
            I => throttle_order_5
        );

    \I__6006\ : InMux
    port map (
            O => \N__34596\,
            I => \N__34593\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__34593\,
            I => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\
        );

    \I__6004\ : InMux
    port map (
            O => \N__34590\,
            I => \ppm_encoder_1.un1_throttle_cry_4\
        );

    \I__6003\ : InMux
    port map (
            O => \N__34587\,
            I => \ppm_encoder_1.un1_throttle_cry_5\
        );

    \I__6002\ : InMux
    port map (
            O => \N__34584\,
            I => \ppm_encoder_1.un1_throttle_cry_6\
        );

    \I__6001\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34576\
        );

    \I__6000\ : InMux
    port map (
            O => \N__34580\,
            I => \N__34571\
        );

    \I__5999\ : InMux
    port map (
            O => \N__34579\,
            I => \N__34571\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__34576\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__34571\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__5996\ : InMux
    port map (
            O => \N__34566\,
            I => \dron_frame_decoder_1.un1_WDT_cry_13\
        );

    \I__5995\ : InMux
    port map (
            O => \N__34563\,
            I => \dron_frame_decoder_1.un1_WDT_cry_14\
        );

    \I__5994\ : CascadeMux
    port map (
            O => \N__34560\,
            I => \N__34556\
        );

    \I__5993\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34552\
        );

    \I__5992\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34547\
        );

    \I__5991\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34547\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__34552\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__34547\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__5988\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34538\
        );

    \I__5987\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34535\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34532\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__34535\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__5984\ : Odrv12
    port map (
            O => \N__34532\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__5983\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34523\
        );

    \I__5982\ : InMux
    port map (
            O => \N__34526\,
            I => \N__34520\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__34523\,
            I => \N__34517\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__34520\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__34517\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__5978\ : CascadeMux
    port map (
            O => \N__34512\,
            I => \N__34509\
        );

    \I__5977\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34505\
        );

    \I__5976\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34502\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34499\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__34502\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__34499\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__5972\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34490\
        );

    \I__5971\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34487\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__34490\,
            I => \N__34484\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__34487\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__5968\ : Odrv4
    port map (
            O => \N__34484\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__5967\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34475\
        );

    \I__5966\ : InMux
    port map (
            O => \N__34478\,
            I => \N__34472\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__34475\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__34472\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__34467\,
            I => \dron_frame_decoder_1.WDT_RNIIVJ1Z0Z_4_cascade_\
        );

    \I__5962\ : InMux
    port map (
            O => \N__34464\,
            I => \N__34458\
        );

    \I__5961\ : InMux
    port map (
            O => \N__34463\,
            I => \N__34458\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__34458\,
            I => \dron_frame_decoder_1.WDT10lt14_0\
        );

    \I__5959\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34451\
        );

    \I__5958\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34448\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__34451\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__34448\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__34443\,
            I => \N__34439\
        );

    \I__5954\ : InMux
    port map (
            O => \N__34442\,
            I => \N__34436\
        );

    \I__5953\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34433\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__34436\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__34433\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__5950\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34425\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__34425\,
            I => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\
        );

    \I__5948\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34417\
        );

    \I__5947\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34412\
        );

    \I__5946\ : InMux
    port map (
            O => \N__34420\,
            I => \N__34412\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__34417\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__34412\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__5943\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34403\
        );

    \I__5942\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34400\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__34403\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__34400\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__5939\ : CascadeMux
    port map (
            O => \N__34395\,
            I => \N__34390\
        );

    \I__5938\ : InMux
    port map (
            O => \N__34394\,
            I => \N__34387\
        );

    \I__5937\ : InMux
    port map (
            O => \N__34393\,
            I => \N__34382\
        );

    \I__5936\ : InMux
    port map (
            O => \N__34390\,
            I => \N__34382\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__34387\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__34382\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__5933\ : InMux
    port map (
            O => \N__34377\,
            I => \N__34374\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__34374\,
            I => \dron_frame_decoder_1.WDT10lto13_1\
        );

    \I__5931\ : CascadeMux
    port map (
            O => \N__34371\,
            I => \N__34367\
        );

    \I__5930\ : CascadeMux
    port map (
            O => \N__34370\,
            I => \N__34363\
        );

    \I__5929\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34360\
        );

    \I__5928\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34357\
        );

    \I__5927\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34354\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__34360\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__34357\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__34354\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__5923\ : InMux
    port map (
            O => \N__34347\,
            I => \dron_frame_decoder_1.un1_WDT_cry_4\
        );

    \I__5922\ : InMux
    port map (
            O => \N__34344\,
            I => \dron_frame_decoder_1.un1_WDT_cry_5\
        );

    \I__5921\ : InMux
    port map (
            O => \N__34341\,
            I => \dron_frame_decoder_1.un1_WDT_cry_6\
        );

    \I__5920\ : InMux
    port map (
            O => \N__34338\,
            I => \bfn_11_11_0_\
        );

    \I__5919\ : InMux
    port map (
            O => \N__34335\,
            I => \dron_frame_decoder_1.un1_WDT_cry_8\
        );

    \I__5918\ : InMux
    port map (
            O => \N__34332\,
            I => \dron_frame_decoder_1.un1_WDT_cry_9\
        );

    \I__5917\ : InMux
    port map (
            O => \N__34329\,
            I => \dron_frame_decoder_1.un1_WDT_cry_10\
        );

    \I__5916\ : InMux
    port map (
            O => \N__34326\,
            I => \dron_frame_decoder_1.un1_WDT_cry_11\
        );

    \I__5915\ : InMux
    port map (
            O => \N__34323\,
            I => \dron_frame_decoder_1.un1_WDT_cry_12\
        );

    \I__5914\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34317\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__34317\,
            I => \uart_drone.data_Auxce_0_1\
        );

    \I__5912\ : InMux
    port map (
            O => \N__34314\,
            I => \N__34310\
        );

    \I__5911\ : InMux
    port map (
            O => \N__34313\,
            I => \N__34307\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__34310\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__34307\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__5908\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34298\
        );

    \I__5907\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34295\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__34298\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__34295\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__34290\,
            I => \N__34287\
        );

    \I__5903\ : InMux
    port map (
            O => \N__34287\,
            I => \N__34283\
        );

    \I__5902\ : InMux
    port map (
            O => \N__34286\,
            I => \N__34280\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__34283\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__34280\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__5899\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34269\
        );

    \I__5898\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34269\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__34269\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__34266\,
            I => \N__34263\
        );

    \I__5895\ : InMux
    port map (
            O => \N__34263\,
            I => \N__34254\
        );

    \I__5894\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34254\
        );

    \I__5893\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34254\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__34254\,
            I => \N__34251\
        );

    \I__5891\ : Span4Mux_h
    port map (
            O => \N__34251\,
            I => \N__34247\
        );

    \I__5890\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34244\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__34247\,
            I => \reset_module_System.reset6_14\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__34244\,
            I => \reset_module_System.reset6_14\
        );

    \I__5887\ : InMux
    port map (
            O => \N__34239\,
            I => \N__34233\
        );

    \I__5886\ : InMux
    port map (
            O => \N__34238\,
            I => \N__34233\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__34233\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__5884\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34226\
        );

    \I__5883\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34223\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__34226\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__34223\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__34218\,
            I => \N__34214\
        );

    \I__5879\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34209\
        );

    \I__5878\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34209\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__34209\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__5876\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34202\
        );

    \I__5875\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34199\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__34202\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__34199\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__5872\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34191\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__34191\,
            I => \reset_module_System.reset6_11\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__34188\,
            I => \N__34184\
        );

    \I__5869\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34181\
        );

    \I__5868\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34178\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__34181\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__34178\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__5865\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34170\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__34170\,
            I => \dron_frame_decoder_1.WDTZ0Z_0\
        );

    \I__5863\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34164\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__34164\,
            I => \dron_frame_decoder_1.WDTZ0Z_1\
        );

    \I__5861\ : InMux
    port map (
            O => \N__34161\,
            I => \dron_frame_decoder_1.un1_WDT_cry_0\
        );

    \I__5860\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34155\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__34155\,
            I => \dron_frame_decoder_1.WDTZ0Z_2\
        );

    \I__5858\ : InMux
    port map (
            O => \N__34152\,
            I => \dron_frame_decoder_1.un1_WDT_cry_1\
        );

    \I__5857\ : InMux
    port map (
            O => \N__34149\,
            I => \N__34146\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__34146\,
            I => \dron_frame_decoder_1.WDTZ0Z_3\
        );

    \I__5855\ : InMux
    port map (
            O => \N__34143\,
            I => \dron_frame_decoder_1.un1_WDT_cry_2\
        );

    \I__5854\ : InMux
    port map (
            O => \N__34140\,
            I => \dron_frame_decoder_1.un1_WDT_cry_3\
        );

    \I__5853\ : InMux
    port map (
            O => \N__34137\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__5852\ : InMux
    port map (
            O => \N__34134\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__5851\ : InMux
    port map (
            O => \N__34131\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__5850\ : InMux
    port map (
            O => \N__34128\,
            I => \N__34124\
        );

    \I__5849\ : InMux
    port map (
            O => \N__34127\,
            I => \N__34121\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__34124\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__34121\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__5846\ : InMux
    port map (
            O => \N__34116\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__5845\ : InMux
    port map (
            O => \N__34113\,
            I => \bfn_11_9_0_\
        );

    \I__5844\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34106\
        );

    \I__5843\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34103\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__34106\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__34103\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__5840\ : InMux
    port map (
            O => \N__34098\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__5839\ : InMux
    port map (
            O => \N__34095\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__34092\,
            I => \N__34089\
        );

    \I__5837\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34085\
        );

    \I__5836\ : InMux
    port map (
            O => \N__34088\,
            I => \N__34082\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__34085\,
            I => \N__34079\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__34082\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__5833\ : Odrv4
    port map (
            O => \N__34079\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__5832\ : InMux
    port map (
            O => \N__34074\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__5831\ : InMux
    port map (
            O => \N__34071\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__5830\ : InMux
    port map (
            O => \N__34068\,
            I => \N__34064\
        );

    \I__5829\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34061\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__34064\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__34061\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__5826\ : InMux
    port map (
            O => \N__34056\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__5825\ : InMux
    port map (
            O => \N__34053\,
            I => \N__34049\
        );

    \I__5824\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34046\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__34049\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__34046\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__5821\ : InMux
    port map (
            O => \N__34041\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__5820\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34034\
        );

    \I__5819\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34031\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__34034\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__34031\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__5816\ : InMux
    port map (
            O => \N__34026\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__5815\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34019\
        );

    \I__5814\ : InMux
    port map (
            O => \N__34022\,
            I => \N__34016\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__34019\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__34016\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__5811\ : InMux
    port map (
            O => \N__34011\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__5810\ : CascadeMux
    port map (
            O => \N__34008\,
            I => \N__34004\
        );

    \I__5809\ : InMux
    port map (
            O => \N__34007\,
            I => \N__34001\
        );

    \I__5808\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33998\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__34001\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__33998\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__5805\ : InMux
    port map (
            O => \N__33993\,
            I => \bfn_11_8_0_\
        );

    \I__5804\ : InMux
    port map (
            O => \N__33990\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__5803\ : InMux
    port map (
            O => \N__33987\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__5802\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33980\
        );

    \I__5801\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33977\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__33980\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__33977\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__5798\ : InMux
    port map (
            O => \N__33972\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__5797\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33965\
        );

    \I__5796\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33962\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__33965\,
            I => \N__33959\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__33962\,
            I => \N__33954\
        );

    \I__5793\ : Span4Mux_v
    port map (
            O => \N__33959\,
            I => \N__33954\
        );

    \I__5792\ : Span4Mux_h
    port map (
            O => \N__33954\,
            I => \N__33951\
        );

    \I__5791\ : Span4Mux_v
    port map (
            O => \N__33951\,
            I => \N__33948\
        );

    \I__5790\ : Odrv4
    port map (
            O => \N__33948\,
            I => \pid_front.error_p_regZ0Z_11\
        );

    \I__5789\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33939\
        );

    \I__5788\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33939\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__33939\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__5786\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33933\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__33933\,
            I => \uart_drone.CO0\
        );

    \I__5784\ : InMux
    port map (
            O => \N__33930\,
            I => \N__33923\
        );

    \I__5783\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33923\
        );

    \I__5782\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33920\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__33923\,
            I => \N__33913\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__33920\,
            I => \N__33913\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__33919\,
            I => \N__33907\
        );

    \I__5778\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33904\
        );

    \I__5777\ : Span4Mux_h
    port map (
            O => \N__33913\,
            I => \N__33901\
        );

    \I__5776\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33898\
        );

    \I__5775\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33891\
        );

    \I__5774\ : InMux
    port map (
            O => \N__33910\,
            I => \N__33891\
        );

    \I__5773\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33891\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__33904\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__33901\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__33898\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__33891\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__33882\,
            I => \N__33878\
        );

    \I__5767\ : CascadeMux
    port map (
            O => \N__33881\,
            I => \N__33875\
        );

    \I__5766\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33869\
        );

    \I__5765\ : InMux
    port map (
            O => \N__33875\,
            I => \N__33869\
        );

    \I__5764\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33866\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__33869\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__33866\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__33861\,
            I => \N__33856\
        );

    \I__5760\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33853\
        );

    \I__5759\ : InMux
    port map (
            O => \N__33859\,
            I => \N__33848\
        );

    \I__5758\ : InMux
    port map (
            O => \N__33856\,
            I => \N__33845\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__33853\,
            I => \N__33842\
        );

    \I__5756\ : InMux
    port map (
            O => \N__33852\,
            I => \N__33837\
        );

    \I__5755\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33837\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33831\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__33845\,
            I => \N__33831\
        );

    \I__5752\ : Span4Mux_v
    port map (
            O => \N__33842\,
            I => \N__33826\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33826\
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__33836\,
            I => \N__33822\
        );

    \I__5749\ : Span4Mux_h
    port map (
            O => \N__33831\,
            I => \N__33818\
        );

    \I__5748\ : Span4Mux_h
    port map (
            O => \N__33826\,
            I => \N__33815\
        );

    \I__5747\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33812\
        );

    \I__5746\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33807\
        );

    \I__5745\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33807\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__33818\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__33815\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__33812\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__33807\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__5740\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33794\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__33797\,
            I => \N__33791\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__33794\,
            I => \N__33782\
        );

    \I__5737\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33777\
        );

    \I__5736\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33777\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__33789\,
            I => \N__33773\
        );

    \I__5734\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33770\
        );

    \I__5733\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33763\
        );

    \I__5732\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33763\
        );

    \I__5731\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33763\
        );

    \I__5730\ : Span4Mux_h
    port map (
            O => \N__33782\,
            I => \N__33760\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__33777\,
            I => \N__33757\
        );

    \I__5728\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33752\
        );

    \I__5727\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33752\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__33770\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__33763\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__33760\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__33757\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__33752\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__5721\ : InMux
    port map (
            O => \N__33741\,
            I => \N__33738\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__33735\,
            I => \N__33731\
        );

    \I__5718\ : InMux
    port map (
            O => \N__33734\,
            I => \N__33728\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__33731\,
            I => \uart_drone.N_144_1\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__33728\,
            I => \uart_drone.N_144_1\
        );

    \I__5715\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33718\
        );

    \I__5714\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33715\
        );

    \I__5713\ : InMux
    port map (
            O => \N__33721\,
            I => \N__33712\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__33718\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__33715\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__33712\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__33705\,
            I => \N__33699\
        );

    \I__5708\ : InMux
    port map (
            O => \N__33704\,
            I => \N__33694\
        );

    \I__5707\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33694\
        );

    \I__5706\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33691\
        );

    \I__5705\ : InMux
    port map (
            O => \N__33699\,
            I => \N__33688\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__33694\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__33691\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__33688\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__5701\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33677\
        );

    \I__5700\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33674\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__33677\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__33674\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__5697\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33666\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__33666\,
            I => \reset_module_System.count_1_2\
        );

    \I__5695\ : InMux
    port map (
            O => \N__33663\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__5694\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33656\
        );

    \I__5693\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33653\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__33656\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__33653\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__5690\ : InMux
    port map (
            O => \N__33648\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__5689\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33641\
        );

    \I__5688\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33638\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__33641\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__33638\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__5685\ : InMux
    port map (
            O => \N__33633\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__5684\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33627\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33624\
        );

    \I__5682\ : Odrv4
    port map (
            O => \N__33624\,
            I => \pid_front.pid_prereg_esr_RNI6FQ75Z0Z_23\
        );

    \I__5681\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33617\
        );

    \I__5680\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33614\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__33617\,
            I => \pid_front.un1_pid_prereg_42\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__33614\,
            I => \pid_front.un1_pid_prereg_42\
        );

    \I__5677\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33606\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__33606\,
            I => \N__33601\
        );

    \I__5675\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33596\
        );

    \I__5674\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33596\
        );

    \I__5673\ : Span4Mux_v
    port map (
            O => \N__33601\,
            I => \N__33593\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33590\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__33593\,
            I => \pid_front.un1_pid_prereg_47\
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__33590\,
            I => \pid_front.un1_pid_prereg_47\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__33585\,
            I => \pid_front.un1_pid_prereg_42_cascade_\
        );

    \I__5668\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33578\
        );

    \I__5667\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33575\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33570\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__33575\,
            I => \N__33570\
        );

    \I__5664\ : Span4Mux_v
    port map (
            O => \N__33570\,
            I => \N__33567\
        );

    \I__5663\ : Span4Mux_h
    port map (
            O => \N__33567\,
            I => \N__33564\
        );

    \I__5662\ : Span4Mux_h
    port map (
            O => \N__33564\,
            I => \N__33561\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__33561\,
            I => \pid_front.error_p_regZ0Z_16\
        );

    \I__5660\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33555\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__33555\,
            I => \N__33551\
        );

    \I__5658\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33548\
        );

    \I__5657\ : Span4Mux_v
    port map (
            O => \N__33551\,
            I => \N__33543\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__33548\,
            I => \N__33543\
        );

    \I__5655\ : Span4Mux_v
    port map (
            O => \N__33543\,
            I => \N__33540\
        );

    \I__5654\ : Odrv4
    port map (
            O => \N__33540\,
            I => \pid_front.error_d_reg_prevZ0Z_16\
        );

    \I__5653\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33530\
        );

    \I__5652\ : InMux
    port map (
            O => \N__33536\,
            I => \N__33530\
        );

    \I__5651\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33527\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__33530\,
            I => \N__33524\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__33527\,
            I => \N__33519\
        );

    \I__5648\ : Span4Mux_h
    port map (
            O => \N__33524\,
            I => \N__33519\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__33519\,
            I => \pid_front.un1_pid_prereg_35\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__33516\,
            I => \pid_front.un1_pid_prereg_36_cascade_\
        );

    \I__5645\ : InMux
    port map (
            O => \N__33513\,
            I => \N__33510\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__33510\,
            I => \N__33506\
        );

    \I__5643\ : InMux
    port map (
            O => \N__33509\,
            I => \N__33503\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__33506\,
            I => \pid_front.un1_pid_prereg_30\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__33503\,
            I => \pid_front.un1_pid_prereg_30\
        );

    \I__5640\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33492\
        );

    \I__5639\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33492\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__33492\,
            I => \N__33489\
        );

    \I__5637\ : Span4Mux_v
    port map (
            O => \N__33489\,
            I => \N__33486\
        );

    \I__5636\ : Sp12to4
    port map (
            O => \N__33486\,
            I => \N__33483\
        );

    \I__5635\ : Span12Mux_h
    port map (
            O => \N__33483\,
            I => \N__33480\
        );

    \I__5634\ : Odrv12
    port map (
            O => \N__33480\,
            I => \pid_front.error_p_regZ0Z_17\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__5632\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33468\
        );

    \I__5631\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33468\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__33468\,
            I => \pid_front.error_d_reg_prevZ0Z_17\
        );

    \I__5629\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33459\
        );

    \I__5628\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33459\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__33459\,
            I => \pid_front.un1_pid_prereg_41\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__33456\,
            I => \pid_front.un1_pid_prereg_41_cascade_\
        );

    \I__5625\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33449\
        );

    \I__5624\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33446\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__33449\,
            I => \pid_front.un1_pid_prereg_36\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__33446\,
            I => \pid_front.un1_pid_prereg_36\
        );

    \I__5621\ : InMux
    port map (
            O => \N__33441\,
            I => \N__33438\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__33438\,
            I => \pid_front.un1_reset_0_i_sn\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__33435\,
            I => \N__33432\
        );

    \I__5618\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33429\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33425\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__33428\,
            I => \N__33421\
        );

    \I__5615\ : Span12Mux_v
    port map (
            O => \N__33425\,
            I => \N__33417\
        );

    \I__5614\ : InMux
    port map (
            O => \N__33424\,
            I => \N__33412\
        );

    \I__5613\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33412\
        );

    \I__5612\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33409\
        );

    \I__5611\ : Odrv12
    port map (
            O => \N__33417\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__33412\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__33409\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__5608\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__5606\ : Span4Mux_h
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__5605\ : Span4Mux_h
    port map (
            O => \N__33393\,
            I => \N__33390\
        );

    \I__5604\ : Span4Mux_v
    port map (
            O => \N__33390\,
            I => \N__33382\
        );

    \I__5603\ : InMux
    port map (
            O => \N__33389\,
            I => \N__33371\
        );

    \I__5602\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33371\
        );

    \I__5601\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33371\
        );

    \I__5600\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33371\
        );

    \I__5599\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33371\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__33382\,
            I => \pid_alt.N_62_mux\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__33371\,
            I => \pid_alt.N_62_mux\
        );

    \I__5596\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33363\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__33363\,
            I => \N__33360\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__33360\,
            I => \N__33357\
        );

    \I__5593\ : Span4Mux_v
    port map (
            O => \N__33357\,
            I => \N__33353\
        );

    \I__5592\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33350\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__33353\,
            I => \N__33347\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__33350\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__33347\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__5588\ : SRMux
    port map (
            O => \N__33342\,
            I => \N__33339\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__33339\,
            I => \N__33335\
        );

    \I__5586\ : SRMux
    port map (
            O => \N__33338\,
            I => \N__33332\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__33335\,
            I => \N__33327\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33324\
        );

    \I__5583\ : SRMux
    port map (
            O => \N__33331\,
            I => \N__33321\
        );

    \I__5582\ : SRMux
    port map (
            O => \N__33330\,
            I => \N__33318\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__33327\,
            I => \N__33315\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__33324\,
            I => \N__33310\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__33321\,
            I => \N__33310\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__33318\,
            I => \N__33307\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__33315\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__33310\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__5575\ : Odrv4
    port map (
            O => \N__33307\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__5574\ : CascadeMux
    port map (
            O => \N__33300\,
            I => \N__33297\
        );

    \I__5573\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__33294\,
            I => \N__33290\
        );

    \I__5571\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33287\
        );

    \I__5570\ : Span4Mux_h
    port map (
            O => \N__33290\,
            I => \N__33284\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__33287\,
            I => \N__33281\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__33284\,
            I => \pid_front.un1_pid_prereg_57\
        );

    \I__5567\ : Odrv4
    port map (
            O => \N__33281\,
            I => \pid_front.un1_pid_prereg_57\
        );

    \I__5566\ : InMux
    port map (
            O => \N__33276\,
            I => \N__33273\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__33273\,
            I => \N__33269\
        );

    \I__5564\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33266\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__33269\,
            I => \N__33263\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__33266\,
            I => \N__33260\
        );

    \I__5561\ : Span4Mux_v
    port map (
            O => \N__33263\,
            I => \N__33257\
        );

    \I__5560\ : Sp12to4
    port map (
            O => \N__33260\,
            I => \N__33254\
        );

    \I__5559\ : Sp12to4
    port map (
            O => \N__33257\,
            I => \N__33249\
        );

    \I__5558\ : Span12Mux_v
    port map (
            O => \N__33254\,
            I => \N__33249\
        );

    \I__5557\ : Odrv12
    port map (
            O => \N__33249\,
            I => \pid_front.error_p_regZ0Z_18\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__33246\,
            I => \N__33242\
        );

    \I__5555\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33238\
        );

    \I__5554\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33233\
        );

    \I__5553\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33233\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33230\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__33233\,
            I => \N__33227\
        );

    \I__5550\ : Span4Mux_h
    port map (
            O => \N__33230\,
            I => \N__33224\
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__33227\,
            I => \pid_front.un1_pid_prereg_18\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__33224\,
            I => \pid_front.un1_pid_prereg_18\
        );

    \I__5547\ : InMux
    port map (
            O => \N__33219\,
            I => \N__33213\
        );

    \I__5546\ : InMux
    port map (
            O => \N__33218\,
            I => \N__33213\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__33213\,
            I => \N__33210\
        );

    \I__5544\ : Span4Mux_v
    port map (
            O => \N__33210\,
            I => \N__33207\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__33207\,
            I => \N__33204\
        );

    \I__5542\ : Sp12to4
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__5541\ : Odrv12
    port map (
            O => \N__33201\,
            I => \pid_front.error_p_regZ0Z_13\
        );

    \I__5540\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33192\
        );

    \I__5539\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33192\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__33192\,
            I => \pid_front.error_d_reg_prevZ0Z_13\
        );

    \I__5537\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33183\
        );

    \I__5536\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33183\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33179\
        );

    \I__5534\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33176\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__33179\,
            I => \pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__33176\,
            I => \pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__33171\,
            I => \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13_cascade_\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__33168\,
            I => \pid_front.pid_prereg_esr_RNICUKFAZ0Z_6_cascade_\
        );

    \I__5529\ : CascadeMux
    port map (
            O => \N__33165\,
            I => \pid_front.un1_reset_0_i_cascade_\
        );

    \I__5528\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33159\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__33159\,
            I => \pid_front.un1_reset_0_i_rn_0\
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__33156\,
            I => \pid_front.m32_1_cascade_\
        );

    \I__5525\ : InMux
    port map (
            O => \N__33153\,
            I => \N__33150\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__33150\,
            I => \N__33147\
        );

    \I__5523\ : Odrv12
    port map (
            O => \N__33147\,
            I => \pid_front.O_0_5\
        );

    \I__5522\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33138\
        );

    \I__5521\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33138\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__33138\,
            I => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\
        );

    \I__5519\ : CascadeMux
    port map (
            O => \N__33135\,
            I => \N__33132\
        );

    \I__5518\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33120\
        );

    \I__5517\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33120\
        );

    \I__5516\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33120\
        );

    \I__5515\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33120\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__33120\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__33117\,
            I => \N__33113\
        );

    \I__5512\ : CascadeMux
    port map (
            O => \N__33116\,
            I => \N__33110\
        );

    \I__5511\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33102\
        );

    \I__5510\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33102\
        );

    \I__5509\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33099\
        );

    \I__5508\ : InMux
    port map (
            O => \N__33108\,
            I => \N__33094\
        );

    \I__5507\ : InMux
    port map (
            O => \N__33107\,
            I => \N__33094\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__33102\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__33099\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__33094\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__5503\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__33084\,
            I => \dron_frame_decoder_1.drone_H_disp_side_10\
        );

    \I__5501\ : CEMux
    port map (
            O => \N__33081\,
            I => \N__33078\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__33078\,
            I => \N__33074\
        );

    \I__5499\ : CEMux
    port map (
            O => \N__33077\,
            I => \N__33071\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__33074\,
            I => \N__33068\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__33071\,
            I => \N__33065\
        );

    \I__5496\ : Odrv4
    port map (
            O => \N__33068\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__33065\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__5494\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33057\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__33057\,
            I => \N__33054\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__33054\,
            I => \dron_frame_decoder_1.N_219_4\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__33051\,
            I => \dron_frame_decoder_1.N_219_4_cascade_\
        );

    \I__5490\ : InMux
    port map (
            O => \N__33048\,
            I => \N__33045\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__33042\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__33042\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_1_3\
        );

    \I__5487\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33036\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__33036\,
            I => \N__33033\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__33033\,
            I => \N__33030\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__33030\,
            I => scaler_4_data_5
        );

    \I__5483\ : CascadeMux
    port map (
            O => \N__33027\,
            I => \N__33023\
        );

    \I__5482\ : InMux
    port map (
            O => \N__33026\,
            I => \N__33020\
        );

    \I__5481\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33017\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__33020\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__33017\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__5478\ : CascadeMux
    port map (
            O => \N__33012\,
            I => \N__33008\
        );

    \I__5477\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33005\
        );

    \I__5476\ : InMux
    port map (
            O => \N__33008\,
            I => \N__33002\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__33005\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__33002\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__5473\ : CEMux
    port map (
            O => \N__32997\,
            I => \N__32993\
        );

    \I__5472\ : CEMux
    port map (
            O => \N__32996\,
            I => \N__32990\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__32993\,
            I => \uart_drone.data_rdyc_1_0\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__32990\,
            I => \uart_drone.data_rdyc_1_0\
        );

    \I__5469\ : SRMux
    port map (
            O => \N__32985\,
            I => \N__32982\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32978\
        );

    \I__5467\ : SRMux
    port map (
            O => \N__32981\,
            I => \N__32975\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__32978\,
            I => \N__32972\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32969\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__32972\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__5463\ : Odrv4
    port map (
            O => \N__32969\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__5462\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32961\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__32961\,
            I => \N__32958\
        );

    \I__5460\ : Odrv12
    port map (
            O => \N__32958\,
            I => \uart_drone.data_Auxce_0_0_4\
        );

    \I__5459\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32952\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__32952\,
            I => \dron_frame_decoder_1.N_263_5\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__32949\,
            I => \dron_frame_decoder_1.N_263_5_cascade_\
        );

    \I__5456\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32942\
        );

    \I__5455\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32938\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__32942\,
            I => \N__32935\
        );

    \I__5453\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32932\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__32938\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__32935\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__32932\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__5449\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__5447\ : Span4Mux_h
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__32916\,
            I => \uart_drone.data_Auxce_0_5\
        );

    \I__5445\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32910\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__32910\,
            I => \N__32907\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__32907\,
            I => \uart_drone.data_Auxce_0_6\
        );

    \I__5442\ : IoInMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__32901\,
            I => \N__32898\
        );

    \I__5440\ : IoSpan4Mux
    port map (
            O => \N__32898\,
            I => \N__32885\
        );

    \I__5439\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32882\
        );

    \I__5438\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32865\
        );

    \I__5437\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32865\
        );

    \I__5436\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32865\
        );

    \I__5435\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32865\
        );

    \I__5434\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32865\
        );

    \I__5433\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32865\
        );

    \I__5432\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32865\
        );

    \I__5431\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32865\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__32888\,
            I => \N__32861\
        );

    \I__5429\ : IoSpan4Mux
    port map (
            O => \N__32885\,
            I => \N__32856\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__32882\,
            I => \N__32851\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32851\
        );

    \I__5426\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32848\
        );

    \I__5425\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32843\
        );

    \I__5424\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32843\
        );

    \I__5423\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32840\
        );

    \I__5422\ : Span4Mux_s2_v
    port map (
            O => \N__32856\,
            I => \N__32835\
        );

    \I__5421\ : Span4Mux_v
    port map (
            O => \N__32851\,
            I => \N__32835\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__32848\,
            I => \N__32832\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__32843\,
            I => \debug_CH0_16A_c\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__32840\,
            I => \debug_CH0_16A_c\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__32835\,
            I => \debug_CH0_16A_c\
        );

    \I__5416\ : Odrv12
    port map (
            O => \N__32832\,
            I => \debug_CH0_16A_c\
        );

    \I__5415\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32807\
        );

    \I__5414\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32807\
        );

    \I__5413\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32807\
        );

    \I__5412\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32807\
        );

    \I__5411\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32798\
        );

    \I__5410\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32798\
        );

    \I__5409\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32798\
        );

    \I__5408\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32798\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32793\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__32798\,
            I => \N__32793\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__32793\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__5404\ : SRMux
    port map (
            O => \N__32790\,
            I => \N__32787\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32784\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__32781\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__32778\,
            I => \N__32774\
        );

    \I__5399\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32771\
        );

    \I__5398\ : InMux
    port map (
            O => \N__32774\,
            I => \N__32768\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__32771\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__32768\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__32763\,
            I => \N__32759\
        );

    \I__5394\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32756\
        );

    \I__5393\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32753\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__32756\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__32753\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__32748\,
            I => \N__32744\
        );

    \I__5389\ : InMux
    port map (
            O => \N__32747\,
            I => \N__32741\
        );

    \I__5388\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32738\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__32741\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__32738\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__32733\,
            I => \N__32729\
        );

    \I__5384\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32726\
        );

    \I__5383\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32723\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__32726\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__32723\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__32718\,
            I => \N__32715\
        );

    \I__5379\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32711\
        );

    \I__5378\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32708\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__32711\,
            I => \N__32705\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__32708\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__32705\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__32700\,
            I => \reset_module_System.reset6_3_cascade_\
        );

    \I__5373\ : InMux
    port map (
            O => \N__32697\,
            I => \N__32694\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__32694\,
            I => \reset_module_System.reset6_13\
        );

    \I__5371\ : CascadeMux
    port map (
            O => \N__32691\,
            I => \reset_module_System.reset6_17_cascade_\
        );

    \I__5370\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32679\
        );

    \I__5369\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32679\
        );

    \I__5368\ : InMux
    port map (
            O => \N__32686\,
            I => \N__32679\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__32679\,
            I => \reset_module_System.reset6_19\
        );

    \I__5366\ : InMux
    port map (
            O => \N__32676\,
            I => \N__32669\
        );

    \I__5365\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32669\
        );

    \I__5364\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32666\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__32669\,
            I => \reset_module_System.reset6_15\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__32666\,
            I => \reset_module_System.reset6_15\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__32661\,
            I => \reset_module_System.reset6_19_cascade_\
        );

    \I__5360\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32655\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__32655\,
            I => \uart_drone.data_Auxce_0_0_0\
        );

    \I__5358\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32649\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__32649\,
            I => \N__32646\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__32646\,
            I => \uart_drone.data_Auxce_0_0_2\
        );

    \I__5355\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32639\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__32642\,
            I => \N__32636\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__32639\,
            I => \N__32633\
        );

    \I__5352\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32630\
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__32633\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__32630\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__5349\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32621\
        );

    \I__5348\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32618\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__32621\,
            I => \uart_drone.N_126_li\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__32618\,
            I => \uart_drone.N_126_li\
        );

    \I__5345\ : CascadeMux
    port map (
            O => \N__32613\,
            I => \uart_drone.state_srsts_0_0_0_cascade_\
        );

    \I__5344\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32603\
        );

    \I__5343\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32599\
        );

    \I__5342\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32592\
        );

    \I__5341\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32592\
        );

    \I__5340\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32592\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__32603\,
            I => \N__32589\
        );

    \I__5338\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32586\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__32599\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__32592\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__32589\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__32586\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__5333\ : InMux
    port map (
            O => \N__32577\,
            I => \N__32571\
        );

    \I__5332\ : InMux
    port map (
            O => \N__32576\,
            I => \N__32571\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__32571\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__32568\,
            I => \N__32563\
        );

    \I__5329\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32560\
        );

    \I__5328\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32555\
        );

    \I__5327\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32555\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__32560\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__32555\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__5324\ : CascadeMux
    port map (
            O => \N__32550\,
            I => \reset_module_System.reset6_15_cascade_\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__32547\,
            I => \reset_module_System.count_1_1_cascade_\
        );

    \I__5322\ : InMux
    port map (
            O => \N__32544\,
            I => \N__32541\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__32541\,
            I => \N__32538\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__32538\,
            I => \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__32535\,
            I => \uart_drone.N_145_cascade_\
        );

    \I__5318\ : CascadeMux
    port map (
            O => \N__32532\,
            I => \uart_drone.un1_state_4_0_cascade_\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__32529\,
            I => \uart_drone.state_srsts_i_0_2_cascade_\
        );

    \I__5316\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32520\
        );

    \I__5315\ : InMux
    port map (
            O => \N__32525\,
            I => \N__32520\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__32520\,
            I => \N__32515\
        );

    \I__5313\ : InMux
    port map (
            O => \N__32519\,
            I => \N__32510\
        );

    \I__5312\ : InMux
    port map (
            O => \N__32518\,
            I => \N__32510\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__32515\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__32510\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__32505\,
            I => \N__32501\
        );

    \I__5308\ : InMux
    port map (
            O => \N__32504\,
            I => \N__32495\
        );

    \I__5307\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32495\
        );

    \I__5306\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32492\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__32495\,
            I => \N__32487\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__32492\,
            I => \N__32484\
        );

    \I__5303\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32481\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__32490\,
            I => \N__32478\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__32487\,
            I => \N__32475\
        );

    \I__5300\ : Span4Mux_h
    port map (
            O => \N__32484\,
            I => \N__32472\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__32481\,
            I => \N__32469\
        );

    \I__5298\ : InMux
    port map (
            O => \N__32478\,
            I => \N__32466\
        );

    \I__5297\ : Odrv4
    port map (
            O => \N__32475\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__32472\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__32469\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__32466\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__32457\,
            I => \pid_front.un1_pid_prereg_48_cascade_\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__5291\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32445\
        );

    \I__5290\ : InMux
    port map (
            O => \N__32450\,
            I => \N__32445\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__32445\,
            I => \pid_front.error_d_reg_prevZ0Z_19\
        );

    \I__5288\ : InMux
    port map (
            O => \N__32442\,
            I => \N__32436\
        );

    \I__5287\ : InMux
    port map (
            O => \N__32441\,
            I => \N__32436\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__32436\,
            I => \N__32433\
        );

    \I__5285\ : Span4Mux_v
    port map (
            O => \N__32433\,
            I => \N__32430\
        );

    \I__5284\ : Span4Mux_v
    port map (
            O => \N__32430\,
            I => \N__32427\
        );

    \I__5283\ : Sp12to4
    port map (
            O => \N__32427\,
            I => \N__32424\
        );

    \I__5282\ : Odrv12
    port map (
            O => \N__32424\,
            I => \pid_front.error_p_regZ0Z_19\
        );

    \I__5281\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32414\
        );

    \I__5279\ : InMux
    port map (
            O => \N__32417\,
            I => \N__32411\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__32414\,
            I => \pid_front.un1_pid_prereg_56\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__32411\,
            I => \pid_front.un1_pid_prereg_56\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__32406\,
            I => \pid_front.un1_pid_prereg_56_cascade_\
        );

    \I__5275\ : InMux
    port map (
            O => \N__32403\,
            I => \N__32400\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32396\
        );

    \I__5273\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32393\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__32396\,
            I => \pid_front.un1_pid_prereg_48\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__32393\,
            I => \pid_front.un1_pid_prereg_48\
        );

    \I__5270\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32385\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__32385\,
            I => \N__32382\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__32382\,
            I => \pid_front.N_1471_i\
        );

    \I__5267\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32372\
        );

    \I__5266\ : InMux
    port map (
            O => \N__32378\,
            I => \N__32372\
        );

    \I__5265\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32369\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__32372\,
            I => \N__32364\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32364\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__32364\,
            I => \pid_front.error_p_reg_esr_RNIA93NZ0Z_12\
        );

    \I__5261\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32352\
        );

    \I__5260\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32352\
        );

    \I__5259\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32352\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__32352\,
            I => \pid_front.error_d_reg_prevZ0Z_12\
        );

    \I__5257\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32344\
        );

    \I__5256\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32339\
        );

    \I__5255\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32339\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__32344\,
            I => \N__32334\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__32339\,
            I => \N__32334\
        );

    \I__5252\ : Span12Mux_v
    port map (
            O => \N__32334\,
            I => \N__32331\
        );

    \I__5251\ : Odrv12
    port map (
            O => \N__32331\,
            I => \pid_front.error_p_regZ0Z_12\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__32328\,
            I => \pid_front.un1_pid_prereg_107_0_cascade_\
        );

    \I__5249\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32322\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__32322\,
            I => drone_altitude_1
        );

    \I__5247\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32316\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__32316\,
            I => \N__32313\
        );

    \I__5245\ : Odrv12
    port map (
            O => \N__32313\,
            I => \pid_alt.error_axbZ0Z_1\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__32310\,
            I => \N__32306\
        );

    \I__5243\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32301\
        );

    \I__5242\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32296\
        );

    \I__5241\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32296\
        );

    \I__5240\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32293\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__32301\,
            I => \N__32288\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32288\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__32293\,
            I => \N__32285\
        );

    \I__5236\ : Span4Mux_v
    port map (
            O => \N__32288\,
            I => \N__32282\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__32285\,
            I => \N__32277\
        );

    \I__5234\ : Span4Mux_h
    port map (
            O => \N__32282\,
            I => \N__32277\
        );

    \I__5233\ : Span4Mux_h
    port map (
            O => \N__32277\,
            I => \N__32274\
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__32274\,
            I => \pid_front.error_p_regZ0Z_8\
        );

    \I__5231\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32268\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__32268\,
            I => \N__32263\
        );

    \I__5229\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32257\
        );

    \I__5228\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32257\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__32263\,
            I => \N__32254\
        );

    \I__5226\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32251\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__32257\,
            I => \N__32248\
        );

    \I__5224\ : Span4Mux_h
    port map (
            O => \N__32254\,
            I => \N__32243\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__32251\,
            I => \N__32243\
        );

    \I__5222\ : Span4Mux_v
    port map (
            O => \N__32248\,
            I => \N__32240\
        );

    \I__5221\ : Odrv4
    port map (
            O => \N__32243\,
            I => \pid_front.error_d_reg_prevZ0Z_8\
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__32240\,
            I => \pid_front.error_d_reg_prevZ0Z_8\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__32235\,
            I => \N__32232\
        );

    \I__5218\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32229\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__32229\,
            I => \pid_front.un1_pid_prereg_80_0\
        );

    \I__5216\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32223\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__32223\,
            I => \pid_front.N_1455_i\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__32220\,
            I => \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11_cascade_\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__32217\,
            I => \pid_front.un1_pid_prereg_57_cascade_\
        );

    \I__5212\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32209\
        );

    \I__5211\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32203\
        );

    \I__5210\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32200\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__32209\,
            I => \N__32197\
        );

    \I__5208\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32192\
        );

    \I__5207\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32192\
        );

    \I__5206\ : InMux
    port map (
            O => \N__32206\,
            I => \N__32189\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__32203\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__32200\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__32197\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__32192\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__32189\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__32178\,
            I => \N__32174\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__32177\,
            I => \N__32171\
        );

    \I__5198\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32167\
        );

    \I__5197\ : InMux
    port map (
            O => \N__32171\,
            I => \N__32164\
        );

    \I__5196\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32161\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__32167\,
            I => \N__32156\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__32164\,
            I => \N__32156\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__32161\,
            I => \N__32151\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__32156\,
            I => \N__32151\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__32151\,
            I => \dron_frame_decoder_1.stateZ0Z_7\
        );

    \I__5190\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32145\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__32145\,
            I => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\
        );

    \I__5188\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__32139\,
            I => \N__32136\
        );

    \I__5186\ : Odrv12
    port map (
            O => \N__32136\,
            I => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__32133\,
            I => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_\
        );

    \I__5184\ : InMux
    port map (
            O => \N__32130\,
            I => \N__32127\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__32127\,
            I => \dron_frame_decoder_1.drone_H_disp_side_9\
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__32124\,
            I => \dron_frame_decoder_1.N_198_cascade_\
        );

    \I__5181\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32118\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__32118\,
            I => \dron_frame_decoder_1.N_200\
        );

    \I__5179\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32112\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__32112\,
            I => \N__32108\
        );

    \I__5177\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32105\
        );

    \I__5176\ : Span4Mux_s3_h
    port map (
            O => \N__32108\,
            I => \N__32102\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32099\
        );

    \I__5174\ : Span4Mux_h
    port map (
            O => \N__32102\,
            I => \N__32096\
        );

    \I__5173\ : Span4Mux_s1_h
    port map (
            O => \N__32099\,
            I => \N__32093\
        );

    \I__5172\ : Span4Mux_h
    port map (
            O => \N__32096\,
            I => \N__32090\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__32093\,
            I => \N__32087\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__32090\,
            I => \N__32084\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__32087\,
            I => \N__32081\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__32084\,
            I => xy_kp_0
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__32081\,
            I => xy_kp_0
        );

    \I__5166\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32072\
        );

    \I__5165\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32069\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__32072\,
            I => \N__32066\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__32063\
        );

    \I__5162\ : Span4Mux_s2_h
    port map (
            O => \N__32066\,
            I => \N__32060\
        );

    \I__5161\ : Span12Mux_s4_h
    port map (
            O => \N__32063\,
            I => \N__32057\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__32060\,
            I => \N__32054\
        );

    \I__5159\ : Span12Mux_h
    port map (
            O => \N__32057\,
            I => \N__32051\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__32054\,
            I => \N__32048\
        );

    \I__5157\ : Odrv12
    port map (
            O => \N__32051\,
            I => xy_kp_1
        );

    \I__5156\ : Odrv4
    port map (
            O => \N__32048\,
            I => xy_kp_1
        );

    \I__5155\ : InMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__5153\ : Span4Mux_s3_h
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__5152\ : Span4Mux_h
    port map (
            O => \N__32034\,
            I => \N__32030\
        );

    \I__5151\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32027\
        );

    \I__5150\ : Span4Mux_h
    port map (
            O => \N__32030\,
            I => \N__32024\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__32021\
        );

    \I__5148\ : Span4Mux_h
    port map (
            O => \N__32024\,
            I => \N__32018\
        );

    \I__5147\ : Span12Mux_s9_h
    port map (
            O => \N__32021\,
            I => \N__32015\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__32018\,
            I => xy_kp_2
        );

    \I__5145\ : Odrv12
    port map (
            O => \N__32015\,
            I => xy_kp_2
        );

    \I__5144\ : InMux
    port map (
            O => \N__32010\,
            I => \N__32007\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__32007\,
            I => \N__32003\
        );

    \I__5142\ : InMux
    port map (
            O => \N__32006\,
            I => \N__32000\
        );

    \I__5141\ : Span4Mux_s3_h
    port map (
            O => \N__32003\,
            I => \N__31997\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__32000\,
            I => \N__31994\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__31997\,
            I => \N__31991\
        );

    \I__5138\ : Span4Mux_v
    port map (
            O => \N__31994\,
            I => \N__31988\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__31991\,
            I => \N__31985\
        );

    \I__5136\ : Span4Mux_h
    port map (
            O => \N__31988\,
            I => \N__31982\
        );

    \I__5135\ : Span4Mux_h
    port map (
            O => \N__31985\,
            I => \N__31979\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__31982\,
            I => \N__31976\
        );

    \I__5133\ : Odrv4
    port map (
            O => \N__31979\,
            I => xy_kp_3
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__31976\,
            I => xy_kp_3
        );

    \I__5131\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31968\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__31968\,
            I => \N__31964\
        );

    \I__5129\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31961\
        );

    \I__5128\ : Span4Mux_s3_h
    port map (
            O => \N__31964\,
            I => \N__31958\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31955\
        );

    \I__5126\ : Span4Mux_h
    port map (
            O => \N__31958\,
            I => \N__31952\
        );

    \I__5125\ : Span4Mux_s1_h
    port map (
            O => \N__31955\,
            I => \N__31949\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__31952\,
            I => \N__31946\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__31949\,
            I => \N__31943\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__31946\,
            I => \N__31940\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__31943\,
            I => \N__31937\
        );

    \I__5120\ : Odrv4
    port map (
            O => \N__31940\,
            I => xy_kp_7
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__31937\,
            I => xy_kp_7
        );

    \I__5118\ : CEMux
    port map (
            O => \N__31932\,
            I => \N__31929\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__31926\,
            I => \N__31922\
        );

    \I__5115\ : CEMux
    port map (
            O => \N__31925\,
            I => \N__31919\
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__31922\,
            I => \Commands_frame_decoder.state_RNIG48SZ0Z_7\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__31919\,
            I => \Commands_frame_decoder.state_RNIG48SZ0Z_7\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__31914\,
            I => \N__31910\
        );

    \I__5111\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31901\
        );

    \I__5110\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31901\
        );

    \I__5109\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31901\
        );

    \I__5108\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31898\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__31901\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__31898\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__5105\ : InMux
    port map (
            O => \N__31893\,
            I => \N__31890\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__31890\,
            I => \dron_frame_decoder_1.state_ns_i_a2_0_0_0\
        );

    \I__5103\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31880\
        );

    \I__5102\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31880\
        );

    \I__5101\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31877\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31874\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__31877\,
            I => \uart_drone.data_rdyc_1\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__31874\,
            I => \uart_drone.data_rdyc_1\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__31869\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__31866\,
            I => \N__31861\
        );

    \I__5095\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31858\
        );

    \I__5094\ : InMux
    port map (
            O => \N__31864\,
            I => \N__31853\
        );

    \I__5093\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31853\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__31858\,
            I => \N__31850\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__31853\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__31850\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__5089\ : InMux
    port map (
            O => \N__31845\,
            I => \N__31842\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__31842\,
            I => \N__31837\
        );

    \I__5087\ : InMux
    port map (
            O => \N__31841\,
            I => \N__31832\
        );

    \I__5086\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31832\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__31837\,
            I => \N__31826\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31826\
        );

    \I__5083\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31823\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__31826\,
            I => \Commands_frame_decoder.stateZ0Z_14\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__31823\,
            I => \Commands_frame_decoder.stateZ0Z_14\
        );

    \I__5080\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31815\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__31815\,
            I => \Commands_frame_decoder.count_1_sqmuxa\
        );

    \I__5078\ : InMux
    port map (
            O => \N__31812\,
            I => \N__31809\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__31809\,
            I => \N__31805\
        );

    \I__5076\ : InMux
    port map (
            O => \N__31808\,
            I => \N__31801\
        );

    \I__5075\ : Span4Mux_v
    port map (
            O => \N__31805\,
            I => \N__31798\
        );

    \I__5074\ : InMux
    port map (
            O => \N__31804\,
            I => \N__31795\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31790\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__31798\,
            I => \N__31790\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__31795\,
            I => \Commands_frame_decoder.stateZ0Z_13\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__31790\,
            I => \Commands_frame_decoder.stateZ0Z_13\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__31785\,
            I => \N__31768\
        );

    \I__5068\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31759\
        );

    \I__5067\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31754\
        );

    \I__5066\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31754\
        );

    \I__5065\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31747\
        );

    \I__5064\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31747\
        );

    \I__5063\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31747\
        );

    \I__5062\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31742\
        );

    \I__5061\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31742\
        );

    \I__5060\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31735\
        );

    \I__5059\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31732\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__31774\,
            I => \N__31729\
        );

    \I__5057\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31722\
        );

    \I__5056\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31719\
        );

    \I__5055\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31716\
        );

    \I__5054\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31713\
        );

    \I__5053\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31704\
        );

    \I__5052\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31704\
        );

    \I__5051\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31704\
        );

    \I__5050\ : InMux
    port map (
            O => \N__31764\,
            I => \N__31704\
        );

    \I__5049\ : InMux
    port map (
            O => \N__31763\,
            I => \N__31701\
        );

    \I__5048\ : InMux
    port map (
            O => \N__31762\,
            I => \N__31698\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__31759\,
            I => \N__31695\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__31754\,
            I => \N__31690\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__31747\,
            I => \N__31690\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__31742\,
            I => \N__31687\
        );

    \I__5043\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31680\
        );

    \I__5042\ : InMux
    port map (
            O => \N__31740\,
            I => \N__31680\
        );

    \I__5041\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31680\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__31738\,
            I => \N__31675\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__31735\,
            I => \N__31671\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__31732\,
            I => \N__31668\
        );

    \I__5037\ : InMux
    port map (
            O => \N__31729\,
            I => \N__31663\
        );

    \I__5036\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31663\
        );

    \I__5035\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31656\
        );

    \I__5034\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31656\
        );

    \I__5033\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31656\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31650\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__31719\,
            I => \N__31650\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__31716\,
            I => \N__31647\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__31713\,
            I => \N__31634\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31634\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__31701\,
            I => \N__31634\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__31698\,
            I => \N__31634\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__31695\,
            I => \N__31634\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__31690\,
            I => \N__31634\
        );

    \I__5023\ : Span4Mux_h
    port map (
            O => \N__31687\,
            I => \N__31629\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__31680\,
            I => \N__31629\
        );

    \I__5021\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31626\
        );

    \I__5020\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31621\
        );

    \I__5019\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31621\
        );

    \I__5018\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31618\
        );

    \I__5017\ : Span4Mux_v
    port map (
            O => \N__31671\,
            I => \N__31613\
        );

    \I__5016\ : Span4Mux_v
    port map (
            O => \N__31668\,
            I => \N__31613\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__31663\,
            I => \N__31608\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__31656\,
            I => \N__31608\
        );

    \I__5013\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31605\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__31650\,
            I => \N__31596\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__31647\,
            I => \N__31596\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__31634\,
            I => \N__31596\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__31629\,
            I => \N__31596\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__31626\,
            I => uart_pc_data_rdy
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__31621\,
            I => uart_pc_data_rdy
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__31618\,
            I => uart_pc_data_rdy
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__31613\,
            I => uart_pc_data_rdy
        );

    \I__5004\ : Odrv12
    port map (
            O => \N__31608\,
            I => uart_pc_data_rdy
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__31605\,
            I => uart_pc_data_rdy
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__31596\,
            I => uart_pc_data_rdy
        );

    \I__5001\ : CascadeMux
    port map (
            O => \N__31581\,
            I => \dron_frame_decoder_1.state_ns_0_a3_0_1Z0Z_1_cascade_\
        );

    \I__5000\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31575\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__31575\,
            I => \dron_frame_decoder_1.N_220\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__31572\,
            I => \dron_frame_decoder_1.N_220_cascade_\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__31569\,
            I => \N__31566\
        );

    \I__4996\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31560\
        );

    \I__4995\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31560\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__31560\,
            I => \dron_frame_decoder_1.N_224\
        );

    \I__4993\ : InMux
    port map (
            O => \N__31557\,
            I => \N__31553\
        );

    \I__4992\ : InMux
    port map (
            O => \N__31556\,
            I => \N__31550\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__31553\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__31550\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__31545\,
            I => \N__31540\
        );

    \I__4988\ : InMux
    port map (
            O => \N__31544\,
            I => \N__31534\
        );

    \I__4987\ : InMux
    port map (
            O => \N__31543\,
            I => \N__31534\
        );

    \I__4986\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31529\
        );

    \I__4985\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31529\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__31534\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__31529\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__31524\,
            I => \N__31521\
        );

    \I__4981\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31518\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__31518\,
            I => \N__31515\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__31515\,
            I => \uart_drone.un1_state_2_0_a3_0\
        );

    \I__4978\ : InMux
    port map (
            O => \N__31512\,
            I => \uart_drone.un4_timer_Count_1_cry_1\
        );

    \I__4977\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__31506\,
            I => \uart_drone.timer_Count_RNO_0_0_3\
        );

    \I__4975\ : InMux
    port map (
            O => \N__31503\,
            I => \uart_drone.un4_timer_Count_1_cry_2\
        );

    \I__4974\ : InMux
    port map (
            O => \N__31500\,
            I => \uart_drone.un4_timer_Count_1_cry_3\
        );

    \I__4973\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31494\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__31494\,
            I => \uart_drone.timer_Count_RNO_0_0_4\
        );

    \I__4971\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31488\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__31488\,
            I => \uart_drone.timer_Count_RNO_0_0_2\
        );

    \I__4969\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31478\
        );

    \I__4968\ : InMux
    port map (
            O => \N__31484\,
            I => \N__31475\
        );

    \I__4967\ : InMux
    port map (
            O => \N__31483\,
            I => \N__31472\
        );

    \I__4966\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31467\
        );

    \I__4965\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31467\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__31478\,
            I => \uart_drone.N_143\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__31475\,
            I => \uart_drone.N_143\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__31472\,
            I => \uart_drone.N_143\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__31467\,
            I => \uart_drone.N_143\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__31458\,
            I => \N__31454\
        );

    \I__4959\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31450\
        );

    \I__4958\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31445\
        );

    \I__4957\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31445\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__31450\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__31445\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__4954\ : InMux
    port map (
            O => \N__31440\,
            I => \N__31437\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__31437\,
            I => \N__31432\
        );

    \I__4952\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31429\
        );

    \I__4951\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31426\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__31432\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__31429\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__31426\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__4947\ : InMux
    port map (
            O => \N__31419\,
            I => \N__31415\
        );

    \I__4946\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31412\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__31415\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__31412\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4943\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31402\
        );

    \I__4942\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31397\
        );

    \I__4941\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31397\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__31402\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__31397\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__4938\ : CascadeMux
    port map (
            O => \N__31392\,
            I => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4_cascade_\
        );

    \I__4937\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31386\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__31386\,
            I => \Commands_frame_decoder.WDT8lto15_N_5L7_1\
        );

    \I__4935\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31380\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__31380\,
            I => \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12\
        );

    \I__4933\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31372\
        );

    \I__4932\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31369\
        );

    \I__4931\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31366\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__31372\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__31369\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__31366\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4927\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31353\
        );

    \I__4926\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31350\
        );

    \I__4925\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31345\
        );

    \I__4924\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31345\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__31353\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__31350\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__31345\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__31338\,
            I => \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12_cascade_\
        );

    \I__4919\ : InMux
    port map (
            O => \N__31335\,
            I => \N__31330\
        );

    \I__4918\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31327\
        );

    \I__4917\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31324\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__31330\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__31327\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__31324\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4913\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31310\
        );

    \I__4912\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31300\
        );

    \I__4911\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31297\
        );

    \I__4910\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31292\
        );

    \I__4909\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31292\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__31310\,
            I => \N__31287\
        );

    \I__4907\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31280\
        );

    \I__4906\ : InMux
    port map (
            O => \N__31308\,
            I => \N__31280\
        );

    \I__4905\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31280\
        );

    \I__4904\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31275\
        );

    \I__4903\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31275\
        );

    \I__4902\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31270\
        );

    \I__4901\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31270\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__31300\,
            I => \N__31264\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31264\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__31292\,
            I => \N__31261\
        );

    \I__4897\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31256\
        );

    \I__4896\ : InMux
    port map (
            O => \N__31290\,
            I => \N__31256\
        );

    \I__4895\ : Span4Mux_v
    port map (
            O => \N__31287\,
            I => \N__31253\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__31280\,
            I => \N__31248\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31248\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__31270\,
            I => \N__31245\
        );

    \I__4891\ : InMux
    port map (
            O => \N__31269\,
            I => \N__31242\
        );

    \I__4890\ : Span4Mux_v
    port map (
            O => \N__31264\,
            I => \N__31239\
        );

    \I__4889\ : Span4Mux_v
    port map (
            O => \N__31261\,
            I => \N__31234\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__31256\,
            I => \N__31234\
        );

    \I__4887\ : Span4Mux_h
    port map (
            O => \N__31253\,
            I => \N__31225\
        );

    \I__4886\ : Span4Mux_v
    port map (
            O => \N__31248\,
            I => \N__31225\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__31245\,
            I => \N__31225\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__31242\,
            I => \N__31225\
        );

    \I__4883\ : Span4Mux_h
    port map (
            O => \N__31239\,
            I => \N__31222\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__31234\,
            I => \N__31219\
        );

    \I__4881\ : Span4Mux_v
    port map (
            O => \N__31225\,
            I => \N__31216\
        );

    \I__4880\ : Odrv4
    port map (
            O => \N__31222\,
            I => \Commands_frame_decoder.WDT8_0\
        );

    \I__4879\ : Odrv4
    port map (
            O => \N__31219\,
            I => \Commands_frame_decoder.WDT8_0\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__31216\,
            I => \Commands_frame_decoder.WDT8_0\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__31209\,
            I => \uart_drone.N_126_li_cascade_\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__31206\,
            I => \uart_drone.N_143_cascade_\
        );

    \I__4875\ : IoInMux
    port map (
            O => \N__31203\,
            I => \N__31200\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31197\
        );

    \I__4873\ : Span4Mux_s3_v
    port map (
            O => \N__31197\,
            I => \N__31194\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__31194\,
            I => \pid_front.state_0_0\
        );

    \I__4871\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31188\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__31188\,
            I => uart_input_pc_c
        );

    \I__4869\ : InMux
    port map (
            O => \N__31185\,
            I => \N__31182\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31179\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__31179\,
            I => \uart_pc_sync.aux_0__0_Z0Z_0\
        );

    \I__4866\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31173\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__31173\,
            I => \N__31170\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__31170\,
            I => \uart_drone_sync.aux_3__0__0_0\
        );

    \I__4863\ : CascadeMux
    port map (
            O => \N__31167\,
            I => \Commands_frame_decoder.state_0_sqmuxa_1_cascade_\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__31164\,
            I => \N__31160\
        );

    \I__4861\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31157\
        );

    \I__4860\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31154\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__31157\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__31154\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__4857\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31146\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__31146\,
            I => \N__31143\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__31143\,
            I => \uart_pc_sync.aux_1__0_Z0Z_0\
        );

    \I__4854\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__31134\,
            I => \uart_pc_sync.aux_2__0_Z0Z_0\
        );

    \I__4851\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31127\
        );

    \I__4850\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31124\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__31127\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__31124\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__4847\ : CascadeMux
    port map (
            O => \N__31119\,
            I => \N__31115\
        );

    \I__4846\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31112\
        );

    \I__4845\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31109\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__31112\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__31109\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4842\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31100\
        );

    \I__4841\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31097\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__31100\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__31097\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__4838\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31088\
        );

    \I__4837\ : InMux
    port map (
            O => \N__31091\,
            I => \N__31085\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__31088\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__31085\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__4834\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31076\
        );

    \I__4833\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31073\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__31076\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__31073\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__31068\,
            I => \N__31064\
        );

    \I__4829\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31061\
        );

    \I__4828\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31058\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__31061\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__31058\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__4825\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31049\
        );

    \I__4824\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31046\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__31049\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__31046\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__31041\,
            I => \pid_front.un1_pid_prereg_23_cascade_\
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__31038\,
            I => \pid_front.un1_pid_prereg_30_cascade_\
        );

    \I__4819\ : InMux
    port map (
            O => \N__31035\,
            I => \N__31029\
        );

    \I__4818\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31029\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__31026\,
            I => \N__31023\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__4814\ : Span4Mux_h
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__31017\,
            I => \pid_front.error_p_regZ0Z_15\
        );

    \I__4812\ : CascadeMux
    port map (
            O => \N__31014\,
            I => \N__31011\
        );

    \I__4811\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31005\
        );

    \I__4810\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31005\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__31005\,
            I => \pid_front.error_d_reg_prevZ0Z_15\
        );

    \I__4808\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30998\
        );

    \I__4807\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30995\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__30998\,
            I => \pid_front.un1_pid_prereg_29\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__30995\,
            I => \pid_front.un1_pid_prereg_29\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__30990\,
            I => \pid_front.un1_pid_prereg_29_cascade_\
        );

    \I__4803\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30983\
        );

    \I__4802\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30980\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__30983\,
            I => \N__30975\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__30980\,
            I => \N__30975\
        );

    \I__4799\ : Span4Mux_v
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__4798\ : Span4Mux_h
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__4797\ : Span4Mux_v
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__30966\,
            I => \pid_front.error_p_regZ0Z_14\
        );

    \I__4795\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30956\
        );

    \I__4794\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30956\
        );

    \I__4793\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30953\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__30956\,
            I => \pid_front.un1_pid_prereg_24\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__30953\,
            I => \pid_front.un1_pid_prereg_24\
        );

    \I__4790\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30945\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__30942\,
            I => \N__30939\
        );

    \I__4787\ : Span4Mux_h
    port map (
            O => \N__30939\,
            I => \N__30936\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__30936\,
            I => \N__30933\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__30933\,
            I => \pid_front.O_0_11\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__30930\,
            I => \pid_front.N_1451_i_cascade_\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__30927\,
            I => \pid_front.error_d_reg_esr_RNINKUFZ0Z_7_cascade_\
        );

    \I__4782\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__30921\,
            I => \pid_front.un1_pid_prereg_70_0\
        );

    \I__4780\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30914\
        );

    \I__4779\ : InMux
    port map (
            O => \N__30917\,
            I => \N__30911\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__30914\,
            I => \N__30908\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__30911\,
            I => \pid_front.un1_pid_prereg_23\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__30908\,
            I => \pid_front.un1_pid_prereg_23\
        );

    \I__4775\ : InMux
    port map (
            O => \N__30903\,
            I => \N__30900\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__30900\,
            I => \dron_frame_decoder_1.drone_altitude_5\
        );

    \I__4773\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__30894\,
            I => \dron_frame_decoder_1.drone_altitude_6\
        );

    \I__4771\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__30888\,
            I => \dron_frame_decoder_1.drone_altitude_7\
        );

    \I__4769\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30882\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__30882\,
            I => \dron_frame_decoder_1.drone_altitude_8\
        );

    \I__4767\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30876\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__30876\,
            I => drone_altitude_14
        );

    \I__4765\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30870\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__30870\,
            I => drone_altitude_13
        );

    \I__4763\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__30864\,
            I => drone_altitude_12
        );

    \I__4761\ : CEMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30855\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__30855\,
            I => \N__30851\
        );

    \I__4758\ : CEMux
    port map (
            O => \N__30854\,
            I => \N__30847\
        );

    \I__4757\ : Span4Mux_h
    port map (
            O => \N__30851\,
            I => \N__30844\
        );

    \I__4756\ : CEMux
    port map (
            O => \N__30850\,
            I => \N__30841\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__30847\,
            I => \N__30838\
        );

    \I__4754\ : Sp12to4
    port map (
            O => \N__30844\,
            I => \N__30833\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__30841\,
            I => \N__30833\
        );

    \I__4752\ : Sp12to4
    port map (
            O => \N__30838\,
            I => \N__30830\
        );

    \I__4751\ : Odrv12
    port map (
            O => \N__30833\,
            I => \dron_frame_decoder_1.N_513_0\
        );

    \I__4750\ : Odrv12
    port map (
            O => \N__30830\,
            I => \dron_frame_decoder_1.N_513_0\
        );

    \I__4749\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30820\
        );

    \I__4748\ : InMux
    port map (
            O => \N__30824\,
            I => \N__30815\
        );

    \I__4747\ : InMux
    port map (
            O => \N__30823\,
            I => \N__30815\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30812\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__30815\,
            I => \N__30809\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__30812\,
            I => \N__30806\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__30809\,
            I => \N__30803\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__30806\,
            I => \N__30800\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__30803\,
            I => \N__30797\
        );

    \I__4740\ : Span4Mux_h
    port map (
            O => \N__30800\,
            I => \N__30794\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__30797\,
            I => \pid_front.error_p_regZ0Z_9\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__30794\,
            I => \pid_front.error_p_regZ0Z_9\
        );

    \I__4737\ : InMux
    port map (
            O => \N__30789\,
            I => \N__30782\
        );

    \I__4736\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30782\
        );

    \I__4735\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30779\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__30782\,
            I => \pid_front.error_d_reg_prevZ0Z_9\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__30779\,
            I => \pid_front.error_d_reg_prevZ0Z_9\
        );

    \I__4732\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30771\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__30771\,
            I => \N__30768\
        );

    \I__4730\ : Span4Mux_v
    port map (
            O => \N__30768\,
            I => \N__30765\
        );

    \I__4729\ : Odrv4
    port map (
            O => \N__30765\,
            I => \pid_front.N_1459_i\
        );

    \I__4728\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30759\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__30759\,
            I => \N__30755\
        );

    \I__4726\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30752\
        );

    \I__4725\ : Span4Mux_v
    port map (
            O => \N__30755\,
            I => \N__30749\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__30752\,
            I => \N__30746\
        );

    \I__4723\ : Sp12to4
    port map (
            O => \N__30749\,
            I => \N__30743\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__30746\,
            I => \N__30740\
        );

    \I__4721\ : Span12Mux_s11_h
    port map (
            O => \N__30743\,
            I => \N__30737\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__30740\,
            I => \N__30734\
        );

    \I__4719\ : Odrv12
    port map (
            O => \N__30737\,
            I => xy_kp_6
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__30734\,
            I => xy_kp_6
        );

    \I__4717\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__30723\,
            I => \N__30719\
        );

    \I__4714\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30716\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__30719\,
            I => \N__30713\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__30716\,
            I => \N__30710\
        );

    \I__4711\ : Span4Mux_h
    port map (
            O => \N__30713\,
            I => \N__30707\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__30710\,
            I => \N__30704\
        );

    \I__4709\ : Sp12to4
    port map (
            O => \N__30707\,
            I => \N__30701\
        );

    \I__4708\ : Span4Mux_h
    port map (
            O => \N__30704\,
            I => \N__30698\
        );

    \I__4707\ : Odrv12
    port map (
            O => \N__30701\,
            I => xy_kp_5
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__30698\,
            I => xy_kp_5
        );

    \I__4705\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30690\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__4703\ : Span4Mux_v
    port map (
            O => \N__30687\,
            I => \N__30682\
        );

    \I__4702\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30679\
        );

    \I__4701\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30676\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__30682\,
            I => \N__30671\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__30679\,
            I => \N__30671\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30668\
        );

    \I__4697\ : Span4Mux_h
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__30668\,
            I => \N__30662\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__30665\,
            I => \N__30659\
        );

    \I__4694\ : Sp12to4
    port map (
            O => \N__30662\,
            I => \N__30656\
        );

    \I__4693\ : Sp12to4
    port map (
            O => \N__30659\,
            I => \N__30650\
        );

    \I__4692\ : Span12Mux_s8_h
    port map (
            O => \N__30656\,
            I => \N__30650\
        );

    \I__4691\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30647\
        );

    \I__4690\ : Odrv12
    port map (
            O => \N__30650\,
            I => drone_altitude_0
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__30647\,
            I => drone_altitude_0
        );

    \I__4688\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__30639\,
            I => \dron_frame_decoder_1.drone_altitude_4\
        );

    \I__4686\ : CascadeMux
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__4685\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__30630\,
            I => \uart_pc.data_Auxce_0_5\
        );

    \I__4683\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30624\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__30624\,
            I => \uart_pc.data_Auxce_0_6\
        );

    \I__4681\ : InMux
    port map (
            O => \N__30621\,
            I => \N__30615\
        );

    \I__4680\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30612\
        );

    \I__4679\ : InMux
    port map (
            O => \N__30619\,
            I => \N__30609\
        );

    \I__4678\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30606\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__30615\,
            I => \N__30603\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__30612\,
            I => \N__30598\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__30609\,
            I => \N__30598\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__30606\,
            I => \uart_pc.N_152\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__30603\,
            I => \uart_pc.N_152\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__30598\,
            I => \uart_pc.N_152\
        );

    \I__4671\ : InMux
    port map (
            O => \N__30591\,
            I => \N__30588\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__30588\,
            I => \N__30585\
        );

    \I__4669\ : Odrv4
    port map (
            O => \N__30585\,
            I => \uart_pc.data_Auxce_0_0_0\
        );

    \I__4668\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30579\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__30579\,
            I => \N__30576\
        );

    \I__4666\ : Odrv4
    port map (
            O => \N__30576\,
            I => \uart_pc.data_Auxce_0_1\
        );

    \I__4665\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30570\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__30570\,
            I => \N__30567\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__30567\,
            I => \uart_pc.data_Auxce_0_0_2\
        );

    \I__4662\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30553\
        );

    \I__4661\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30546\
        );

    \I__4660\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30546\
        );

    \I__4659\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30546\
        );

    \I__4658\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30535\
        );

    \I__4657\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30535\
        );

    \I__4656\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30535\
        );

    \I__4655\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30535\
        );

    \I__4654\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30535\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__30553\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__30546\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__30535\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__4650\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30505\
        );

    \I__4649\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30505\
        );

    \I__4648\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30505\
        );

    \I__4647\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30505\
        );

    \I__4646\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30505\
        );

    \I__4645\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30505\
        );

    \I__4644\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30494\
        );

    \I__4643\ : InMux
    port map (
            O => \N__30521\,
            I => \N__30494\
        );

    \I__4642\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30494\
        );

    \I__4641\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30494\
        );

    \I__4640\ : InMux
    port map (
            O => \N__30518\,
            I => \N__30494\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__30505\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__30494\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__30489\,
            I => \N__30482\
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__30488\,
            I => \N__30478\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__30487\,
            I => \N__30473\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__30486\,
            I => \N__30469\
        );

    \I__4633\ : InMux
    port map (
            O => \N__30485\,
            I => \N__30457\
        );

    \I__4632\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30457\
        );

    \I__4631\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30457\
        );

    \I__4630\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30457\
        );

    \I__4629\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30457\
        );

    \I__4628\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30446\
        );

    \I__4627\ : InMux
    port map (
            O => \N__30473\,
            I => \N__30446\
        );

    \I__4626\ : InMux
    port map (
            O => \N__30472\,
            I => \N__30446\
        );

    \I__4625\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30446\
        );

    \I__4624\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30446\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__30457\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__30446\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__4620\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30435\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__30435\,
            I => \N__30432\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__30432\,
            I => \uart_pc.data_Auxce_0_3\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__30429\,
            I => \N__30426\
        );

    \I__4616\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30423\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__30423\,
            I => \N__30419\
        );

    \I__4614\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30416\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__30419\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__30416\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__4611\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__30408\,
            I => \N__30404\
        );

    \I__4609\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30401\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__30404\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__30401\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__4606\ : CascadeMux
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__4605\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30389\
        );

    \I__4604\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30386\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__30389\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__30386\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__4601\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30357\
        );

    \I__4600\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30357\
        );

    \I__4599\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30357\
        );

    \I__4598\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30357\
        );

    \I__4597\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30357\
        );

    \I__4596\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30357\
        );

    \I__4595\ : InMux
    port map (
            O => \N__30375\,
            I => \N__30357\
        );

    \I__4594\ : InMux
    port map (
            O => \N__30374\,
            I => \N__30357\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__30357\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__4592\ : IoInMux
    port map (
            O => \N__30354\,
            I => \N__30351\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__30351\,
            I => \N__30348\
        );

    \I__4590\ : Span4Mux_s3_v
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__30345\,
            I => \N__30341\
        );

    \I__4588\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30330\
        );

    \I__4587\ : Span4Mux_h
    port map (
            O => \N__30341\,
            I => \N__30323\
        );

    \I__4586\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30314\
        );

    \I__4585\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30314\
        );

    \I__4584\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30314\
        );

    \I__4583\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30314\
        );

    \I__4582\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30305\
        );

    \I__4581\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30305\
        );

    \I__4580\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30305\
        );

    \I__4579\ : InMux
    port map (
            O => \N__30333\,
            I => \N__30305\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__30330\,
            I => \N__30302\
        );

    \I__4577\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30295\
        );

    \I__4576\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30295\
        );

    \I__4575\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30295\
        );

    \I__4574\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30292\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__30323\,
            I => \debug_CH2_18A_c\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__30314\,
            I => \debug_CH2_18A_c\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__30305\,
            I => \debug_CH2_18A_c\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__30302\,
            I => \debug_CH2_18A_c\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__30295\,
            I => \debug_CH2_18A_c\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__30292\,
            I => \debug_CH2_18A_c\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__30279\,
            I => \N__30275\
        );

    \I__4566\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30272\
        );

    \I__4565\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30269\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__30272\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__30269\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__4562\ : SRMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__30261\,
            I => \N__30258\
        );

    \I__4560\ : Span4Mux_h
    port map (
            O => \N__30258\,
            I => \N__30255\
        );

    \I__4559\ : Span4Mux_h
    port map (
            O => \N__30255\,
            I => \N__30252\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__30252\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__4557\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30245\
        );

    \I__4556\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30242\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__30245\,
            I => \N__30239\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__30242\,
            I => \N__30230\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__30239\,
            I => \N__30227\
        );

    \I__4552\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30224\
        );

    \I__4551\ : InMux
    port map (
            O => \N__30237\,
            I => \N__30219\
        );

    \I__4550\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30219\
        );

    \I__4549\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30212\
        );

    \I__4548\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30212\
        );

    \I__4547\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30212\
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__30230\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__30227\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__30224\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__30219\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__30212\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__30201\,
            I => \uart_pc.CO0_cascade_\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__30198\,
            I => \N__30194\
        );

    \I__4539\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30186\
        );

    \I__4538\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30186\
        );

    \I__4537\ : InMux
    port map (
            O => \N__30193\,
            I => \N__30186\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__30186\,
            I => \N__30183\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__30183\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__4534\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30174\
        );

    \I__4533\ : InMux
    port map (
            O => \N__30179\,
            I => \N__30174\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__30174\,
            I => \N__30171\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__30171\,
            I => \uart_pc.un1_state_7_0\
        );

    \I__4530\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30165\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__30165\,
            I => \N__30162\
        );

    \I__4528\ : Odrv12
    port map (
            O => \N__30162\,
            I => \uart_pc.data_Auxce_0_0_4\
        );

    \I__4527\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__30156\,
            I => \uart_pc.N_144_1\
        );

    \I__4525\ : CascadeMux
    port map (
            O => \N__30153\,
            I => \uart_pc.N_145_cascade_\
        );

    \I__4524\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30145\
        );

    \I__4523\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30141\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__30148\,
            I => \N__30138\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__30145\,
            I => \N__30135\
        );

    \I__4520\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30132\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__30141\,
            I => \N__30129\
        );

    \I__4518\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30126\
        );

    \I__4517\ : Odrv12
    port map (
            O => \N__30135\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__30132\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__30129\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__30126\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__4513\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__30114\,
            I => \uart_pc_sync.aux_3__0_Z0Z_0\
        );

    \I__4511\ : CascadeMux
    port map (
            O => \N__30111\,
            I => \uart_drone.timer_Count_RNO_0_0_1_cascade_\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__30108\,
            I => \N__30104\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__30107\,
            I => \N__30101\
        );

    \I__4508\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30098\
        );

    \I__4507\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30095\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__30098\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__30095\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__4504\ : CascadeMux
    port map (
            O => \N__30090\,
            I => \N__30086\
        );

    \I__4503\ : InMux
    port map (
            O => \N__30089\,
            I => \N__30083\
        );

    \I__4502\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30080\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__30083\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__30080\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__30075\,
            I => \N__30071\
        );

    \I__4498\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30068\
        );

    \I__4497\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30065\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__30068\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__30065\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__4494\ : CascadeMux
    port map (
            O => \N__30060\,
            I => \N__30057\
        );

    \I__4493\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30053\
        );

    \I__4492\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30050\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__30053\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__30050\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__30045\,
            I => \N__30040\
        );

    \I__4488\ : InMux
    port map (
            O => \N__30044\,
            I => \N__30033\
        );

    \I__4487\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30033\
        );

    \I__4486\ : InMux
    port map (
            O => \N__30040\,
            I => \N__30033\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__30033\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__4484\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30026\
        );

    \I__4483\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30023\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__30026\,
            I => \uart_pc.N_126_li\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__30023\,
            I => \uart_pc.N_126_li\
        );

    \I__4480\ : CascadeMux
    port map (
            O => \N__30018\,
            I => \uart_pc.state_srsts_0_0_0_cascade_\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__30015\,
            I => \N__30012\
        );

    \I__4478\ : InMux
    port map (
            O => \N__30012\,
            I => \N__30006\
        );

    \I__4477\ : InMux
    port map (
            O => \N__30011\,
            I => \N__30006\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__30006\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__30003\,
            I => \N__30000\
        );

    \I__4474\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29993\
        );

    \I__4473\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29993\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__29998\,
            I => \N__29988\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__29993\,
            I => \N__29985\
        );

    \I__4470\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29978\
        );

    \I__4469\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29978\
        );

    \I__4468\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29978\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__29985\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__29978\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4465\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29969\
        );

    \I__4464\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29962\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__29969\,
            I => \N__29959\
        );

    \I__4462\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29956\
        );

    \I__4461\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29949\
        );

    \I__4460\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29949\
        );

    \I__4459\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29949\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__29962\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__29959\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__29956\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__29949\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__4454\ : CascadeMux
    port map (
            O => \N__29940\,
            I => \uart_pc.un1_state_4_0_cascade_\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__29937\,
            I => \N__29927\
        );

    \I__4452\ : InMux
    port map (
            O => \N__29936\,
            I => \N__29920\
        );

    \I__4451\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29920\
        );

    \I__4450\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29920\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__29933\,
            I => \N__29916\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__29932\,
            I => \N__29913\
        );

    \I__4447\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29906\
        );

    \I__4446\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29906\
        );

    \I__4445\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29906\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__29920\,
            I => \N__29903\
        );

    \I__4443\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29900\
        );

    \I__4442\ : InMux
    port map (
            O => \N__29916\,
            I => \N__29895\
        );

    \I__4441\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29895\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__29906\,
            I => \N__29892\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__29903\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__29900\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__29895\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__29892\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4435\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29871\
        );

    \I__4434\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29871\
        );

    \I__4433\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29868\
        );

    \I__4432\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29863\
        );

    \I__4431\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29863\
        );

    \I__4430\ : InMux
    port map (
            O => \N__29878\,
            I => \N__29856\
        );

    \I__4429\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29856\
        );

    \I__4428\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29856\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__29871\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__29868\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__29863\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__29856\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4423\ : InMux
    port map (
            O => \N__29847\,
            I => \bfn_8_6_0_\
        );

    \I__4422\ : InMux
    port map (
            O => \N__29844\,
            I => \Commands_frame_decoder.un1_WDT_cry_8\
        );

    \I__4421\ : InMux
    port map (
            O => \N__29841\,
            I => \Commands_frame_decoder.un1_WDT_cry_9\
        );

    \I__4420\ : InMux
    port map (
            O => \N__29838\,
            I => \Commands_frame_decoder.un1_WDT_cry_10\
        );

    \I__4419\ : InMux
    port map (
            O => \N__29835\,
            I => \Commands_frame_decoder.un1_WDT_cry_11\
        );

    \I__4418\ : InMux
    port map (
            O => \N__29832\,
            I => \Commands_frame_decoder.un1_WDT_cry_12\
        );

    \I__4417\ : InMux
    port map (
            O => \N__29829\,
            I => \Commands_frame_decoder.un1_WDT_cry_13\
        );

    \I__4416\ : InMux
    port map (
            O => \N__29826\,
            I => \Commands_frame_decoder.un1_WDT_cry_14\
        );

    \I__4415\ : SRMux
    port map (
            O => \N__29823\,
            I => \N__29820\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29816\
        );

    \I__4413\ : SRMux
    port map (
            O => \N__29819\,
            I => \N__29813\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__29816\,
            I => \N__29808\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__29813\,
            I => \N__29808\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__29808\,
            I => \N__29805\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__29805\,
            I => \Commands_frame_decoder.un1_state57_iZ0\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__29802\,
            I => \uart_pc.state_srsts_i_0_2_cascade_\
        );

    \I__4407\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29796\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__29796\,
            I => \Commands_frame_decoder.WDTZ0Z_0\
        );

    \I__4405\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__29790\,
            I => \Commands_frame_decoder.WDTZ0Z_1\
        );

    \I__4403\ : InMux
    port map (
            O => \N__29787\,
            I => \Commands_frame_decoder.un1_WDT_cry_0\
        );

    \I__4402\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__29781\,
            I => \Commands_frame_decoder.WDTZ0Z_2\
        );

    \I__4400\ : InMux
    port map (
            O => \N__29778\,
            I => \Commands_frame_decoder.un1_WDT_cry_1\
        );

    \I__4399\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29772\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__29772\,
            I => \Commands_frame_decoder.WDTZ0Z_3\
        );

    \I__4397\ : InMux
    port map (
            O => \N__29769\,
            I => \Commands_frame_decoder.un1_WDT_cry_2\
        );

    \I__4396\ : InMux
    port map (
            O => \N__29766\,
            I => \Commands_frame_decoder.un1_WDT_cry_3\
        );

    \I__4395\ : InMux
    port map (
            O => \N__29763\,
            I => \Commands_frame_decoder.un1_WDT_cry_4\
        );

    \I__4394\ : InMux
    port map (
            O => \N__29760\,
            I => \Commands_frame_decoder.un1_WDT_cry_5\
        );

    \I__4393\ : InMux
    port map (
            O => \N__29757\,
            I => \Commands_frame_decoder.un1_WDT_cry_6\
        );

    \I__4392\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29751\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__29751\,
            I => \N__29748\
        );

    \I__4390\ : Odrv12
    port map (
            O => \N__29748\,
            I => drone_altitude_i_7
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__29745\,
            I => \N__29742\
        );

    \I__4388\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29739\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__29739\,
            I => \N__29735\
        );

    \I__4386\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29732\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__29735\,
            I => \N__29729\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__29732\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__29729\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__4382\ : InMux
    port map (
            O => \N__29724\,
            I => \N__29721\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__29721\,
            I => \N__29718\
        );

    \I__4380\ : Odrv12
    port map (
            O => \N__29718\,
            I => \pid_alt.error_axbZ0Z_13\
        );

    \I__4379\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29712\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__29712\,
            I => \N__29709\
        );

    \I__4377\ : Odrv12
    port map (
            O => \N__29709\,
            I => \pid_alt.error_axbZ0Z_14\
        );

    \I__4376\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29703\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__29703\,
            I => \N__29700\
        );

    \I__4374\ : Odrv12
    port map (
            O => \N__29700\,
            I => \pid_alt.error_axbZ0Z_12\
        );

    \I__4373\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29694\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__29694\,
            I => uart_input_drone_c
        );

    \I__4371\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29688\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__29688\,
            I => \uart_drone_sync.aux_0__0__0_0\
        );

    \I__4369\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29682\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__29682\,
            I => \uart_drone_sync.aux_1__0__0_0\
        );

    \I__4367\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29676\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__29676\,
            I => \uart_drone_sync.aux_2__0__0_0\
        );

    \I__4365\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29670\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__4363\ : Span4Mux_v
    port map (
            O => \N__29667\,
            I => \N__29664\
        );

    \I__4362\ : Span4Mux_h
    port map (
            O => \N__29664\,
            I => \N__29661\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__29661\,
            I => drone_altitude_15
        );

    \I__4360\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29655\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__29655\,
            I => \N__29652\
        );

    \I__4358\ : Span4Mux_v
    port map (
            O => \N__29652\,
            I => \N__29649\
        );

    \I__4357\ : Span4Mux_h
    port map (
            O => \N__29649\,
            I => \N__29646\
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__29646\,
            I => drone_altitude_i_4
        );

    \I__4355\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29640\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__29640\,
            I => \N__29637\
        );

    \I__4353\ : Span4Mux_v
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__4352\ : Span4Mux_h
    port map (
            O => \N__29634\,
            I => \N__29631\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__29631\,
            I => drone_altitude_i_5
        );

    \I__4350\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29625\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__29625\,
            I => \N__29622\
        );

    \I__4348\ : Span4Mux_s3_h
    port map (
            O => \N__29622\,
            I => \N__29619\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__29619\,
            I => \N__29616\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__29616\,
            I => drone_altitude_i_6
        );

    \I__4345\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29610\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__29610\,
            I => \dron_frame_decoder_1.drone_altitude_9\
        );

    \I__4343\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29604\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__29604\,
            I => \N__29601\
        );

    \I__4341\ : Span4Mux_s3_h
    port map (
            O => \N__29601\,
            I => \N__29598\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__29598\,
            I => \N__29595\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__29595\,
            I => drone_altitude_i_9
        );

    \I__4338\ : InMux
    port map (
            O => \N__29592\,
            I => \N__29589\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__29589\,
            I => \N__29586\
        );

    \I__4336\ : Span4Mux_s3_h
    port map (
            O => \N__29586\,
            I => \N__29583\
        );

    \I__4335\ : Span4Mux_h
    port map (
            O => \N__29583\,
            I => \N__29580\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__29580\,
            I => drone_altitude_i_8
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__29577\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_\
        );

    \I__4332\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29570\
        );

    \I__4331\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29567\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29564\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__29567\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__29564\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__4327\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29556\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__4325\ : Odrv4
    port map (
            O => \N__29553\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__4324\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29544\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__29549\,
            I => \N__29541\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__29548\,
            I => \N__29538\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \N__29535\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__29544\,
            I => \N__29532\
        );

    \I__4319\ : InMux
    port map (
            O => \N__29541\,
            I => \N__29529\
        );

    \I__4318\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29524\
        );

    \I__4317\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29524\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__29532\,
            I => \N__29521\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__29529\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__29524\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__29521\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4312\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29510\
        );

    \I__4311\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29507\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__29510\,
            I => \Commands_frame_decoder.stateZ0Z_4\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__29507\,
            I => \Commands_frame_decoder.stateZ0Z_4\
        );

    \I__4308\ : InMux
    port map (
            O => \N__29502\,
            I => \N__29499\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__29499\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__4306\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29493\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__4304\ : Odrv12
    port map (
            O => \N__29490\,
            I => \pid_front.O_0_6\
        );

    \I__4303\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__4301\ : Span4Mux_h
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__4300\ : Odrv4
    port map (
            O => \N__29478\,
            I => \pid_front.O_0_4\
        );

    \I__4299\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29472\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__29472\,
            I => \N__29469\
        );

    \I__4297\ : Span4Mux_v
    port map (
            O => \N__29469\,
            I => \N__29466\
        );

    \I__4296\ : Span4Mux_h
    port map (
            O => \N__29466\,
            I => \N__29463\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__29463\,
            I => \pid_front.O_0_9\
        );

    \I__4294\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__29454\,
            I => \N__29451\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__29451\,
            I => \N__29448\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__29448\,
            I => \pid_front.O_0_15\
        );

    \I__4289\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__4287\ : Odrv12
    port map (
            O => \N__29439\,
            I => \dron_frame_decoder_1.drone_altitude_11\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__29436\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\
        );

    \I__4285\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29427\
        );

    \I__4283\ : Span4Mux_v
    port map (
            O => \N__29427\,
            I => \N__29424\
        );

    \I__4282\ : Span4Mux_h
    port map (
            O => \N__29424\,
            I => \N__29420\
        );

    \I__4281\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29417\
        );

    \I__4280\ : Span4Mux_h
    port map (
            O => \N__29420\,
            I => \N__29414\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__29417\,
            I => \N__29411\
        );

    \I__4278\ : Span4Mux_h
    port map (
            O => \N__29414\,
            I => \N__29407\
        );

    \I__4277\ : Span4Mux_v
    port map (
            O => \N__29411\,
            I => \N__29404\
        );

    \I__4276\ : InMux
    port map (
            O => \N__29410\,
            I => \N__29401\
        );

    \I__4275\ : Span4Mux_h
    port map (
            O => \N__29407\,
            I => \N__29396\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__29404\,
            I => \N__29396\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__29401\,
            I => xy_kp_4
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__29396\,
            I => xy_kp_4
        );

    \I__4271\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29388\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__29388\,
            I => \N__29384\
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__29387\,
            I => \N__29380\
        );

    \I__4268\ : Span4Mux_v
    port map (
            O => \N__29384\,
            I => \N__29376\
        );

    \I__4267\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29369\
        );

    \I__4266\ : InMux
    port map (
            O => \N__29380\,
            I => \N__29369\
        );

    \I__4265\ : InMux
    port map (
            O => \N__29379\,
            I => \N__29369\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__29376\,
            I => \Commands_frame_decoder.stateZ0Z_7\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__29369\,
            I => \Commands_frame_decoder.stateZ0Z_7\
        );

    \I__4262\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29358\
        );

    \I__4261\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29358\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__29358\,
            I => \N__29355\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__29355\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__4258\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29348\
        );

    \I__4257\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29344\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__29348\,
            I => \N__29341\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__29347\,
            I => \N__29338\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__29344\,
            I => \N__29335\
        );

    \I__4253\ : Span4Mux_h
    port map (
            O => \N__29341\,
            I => \N__29332\
        );

    \I__4252\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29329\
        );

    \I__4251\ : Span12Mux_s11_v
    port map (
            O => \N__29335\,
            I => \N__29326\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__29332\,
            I => \N__29323\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__29329\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__4248\ : Odrv12
    port map (
            O => \N__29326\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__29323\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__4246\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29313\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__29313\,
            I => \N__29310\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__4243\ : Sp12to4
    port map (
            O => \N__29307\,
            I => \N__29303\
        );

    \I__4242\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29300\
        );

    \I__4241\ : Span12Mux_s7_h
    port map (
            O => \N__29303\,
            I => \N__29297\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__29300\,
            I => alt_kp_4
        );

    \I__4239\ : Odrv12
    port map (
            O => \N__29297\,
            I => alt_kp_4
        );

    \I__4238\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29289\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__29289\,
            I => \N__29283\
        );

    \I__4236\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29276\
        );

    \I__4235\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29276\
        );

    \I__4234\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29276\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__29283\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__29276\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__29271\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_\
        );

    \I__4230\ : InMux
    port map (
            O => \N__29268\,
            I => \N__29262\
        );

    \I__4229\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29262\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29259\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__29259\,
            I => \Commands_frame_decoder.N_378\
        );

    \I__4226\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29243\
        );

    \I__4225\ : InMux
    port map (
            O => \N__29255\,
            I => \N__29243\
        );

    \I__4224\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29243\
        );

    \I__4223\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29234\
        );

    \I__4222\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29234\
        );

    \I__4221\ : InMux
    port map (
            O => \N__29251\,
            I => \N__29234\
        );

    \I__4220\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29234\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__29243\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__29234\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__4217\ : CascadeMux
    port map (
            O => \N__29229\,
            I => \N__29224\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__29228\,
            I => \N__29219\
        );

    \I__4215\ : InMux
    port map (
            O => \N__29227\,
            I => \N__29211\
        );

    \I__4214\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29211\
        );

    \I__4213\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29211\
        );

    \I__4212\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29204\
        );

    \I__4211\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29204\
        );

    \I__4210\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29204\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__29211\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__29204\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__29199\,
            I => \N__29195\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__29198\,
            I => \N__29192\
        );

    \I__4205\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29189\
        );

    \I__4204\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29186\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__29189\,
            I => \N__29183\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__29186\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__4201\ : Odrv4
    port map (
            O => \N__29183\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__4200\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29175\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__29175\,
            I => \N__29172\
        );

    \I__4198\ : Span4Mux_h
    port map (
            O => \N__29172\,
            I => \N__29169\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__29169\,
            I => \Commands_frame_decoder.state_ns_0_i_1_1\
        );

    \I__4196\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__29163\,
            I => \N__29160\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__29160\,
            I => \N__29156\
        );

    \I__4193\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29153\
        );

    \I__4192\ : Span4Mux_v
    port map (
            O => \N__29156\,
            I => \N__29150\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29147\
        );

    \I__4190\ : Span4Mux_h
    port map (
            O => \N__29150\,
            I => \N__29144\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__29147\,
            I => \N__29141\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__29144\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__29141\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\
        );

    \I__4186\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29131\
        );

    \I__4185\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29126\
        );

    \I__4184\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29126\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__29131\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__29126\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__29121\,
            I => \uart_pc.N_126_li_cascade_\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__29118\,
            I => \N__29114\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__29117\,
            I => \N__29111\
        );

    \I__4178\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29101\
        );

    \I__4177\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29101\
        );

    \I__4176\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29101\
        );

    \I__4175\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29096\
        );

    \I__4174\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29096\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__29101\,
            I => \uart_pc.N_143\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__29096\,
            I => \uart_pc.N_143\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__29091\,
            I => \uart_pc.N_143_cascade_\
        );

    \I__4170\ : CascadeMux
    port map (
            O => \N__29088\,
            I => \N__29082\
        );

    \I__4169\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29079\
        );

    \I__4168\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29072\
        );

    \I__4167\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29072\
        );

    \I__4166\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29072\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__29079\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__29072\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__29067\,
            I => \N__29064\
        );

    \I__4162\ : InMux
    port map (
            O => \N__29064\,
            I => \N__29061\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__29061\,
            I => \N__29058\
        );

    \I__4160\ : Span4Mux_h
    port map (
            O => \N__29058\,
            I => \N__29055\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__29055\,
            I => \Commands_frame_decoder.state_ns_i_a2_0_2_0\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__29052\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\
        );

    \I__4157\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29046\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__29046\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_4\
        );

    \I__4155\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__29040\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_1\
        );

    \I__4153\ : InMux
    port map (
            O => \N__29037\,
            I => \N__29031\
        );

    \I__4152\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29031\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__29031\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__4150\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__29025\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_3\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__29022\,
            I => \uart_pc.N_144_1_cascade_\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__4146\ : InMux
    port map (
            O => \N__29016\,
            I => \N__29013\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__29013\,
            I => \uart_pc.un1_state_2_0_a3_0\
        );

    \I__4144\ : InMux
    port map (
            O => \N__29010\,
            I => \N__29007\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__29007\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_2\
        );

    \I__4142\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28998\
        );

    \I__4141\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28998\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__28998\,
            I => \N__28995\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__28995\,
            I => \pid_alt.N_44\
        );

    \I__4138\ : InMux
    port map (
            O => \N__28992\,
            I => \N__28988\
        );

    \I__4137\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28985\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28982\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28979\
        );

    \I__4134\ : Span4Mux_v
    port map (
            O => \N__28982\,
            I => \N__28976\
        );

    \I__4133\ : Span4Mux_h
    port map (
            O => \N__28979\,
            I => \N__28973\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__28976\,
            I => \pid_alt.pid_preregZ0Z_5\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__28973\,
            I => \pid_alt.pid_preregZ0Z_5\
        );

    \I__4130\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28962\
        );

    \I__4129\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28962\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N__28956\
        );

    \I__4127\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28953\
        );

    \I__4126\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28950\
        );

    \I__4125\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28947\
        );

    \I__4124\ : Span4Mux_v
    port map (
            O => \N__28956\,
            I => \N__28942\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__28953\,
            I => \N__28942\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__28950\,
            I => \N__28938\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__28947\,
            I => \N__28935\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__28942\,
            I => \N__28932\
        );

    \I__4119\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28929\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__28938\,
            I => \N__28926\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__28935\,
            I => \N__28923\
        );

    \I__4116\ : Span4Mux_h
    port map (
            O => \N__28932\,
            I => \N__28918\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__28929\,
            I => \N__28918\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__28926\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__28923\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__28918\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__28911\,
            I => \N__28907\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__28910\,
            I => \N__28896\
        );

    \I__4109\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28891\
        );

    \I__4108\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28891\
        );

    \I__4107\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28888\
        );

    \I__4106\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28881\
        );

    \I__4105\ : InMux
    port map (
            O => \N__28903\,
            I => \N__28881\
        );

    \I__4104\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28881\
        );

    \I__4103\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28876\
        );

    \I__4102\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28876\
        );

    \I__4101\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28873\
        );

    \I__4100\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28870\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N__28867\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__28888\,
            I => \N__28862\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__28881\,
            I => \N__28862\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__28876\,
            I => \N__28855\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28855\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28855\
        );

    \I__4093\ : Span4Mux_h
    port map (
            O => \N__28867\,
            I => \N__28848\
        );

    \I__4092\ : Span4Mux_v
    port map (
            O => \N__28862\,
            I => \N__28848\
        );

    \I__4091\ : Span4Mux_v
    port map (
            O => \N__28855\,
            I => \N__28848\
        );

    \I__4090\ : Sp12to4
    port map (
            O => \N__28848\,
            I => \N__28845\
        );

    \I__4089\ : Span12Mux_s3_h
    port map (
            O => \N__28845\,
            I => \N__28842\
        );

    \I__4088\ : Odrv12
    port map (
            O => \N__28842\,
            I => \pid_alt.pid_preregZ0Z_24\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__28839\,
            I => \N__28829\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__28838\,
            I => \N__28826\
        );

    \I__4085\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28815\
        );

    \I__4084\ : InMux
    port map (
            O => \N__28836\,
            I => \N__28815\
        );

    \I__4083\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28815\
        );

    \I__4082\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28815\
        );

    \I__4081\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28812\
        );

    \I__4080\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28809\
        );

    \I__4079\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28799\
        );

    \I__4078\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28799\
        );

    \I__4077\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28799\
        );

    \I__4076\ : InMux
    port map (
            O => \N__28824\,
            I => \N__28799\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__28815\,
            I => \N__28794\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__28812\,
            I => \N__28794\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28791\
        );

    \I__4072\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28788\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__28799\,
            I => \pid_alt.N_305\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__28794\,
            I => \pid_alt.N_305\
        );

    \I__4069\ : Odrv12
    port map (
            O => \N__28791\,
            I => \pid_alt.N_305\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__28788\,
            I => \pid_alt.N_305\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__28779\,
            I => \N__28775\
        );

    \I__4066\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28771\
        );

    \I__4065\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28768\
        );

    \I__4064\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28765\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__28771\,
            I => \N__28761\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28758\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__28765\,
            I => \N__28755\
        );

    \I__4060\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28752\
        );

    \I__4059\ : Span4Mux_v
    port map (
            O => \N__28761\,
            I => \N__28749\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__28758\,
            I => \N__28746\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__28755\,
            I => \N__28743\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28740\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__28749\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__28746\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__28743\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__4052\ : Odrv12
    port map (
            O => \N__28740\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__4051\ : CEMux
    port map (
            O => \N__28731\,
            I => \N__28727\
        );

    \I__4050\ : CEMux
    port map (
            O => \N__28730\,
            I => \N__28724\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28719\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__28724\,
            I => \N__28719\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__28719\,
            I => \pid_alt.N_72_i_1\
        );

    \I__4046\ : SRMux
    port map (
            O => \N__28716\,
            I => \N__28712\
        );

    \I__4045\ : SRMux
    port map (
            O => \N__28715\,
            I => \N__28709\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__28712\,
            I => \N__28703\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__28709\,
            I => \N__28703\
        );

    \I__4042\ : SRMux
    port map (
            O => \N__28708\,
            I => \N__28700\
        );

    \I__4041\ : Sp12to4
    port map (
            O => \N__28703\,
            I => \N__28694\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__28700\,
            I => \N__28694\
        );

    \I__4039\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28691\
        );

    \I__4038\ : Odrv12
    port map (
            O => \N__28694\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__28691\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4036\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28682\
        );

    \I__4035\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28679\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28674\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__28679\,
            I => \N__28674\
        );

    \I__4032\ : Span4Mux_v
    port map (
            O => \N__28674\,
            I => \N__28671\
        );

    \I__4031\ : Span4Mux_v
    port map (
            O => \N__28671\,
            I => \N__28668\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__28668\,
            I => \pid_alt.error_d_reg_prevZ0Z_17\
        );

    \I__4029\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28662\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__28662\,
            I => \N__28658\
        );

    \I__4027\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28655\
        );

    \I__4026\ : Span4Mux_v
    port map (
            O => \N__28658\,
            I => \N__28650\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__28655\,
            I => \N__28650\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__28650\,
            I => \N__28647\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__28647\,
            I => \pid_alt.error_p_regZ0Z_17\
        );

    \I__4022\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28641\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__28641\,
            I => \N__28637\
        );

    \I__4020\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28634\
        );

    \I__4019\ : Span4Mux_v
    port map (
            O => \N__28637\,
            I => \N__28628\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__28634\,
            I => \N__28628\
        );

    \I__4017\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28625\
        );

    \I__4016\ : Span4Mux_h
    port map (
            O => \N__28628\,
            I => \N__28622\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__28625\,
            I => \N__28619\
        );

    \I__4014\ : Span4Mux_v
    port map (
            O => \N__28622\,
            I => \N__28616\
        );

    \I__4013\ : Span4Mux_h
    port map (
            O => \N__28619\,
            I => \N__28611\
        );

    \I__4012\ : Span4Mux_v
    port map (
            O => \N__28616\,
            I => \N__28611\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__4010\ : Odrv4
    port map (
            O => \N__28608\,
            I => \pid_alt.error_d_regZ0Z_17\
        );

    \I__4009\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28601\
        );

    \I__4008\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28598\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28595\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__28598\,
            I => \N__28592\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__28595\,
            I => \N__28589\
        );

    \I__4004\ : Span4Mux_h
    port map (
            O => \N__28592\,
            I => \N__28586\
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__28589\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__28586\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\
        );

    \I__4001\ : InMux
    port map (
            O => \N__28581\,
            I => \uart_pc.un4_timer_Count_1_cry_1\
        );

    \I__4000\ : InMux
    port map (
            O => \N__28578\,
            I => \uart_pc.un4_timer_Count_1_cry_2\
        );

    \I__3999\ : InMux
    port map (
            O => \N__28575\,
            I => \uart_pc.un4_timer_Count_1_cry_3\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__28572\,
            I => \pid_alt.N_90_cascade_\
        );

    \I__3997\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28563\
        );

    \I__3996\ : InMux
    port map (
            O => \N__28568\,
            I => \N__28563\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__28563\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0_2\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__28560\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_\
        );

    \I__3993\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28553\
        );

    \I__3992\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28550\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__28553\,
            I => \pid_alt.N_43\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__28550\,
            I => \pid_alt.N_43\
        );

    \I__3989\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28542\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__28542\,
            I => \N__28539\
        );

    \I__3987\ : Odrv12
    port map (
            O => \N__28539\,
            I => \pid_alt.N_48\
        );

    \I__3986\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__28533\,
            I => \N__28530\
        );

    \I__3984\ : Odrv12
    port map (
            O => \N__28530\,
            I => \pid_alt.pid_preregZ0Z_15\
        );

    \I__3983\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__28521\,
            I => \N__28518\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__28518\,
            I => \pid_alt.pid_preregZ0Z_23\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__28515\,
            I => \N__28512\
        );

    \I__3978\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28509\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__28509\,
            I => \N__28506\
        );

    \I__3976\ : Span4Mux_h
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__28503\,
            I => \pid_alt.pid_preregZ0Z_21\
        );

    \I__3974\ : InMux
    port map (
            O => \N__28500\,
            I => \N__28497\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__28497\,
            I => \N__28494\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__28494\,
            I => \pid_alt.pid_preregZ0Z_18\
        );

    \I__3971\ : InMux
    port map (
            O => \N__28491\,
            I => \N__28488\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__28488\,
            I => \N__28485\
        );

    \I__3969\ : Span4Mux_h
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__28482\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3967\ : InMux
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__28476\,
            I => \N__28473\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__28473\,
            I => \pid_alt.pid_preregZ0Z_20\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__28470\,
            I => \N__28467\
        );

    \I__3963\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28464\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__28464\,
            I => \N__28461\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__28461\,
            I => \pid_alt.pid_preregZ0Z_17\
        );

    \I__3960\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__28452\,
            I => \pid_alt.pid_preregZ0Z_19\
        );

    \I__3957\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__28446\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_2_6\
        );

    \I__3955\ : InMux
    port map (
            O => \N__28443\,
            I => \N__28440\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__28440\,
            I => \N__28437\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__3952\ : Odrv4
    port map (
            O => \N__28434\,
            I => \pid_alt.pid_preregZ0Z_14\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__28431\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_\
        );

    \I__3950\ : InMux
    port map (
            O => \N__28428\,
            I => \N__28425\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__28422\,
            I => \pid_alt.pid_preregZ0Z_16\
        );

    \I__3947\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28416\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__28416\,
            I => \N__28411\
        );

    \I__3945\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28408\
        );

    \I__3944\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28405\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__28411\,
            I => \pid_alt.N_90\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__28408\,
            I => \pid_alt.N_90\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__28405\,
            I => \pid_alt.N_90\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__28398\,
            I => \pid_alt.N_305_cascade_\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__28395\,
            I => \pid_alt.source_pid_9_0_0_4_cascade_\
        );

    \I__3938\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28383\
        );

    \I__3937\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28383\
        );

    \I__3936\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28378\
        );

    \I__3935\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28378\
        );

    \I__3934\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28375\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__28383\,
            I => \N__28372\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__28378\,
            I => \N__28369\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__28375\,
            I => \N__28366\
        );

    \I__3930\ : Span4Mux_v
    port map (
            O => \N__28372\,
            I => \N__28361\
        );

    \I__3929\ : Span4Mux_v
    port map (
            O => \N__28369\,
            I => \N__28361\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__28366\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__28361\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__3926\ : CascadeMux
    port map (
            O => \N__28356\,
            I => \pid_alt.N_44_cascade_\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__3924\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28341\
        );

    \I__3923\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28341\
        );

    \I__3922\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28341\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__28341\,
            I => \pid_alt.N_46\
        );

    \I__3920\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28332\
        );

    \I__3919\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28332\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__28332\,
            I => \N__28329\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__28329\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__28326\,
            I => \pid_alt.N_46_cascade_\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__28323\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_\
        );

    \I__3914\ : InMux
    port map (
            O => \N__28320\,
            I => \N__28317\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__28317\,
            I => \N__28314\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__28314\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_1_7\
        );

    \I__3911\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__28308\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_1_4\
        );

    \I__3909\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28302\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__28302\,
            I => \N__28297\
        );

    \I__3907\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28292\
        );

    \I__3906\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28292\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__28297\,
            I => \N__28289\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__28292\,
            I => \N__28286\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__28289\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__28286\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__3901\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28277\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__28280\,
            I => \N__28274\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__28277\,
            I => \N__28270\
        );

    \I__3898\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28265\
        );

    \I__3897\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28265\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__28270\,
            I => \N__28260\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__28265\,
            I => \N__28260\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__28260\,
            I => \pid_alt.pid_preregZ0Z_9\
        );

    \I__3893\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28253\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__28256\,
            I => \N__28249\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__28253\,
            I => \N__28246\
        );

    \I__3890\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28243\
        );

    \I__3889\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28240\
        );

    \I__3888\ : Span4Mux_v
    port map (
            O => \N__28246\,
            I => \N__28233\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__28243\,
            I => \N__28233\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28233\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__28233\,
            I => \pid_alt.pid_preregZ0Z_10\
        );

    \I__3884\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28227\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__28227\,
            I => \N__28222\
        );

    \I__3882\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28217\
        );

    \I__3881\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28217\
        );

    \I__3880\ : Span4Mux_h
    port map (
            O => \N__28222\,
            I => \N__28214\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__28217\,
            I => \N__28211\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__28214\,
            I => \pid_alt.pid_preregZ0Z_8\
        );

    \I__3877\ : Odrv12
    port map (
            O => \N__28211\,
            I => \pid_alt.pid_preregZ0Z_8\
        );

    \I__3876\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28202\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__28205\,
            I => \N__28199\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__28202\,
            I => \N__28195\
        );

    \I__3873\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28190\
        );

    \I__3872\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28190\
        );

    \I__3871\ : Span4Mux_v
    port map (
            O => \N__28195\,
            I => \N__28185\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28185\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__28185\,
            I => \pid_alt.pid_preregZ0Z_7\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__28182\,
            I => \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_\
        );

    \I__3867\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28174\
        );

    \I__3866\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28169\
        );

    \I__3865\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28169\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__28174\,
            I => \N__28166\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__28169\,
            I => \N__28163\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__28166\,
            I => \N__28160\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__28163\,
            I => \N__28157\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__28160\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__28157\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__3858\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28137\
        );

    \I__3857\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28137\
        );

    \I__3856\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28137\
        );

    \I__3855\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28137\
        );

    \I__3854\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28137\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__28137\,
            I => \pid_alt.source_pid_9_0_tz_6\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__3851\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28125\
        );

    \I__3850\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28125\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__28122\,
            I => \pid_alt.pid_preregZ0Z_2\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__28119\,
            I => \N__28115\
        );

    \I__3846\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28110\
        );

    \I__3845\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28110\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__28110\,
            I => \N__28107\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__28107\,
            I => \pid_alt.pid_preregZ0Z_3\
        );

    \I__3842\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28098\
        );

    \I__3841\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28098\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__28098\,
            I => \N__28095\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__28095\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__3838\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28089\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__28089\,
            I => \N__28086\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__28086\,
            I => \pid_alt.m21_e_9\
        );

    \I__3835\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__28080\,
            I => \pid_alt.m21_e_10\
        );

    \I__3833\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28073\
        );

    \I__3832\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28070\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__28073\,
            I => \pid_alt.N_9_0\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__28070\,
            I => \pid_alt.N_9_0\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__28065\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNIO7B05Z0Z_21_cascade_\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__28062\,
            I => \pid_alt.un1_reset_1_0_i_cascade_\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__28059\,
            I => \N__28055\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__28058\,
            I => \N__28051\
        );

    \I__3825\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28048\
        );

    \I__3824\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28043\
        );

    \I__3823\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28043\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__28048\,
            I => \N__28040\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28034\
        );

    \I__3820\ : Span4Mux_h
    port map (
            O => \N__28040\,
            I => \N__28034\
        );

    \I__3819\ : InMux
    port map (
            O => \N__28039\,
            I => \N__28031\
        );

    \I__3818\ : Span4Mux_v
    port map (
            O => \N__28034\,
            I => \N__28028\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__28031\,
            I => \N__28025\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__28028\,
            I => \N__28022\
        );

    \I__3815\ : Span12Mux_v
    port map (
            O => \N__28025\,
            I => \N__28019\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__28022\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__3813\ : Odrv12
    port map (
            O => \N__28019\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__3812\ : InMux
    port map (
            O => \N__28014\,
            I => \N__28010\
        );

    \I__3811\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28007\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__28010\,
            I => \N__28001\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__28007\,
            I => \N__28001\
        );

    \I__3808\ : InMux
    port map (
            O => \N__28006\,
            I => \N__27998\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__28001\,
            I => \N__27995\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__27998\,
            I => \N__27992\
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__27995\,
            I => \pid_alt.error_i_acumm7lto13\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__27992\,
            I => \pid_alt.error_i_acumm7lto13\
        );

    \I__3803\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27984\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27980\
        );

    \I__3801\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27976\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__27980\,
            I => \N__27973\
        );

    \I__3799\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27970\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__27976\,
            I => \N__27967\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__27973\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__27970\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__27967\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14\
        );

    \I__3794\ : InMux
    port map (
            O => \N__27960\,
            I => \N__27957\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__27957\,
            I => \N__27954\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__27954\,
            I => \pid_alt.error_i_acummZ0Z_13\
        );

    \I__3791\ : CEMux
    port map (
            O => \N__27951\,
            I => \N__27947\
        );

    \I__3790\ : CEMux
    port map (
            O => \N__27950\,
            I => \N__27944\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__27947\,
            I => \pid_alt.N_72_i_0\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__27944\,
            I => \pid_alt.N_72_i_0\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__27939\,
            I => \pid_alt.un1_reset_1_cascade_\
        );

    \I__3786\ : CascadeMux
    port map (
            O => \N__27936\,
            I => \pid_alt.source_pid_9_0_tz_6_cascade_\
        );

    \I__3785\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27929\
        );

    \I__3784\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27926\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27922\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27919\
        );

    \I__3781\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27916\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__27922\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__27919\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__27916\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__3777\ : CascadeMux
    port map (
            O => \N__27909\,
            I => \pid_alt.m21_e_0_cascade_\
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__27906\,
            I => \N__27901\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__27905\,
            I => \N__27897\
        );

    \I__3774\ : InMux
    port map (
            O => \N__27904\,
            I => \N__27888\
        );

    \I__3773\ : InMux
    port map (
            O => \N__27901\,
            I => \N__27888\
        );

    \I__3772\ : InMux
    port map (
            O => \N__27900\,
            I => \N__27888\
        );

    \I__3771\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27883\
        );

    \I__3770\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27883\
        );

    \I__3769\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27880\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__27888\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__27883\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__27880\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__3765\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27870\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__27870\,
            I => \pid_alt.m35_e_3\
        );

    \I__3763\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27862\
        );

    \I__3762\ : InMux
    port map (
            O => \N__27866\,
            I => \N__27857\
        );

    \I__3761\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27857\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__27862\,
            I => \N__27854\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__27857\,
            I => \N__27851\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__27854\,
            I => \N__27848\
        );

    \I__3757\ : Span4Mux_v
    port map (
            O => \N__27851\,
            I => \N__27845\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__27848\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__27845\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\
        );

    \I__3754\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27837\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__27837\,
            I => \N__27832\
        );

    \I__3752\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27827\
        );

    \I__3751\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27827\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__27832\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__27827\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\
        );

    \I__3748\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__3746\ : Span4Mux_v
    port map (
            O => \N__27816\,
            I => \N__27811\
        );

    \I__3745\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27806\
        );

    \I__3744\ : InMux
    port map (
            O => \N__27814\,
            I => \N__27806\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__27811\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__27806\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__27801\,
            I => \N__27798\
        );

    \I__3740\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27793\
        );

    \I__3739\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27788\
        );

    \I__3738\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27788\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__27793\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__27788\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__3735\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27778\
        );

    \I__3734\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27773\
        );

    \I__3733\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27773\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__27778\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__27773\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__27768\,
            I => \N__27763\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__27767\,
            I => \N__27760\
        );

    \I__3728\ : InMux
    port map (
            O => \N__27766\,
            I => \N__27757\
        );

    \I__3727\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27752\
        );

    \I__3726\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27752\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__27757\,
            I => \N__27749\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__27752\,
            I => \N__27746\
        );

    \I__3723\ : Span4Mux_h
    port map (
            O => \N__27749\,
            I => \N__27743\
        );

    \I__3722\ : Span4Mux_h
    port map (
            O => \N__27746\,
            I => \N__27740\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__27743\,
            I => \pid_alt.error_i_acumm_preregZ0Z_11\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__27740\,
            I => \pid_alt.error_i_acumm_preregZ0Z_11\
        );

    \I__3719\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27728\
        );

    \I__3718\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27728\
        );

    \I__3717\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27725\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__27728\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__27725\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__3714\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27716\
        );

    \I__3713\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27713\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__27716\,
            I => \N__27708\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__27713\,
            I => \N__27708\
        );

    \I__3710\ : Span4Mux_h
    port map (
            O => \N__27708\,
            I => \N__27705\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__27705\,
            I => \pid_alt.error_i_acumm_preregZ0Z_1\
        );

    \I__3708\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27698\
        );

    \I__3707\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27695\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__27698\,
            I => \N__27692\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__27695\,
            I => \N__27689\
        );

    \I__3704\ : Odrv12
    port map (
            O => \N__27692\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__3703\ : Odrv4
    port map (
            O => \N__27689\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__27684\,
            I => \pid_alt.m21_e_8_cascade_\
        );

    \I__3701\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__27678\,
            I => \N__27673\
        );

    \I__3699\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27670\
        );

    \I__3698\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27667\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__27673\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__27670\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__27667\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__3694\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27657\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__27657\,
            I => \pid_alt.m21_e_2\
        );

    \I__3692\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27651\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__27651\,
            I => \N__27648\
        );

    \I__3690\ : Span4Mux_h
    port map (
            O => \N__27648\,
            I => \N__27643\
        );

    \I__3689\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27640\
        );

    \I__3688\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27637\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__27643\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__27640\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__27637\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__3684\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27625\
        );

    \I__3683\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27620\
        );

    \I__3682\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27620\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__27625\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__27620\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__3679\ : CEMux
    port map (
            O => \N__27615\,
            I => \N__27546\
        );

    \I__3678\ : CEMux
    port map (
            O => \N__27614\,
            I => \N__27546\
        );

    \I__3677\ : CEMux
    port map (
            O => \N__27613\,
            I => \N__27546\
        );

    \I__3676\ : CEMux
    port map (
            O => \N__27612\,
            I => \N__27546\
        );

    \I__3675\ : CEMux
    port map (
            O => \N__27611\,
            I => \N__27546\
        );

    \I__3674\ : CEMux
    port map (
            O => \N__27610\,
            I => \N__27546\
        );

    \I__3673\ : CEMux
    port map (
            O => \N__27609\,
            I => \N__27546\
        );

    \I__3672\ : CEMux
    port map (
            O => \N__27608\,
            I => \N__27546\
        );

    \I__3671\ : CEMux
    port map (
            O => \N__27607\,
            I => \N__27546\
        );

    \I__3670\ : CEMux
    port map (
            O => \N__27606\,
            I => \N__27546\
        );

    \I__3669\ : CEMux
    port map (
            O => \N__27605\,
            I => \N__27546\
        );

    \I__3668\ : CEMux
    port map (
            O => \N__27604\,
            I => \N__27546\
        );

    \I__3667\ : CEMux
    port map (
            O => \N__27603\,
            I => \N__27546\
        );

    \I__3666\ : CEMux
    port map (
            O => \N__27602\,
            I => \N__27546\
        );

    \I__3665\ : CEMux
    port map (
            O => \N__27601\,
            I => \N__27546\
        );

    \I__3664\ : CEMux
    port map (
            O => \N__27600\,
            I => \N__27546\
        );

    \I__3663\ : CEMux
    port map (
            O => \N__27599\,
            I => \N__27546\
        );

    \I__3662\ : CEMux
    port map (
            O => \N__27598\,
            I => \N__27546\
        );

    \I__3661\ : CEMux
    port map (
            O => \N__27597\,
            I => \N__27546\
        );

    \I__3660\ : CEMux
    port map (
            O => \N__27596\,
            I => \N__27546\
        );

    \I__3659\ : CEMux
    port map (
            O => \N__27595\,
            I => \N__27546\
        );

    \I__3658\ : CEMux
    port map (
            O => \N__27594\,
            I => \N__27546\
        );

    \I__3657\ : CEMux
    port map (
            O => \N__27593\,
            I => \N__27546\
        );

    \I__3656\ : GlobalMux
    port map (
            O => \N__27546\,
            I => \N__27543\
        );

    \I__3655\ : gio2CtrlBuf
    port map (
            O => \N__27543\,
            I => \pid_alt.state_0_g_0\
        );

    \I__3654\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27536\
        );

    \I__3653\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27533\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__27536\,
            I => \Commands_frame_decoder.N_416\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__27533\,
            I => \Commands_frame_decoder.N_416\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__27528\,
            I => \Commands_frame_decoder.N_379_cascade_\
        );

    \I__3649\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27517\
        );

    \I__3648\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27517\
        );

    \I__3647\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27512\
        );

    \I__3646\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27512\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__27517\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__27512\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__3643\ : InMux
    port map (
            O => \N__27507\,
            I => \N__27504\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__27504\,
            I => \Commands_frame_decoder.N_412\
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__27501\,
            I => \N__27498\
        );

    \I__3640\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27492\
        );

    \I__3639\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27492\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__27492\,
            I => \Commands_frame_decoder.stateZ0Z_8\
        );

    \I__3637\ : CEMux
    port map (
            O => \N__27489\,
            I => \N__27485\
        );

    \I__3636\ : CEMux
    port map (
            O => \N__27488\,
            I => \N__27480\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__27485\,
            I => \N__27477\
        );

    \I__3634\ : CEMux
    port map (
            O => \N__27484\,
            I => \N__27474\
        );

    \I__3633\ : CEMux
    port map (
            O => \N__27483\,
            I => \N__27471\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__27480\,
            I => \N__27468\
        );

    \I__3631\ : Span4Mux_v
    port map (
            O => \N__27477\,
            I => \N__27463\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__27474\,
            I => \N__27463\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__27471\,
            I => \N__27460\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__27468\,
            I => \N__27457\
        );

    \I__3627\ : Span4Mux_v
    port map (
            O => \N__27463\,
            I => \N__27454\
        );

    \I__3626\ : Span4Mux_h
    port map (
            O => \N__27460\,
            I => \N__27451\
        );

    \I__3625\ : Span4Mux_v
    port map (
            O => \N__27457\,
            I => \N__27448\
        );

    \I__3624\ : Span4Mux_v
    port map (
            O => \N__27454\,
            I => \N__27445\
        );

    \I__3623\ : Span4Mux_v
    port map (
            O => \N__27451\,
            I => \N__27442\
        );

    \I__3622\ : Span4Mux_v
    port map (
            O => \N__27448\,
            I => \N__27439\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__27445\,
            I => \N__27436\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__27442\,
            I => \N__27433\
        );

    \I__3619\ : Odrv4
    port map (
            O => \N__27439\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__27436\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__27433\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__3616\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27422\
        );

    \I__3615\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27419\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__27422\,
            I => \Commands_frame_decoder.stateZ0Z_9\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__27419\,
            I => \Commands_frame_decoder.stateZ0Z_9\
        );

    \I__3612\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27396\
        );

    \I__3611\ : InMux
    port map (
            O => \N__27413\,
            I => \N__27396\
        );

    \I__3610\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27396\
        );

    \I__3609\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27396\
        );

    \I__3608\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27396\
        );

    \I__3607\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27396\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__27396\,
            I => \N__27390\
        );

    \I__3605\ : InMux
    port map (
            O => \N__27395\,
            I => \N__27383\
        );

    \I__3604\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27383\
        );

    \I__3603\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27383\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__27390\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__27383\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12\
        );

    \I__3600\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27374\
        );

    \I__3599\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27371\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__27374\,
            I => \pid_alt.error_i_acumm_preregZ0Z_3\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__27371\,
            I => \pid_alt.error_i_acumm_preregZ0Z_3\
        );

    \I__3596\ : InMux
    port map (
            O => \N__27366\,
            I => \N__27363\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__27363\,
            I => \N__27359\
        );

    \I__3594\ : InMux
    port map (
            O => \N__27362\,
            I => \N__27356\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__27359\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__27356\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__27351\,
            I => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__27348\,
            I => \Commands_frame_decoder.N_416_cascade_\
        );

    \I__3589\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__27342\,
            I => \Commands_frame_decoder.N_382\
        );

    \I__3587\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27336\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__27336\,
            I => \Commands_frame_decoder.state_ns_0_a3_0_2_2\
        );

    \I__3585\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27329\
        );

    \I__3584\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27326\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__27329\,
            I => \Commands_frame_decoder.N_376_2\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__27326\,
            I => \Commands_frame_decoder.N_376_2\
        );

    \I__3581\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27318\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__27318\,
            I => \Commands_frame_decoder.N_377\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__27315\,
            I => \Commands_frame_decoder.N_376_cascade_\
        );

    \I__3578\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27309\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__27309\,
            I => \Commands_frame_decoder.N_379\
        );

    \I__3576\ : InMux
    port map (
            O => \N__27306\,
            I => \N__27302\
        );

    \I__3575\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27299\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__27302\,
            I => \N__27296\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__27299\,
            I => \N__27293\
        );

    \I__3572\ : Span4Mux_v
    port map (
            O => \N__27296\,
            I => \N__27290\
        );

    \I__3571\ : Span4Mux_v
    port map (
            O => \N__27293\,
            I => \N__27287\
        );

    \I__3570\ : Odrv4
    port map (
            O => \N__27290\,
            I => \pid_alt.error_p_regZ0Z_19\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__27287\,
            I => \pid_alt.error_p_regZ0Z_19\
        );

    \I__3568\ : InMux
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__27279\,
            I => \N__27276\
        );

    \I__3566\ : Span4Mux_h
    port map (
            O => \N__27276\,
            I => \N__27272\
        );

    \I__3565\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27269\
        );

    \I__3564\ : Sp12to4
    port map (
            O => \N__27272\,
            I => \N__27266\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__27269\,
            I => \pid_alt.error_d_reg_prevZ0Z_19\
        );

    \I__3562\ : Odrv12
    port map (
            O => \N__27266\,
            I => \pid_alt.error_d_reg_prevZ0Z_19\
        );

    \I__3561\ : InMux
    port map (
            O => \N__27261\,
            I => \N__27255\
        );

    \I__3560\ : InMux
    port map (
            O => \N__27260\,
            I => \N__27255\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__3558\ : Span4Mux_v
    port map (
            O => \N__27252\,
            I => \N__27248\
        );

    \I__3557\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27245\
        );

    \I__3556\ : Sp12to4
    port map (
            O => \N__27248\,
            I => \N__27240\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__27245\,
            I => \N__27240\
        );

    \I__3554\ : Span12Mux_s7_h
    port map (
            O => \N__27240\,
            I => \N__27237\
        );

    \I__3553\ : Span12Mux_v
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__3552\ : Odrv12
    port map (
            O => \N__27234\,
            I => \pid_alt.error_d_regZ0Z_19\
        );

    \I__3551\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27228\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__27228\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\
        );

    \I__3549\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27222\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__27222\,
            I => \N__27218\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__27221\,
            I => \N__27215\
        );

    \I__3546\ : Span12Mux_h
    port map (
            O => \N__27218\,
            I => \N__27212\
        );

    \I__3545\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27209\
        );

    \I__3544\ : Odrv12
    port map (
            O => \N__27212\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__27209\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__27204\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_\
        );

    \I__3541\ : InMux
    port map (
            O => \N__27201\,
            I => \N__27194\
        );

    \I__3540\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27194\
        );

    \I__3539\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27191\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__27194\,
            I => \N__27188\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__27191\,
            I => \N__27185\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__27188\,
            I => \N__27182\
        );

    \I__3535\ : Odrv12
    port map (
            O => \N__27185\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__27182\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\
        );

    \I__3533\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__27174\,
            I => \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\
        );

    \I__3531\ : InMux
    port map (
            O => \N__27171\,
            I => \N__27165\
        );

    \I__3530\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27165\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__27165\,
            I => \N__27162\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__27162\,
            I => \N__27159\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__27159\,
            I => \pid_alt.error_p_regZ0Z_20\
        );

    \I__3526\ : InMux
    port map (
            O => \N__27156\,
            I => \N__27150\
        );

    \I__3525\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27150\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__27150\,
            I => \pid_alt.error_d_reg_prevZ0Z_20\
        );

    \I__3523\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27138\
        );

    \I__3522\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27138\
        );

    \I__3521\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27138\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__27138\,
            I => \N__27135\
        );

    \I__3519\ : Span4Mux_h
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__3518\ : Sp12to4
    port map (
            O => \N__27132\,
            I => \N__27129\
        );

    \I__3517\ : Span12Mux_v
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__3516\ : Odrv12
    port map (
            O => \N__27126\,
            I => \pid_alt.error_d_regZ0Z_20\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__3514\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27114\
        );

    \I__3513\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27107\
        );

    \I__3512\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27107\
        );

    \I__3511\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27107\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__27114\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__27107\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__27102\,
            I => \N__27098\
        );

    \I__3507\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27095\
        );

    \I__3506\ : InMux
    port map (
            O => \N__27098\,
            I => \N__27092\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__27095\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__27092\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__27087\,
            I => \N__27083\
        );

    \I__3502\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27076\
        );

    \I__3501\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27069\
        );

    \I__3500\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27069\
        );

    \I__3499\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27069\
        );

    \I__3498\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27064\
        );

    \I__3497\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27064\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__27076\,
            I => \pid_alt.un1_pid_prereg_236_1\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__27069\,
            I => \pid_alt.un1_pid_prereg_236_1\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__27064\,
            I => \pid_alt.un1_pid_prereg_236_1\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__27057\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20_cascade_\
        );

    \I__3492\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27046\
        );

    \I__3491\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27043\
        );

    \I__3490\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27034\
        );

    \I__3489\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27034\
        );

    \I__3488\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27034\
        );

    \I__3487\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27034\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__27046\,
            I => \N__27031\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__27043\,
            I => \N__27026\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__27034\,
            I => \N__27026\
        );

    \I__3483\ : Span4Mux_v
    port map (
            O => \N__27031\,
            I => \N__27023\
        );

    \I__3482\ : Odrv12
    port map (
            O => \N__27026\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__27023\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__3480\ : InMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__27015\,
            I => \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__27012\,
            I => \N__27008\
        );

    \I__3477\ : InMux
    port map (
            O => \N__27011\,
            I => \N__27005\
        );

    \I__3476\ : InMux
    port map (
            O => \N__27008\,
            I => \N__27001\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__27005\,
            I => \N__26998\
        );

    \I__3474\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26995\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__27001\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__26998\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__26995\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__26988\,
            I => \N__26984\
        );

    \I__3469\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26979\
        );

    \I__3468\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26979\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__26979\,
            I => \Commands_frame_decoder.stateZ0Z_12\
        );

    \I__3466\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26970\
        );

    \I__3465\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26970\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__26970\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__26967\,
            I => \N__26964\
        );

    \I__3462\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26960\
        );

    \I__3461\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26957\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__26960\,
            I => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__26957\,
            I => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\
        );

    \I__3458\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26943\
        );

    \I__3457\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26943\
        );

    \I__3456\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26943\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__26943\,
            I => \N__26940\
        );

    \I__3454\ : Span4Mux_v
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__26934\,
            I => \N__26931\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__26931\,
            I => \N__26928\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__26928\,
            I => \pid_alt.error_d_regZ0Z_16\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__26925\,
            I => \N__26922\
        );

    \I__3448\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26916\
        );

    \I__3447\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26916\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__26916\,
            I => \pid_alt.error_d_reg_prevZ0Z_16\
        );

    \I__3445\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26907\
        );

    \I__3444\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26907\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__26904\,
            I => \N__26901\
        );

    \I__3441\ : Span4Mux_s1_h
    port map (
            O => \N__26901\,
            I => \N__26898\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__26898\,
            I => \pid_alt.error_p_regZ0Z_16\
        );

    \I__3439\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__26892\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__26889\,
            I => \N__26885\
        );

    \I__3436\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26882\
        );

    \I__3435\ : InMux
    port map (
            O => \N__26885\,
            I => \N__26879\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__26882\,
            I => \N__26874\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__26879\,
            I => \N__26874\
        );

    \I__3432\ : Span4Mux_v
    port map (
            O => \N__26874\,
            I => \N__26871\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__26871\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__26868\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\
        );

    \I__3429\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26860\
        );

    \I__3428\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26855\
        );

    \I__3427\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26855\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26852\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__26855\,
            I => \N__26849\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__26852\,
            I => \N__26846\
        );

    \I__3423\ : Span4Mux_v
    port map (
            O => \N__26849\,
            I => \N__26843\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__26846\,
            I => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__26843\,
            I => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\
        );

    \I__3420\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__26835\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__26832\,
            I => \pid_alt.un1_pid_prereg_236_1_cascade_\
        );

    \I__3417\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26825\
        );

    \I__3416\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26822\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26819\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__26822\,
            I => \pid_alt.error_d_reg_prevZ0Z_8\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__26819\,
            I => \pid_alt.error_d_reg_prevZ0Z_8\
        );

    \I__3412\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26810\
        );

    \I__3411\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26807\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__26810\,
            I => \N__26804\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__26807\,
            I => \N__26801\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__26804\,
            I => \N__26798\
        );

    \I__3407\ : Span4Mux_h
    port map (
            O => \N__26801\,
            I => \N__26795\
        );

    \I__3406\ : Span4Mux_v
    port map (
            O => \N__26798\,
            I => \N__26792\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__26795\,
            I => \pid_alt.error_p_regZ0Z_8\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__26792\,
            I => \pid_alt.error_p_regZ0Z_8\
        );

    \I__3403\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26781\
        );

    \I__3402\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26781\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26777\
        );

    \I__3400\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26774\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__26777\,
            I => \N__26769\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__26774\,
            I => \N__26769\
        );

    \I__3397\ : Span4Mux_v
    port map (
            O => \N__26769\,
            I => \N__26766\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__26763\,
            I => \pid_alt.error_d_regZ0Z_8\
        );

    \I__3394\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26754\
        );

    \I__3393\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26754\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__26754\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__26751\,
            I => \N__26747\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__26750\,
            I => \N__26744\
        );

    \I__3389\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26741\
        );

    \I__3388\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26738\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__26741\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__26738\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\
        );

    \I__3385\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26724\
        );

    \I__3384\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26724\
        );

    \I__3383\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26724\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__26724\,
            I => \N__26721\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__26721\,
            I => \N__26718\
        );

    \I__3380\ : Span4Mux_v
    port map (
            O => \N__26718\,
            I => \N__26715\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__26715\,
            I => \pid_alt.error_d_regZ0Z_7\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__3377\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26703\
        );

    \I__3376\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26703\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__26703\,
            I => \pid_alt.error_d_reg_prevZ0Z_7\
        );

    \I__3374\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26694\
        );

    \I__3373\ : InMux
    port map (
            O => \N__26699\,
            I => \N__26694\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__3371\ : Span4Mux_h
    port map (
            O => \N__26691\,
            I => \N__26688\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__26688\,
            I => \pid_alt.error_p_regZ0Z_7\
        );

    \I__3369\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26682\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__26682\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\
        );

    \I__3367\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26673\
        );

    \I__3366\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26673\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__3364\ : Span4Mux_v
    port map (
            O => \N__26670\,
            I => \N__26667\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__26667\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\
        );

    \I__3362\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26660\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__26663\,
            I => \N__26657\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__26660\,
            I => \N__26654\
        );

    \I__3359\ : InMux
    port map (
            O => \N__26657\,
            I => \N__26651\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__26654\,
            I => \N__26648\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__26651\,
            I => \N__26645\
        );

    \I__3356\ : Span4Mux_v
    port map (
            O => \N__26648\,
            I => \N__26642\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__26645\,
            I => \N__26639\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__26642\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__26639\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__26634\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_\
        );

    \I__3351\ : InMux
    port map (
            O => \N__26631\,
            I => \N__26625\
        );

    \I__3350\ : InMux
    port map (
            O => \N__26630\,
            I => \N__26625\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__26625\,
            I => \N__26621\
        );

    \I__3348\ : InMux
    port map (
            O => \N__26624\,
            I => \N__26618\
        );

    \I__3347\ : Span4Mux_v
    port map (
            O => \N__26621\,
            I => \N__26615\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__26618\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__26615\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\
        );

    \I__3344\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__26607\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__3341\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__26598\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\
        );

    \I__3339\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__26592\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__26589\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_\
        );

    \I__3336\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26581\
        );

    \I__3335\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26576\
        );

    \I__3334\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26576\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26573\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__26576\,
            I => \N__26570\
        );

    \I__3331\ : Span4Mux_v
    port map (
            O => \N__26573\,
            I => \N__26565\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__26570\,
            I => \N__26565\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__26565\,
            I => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__26562\,
            I => \N__26558\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__26561\,
            I => \N__26555\
        );

    \I__3326\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26552\
        );

    \I__3325\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26549\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__26552\,
            I => \N__26546\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26543\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__26546\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__26543\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\
        );

    \I__3320\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26535\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__26535\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__26532\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_\
        );

    \I__3317\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26526\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__26526\,
            I => \N__26521\
        );

    \I__3315\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26516\
        );

    \I__3314\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26516\
        );

    \I__3313\ : Span4Mux_v
    port map (
            O => \N__26521\,
            I => \N__26511\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__26516\,
            I => \N__26511\
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__26511\,
            I => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\
        );

    \I__3310\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26502\
        );

    \I__3309\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26502\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__26502\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\
        );

    \I__3307\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26493\
        );

    \I__3306\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26493\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__26493\,
            I => \N__26490\
        );

    \I__3304\ : Span4Mux_v
    port map (
            O => \N__26490\,
            I => \N__26487\
        );

    \I__3303\ : Span4Mux_h
    port map (
            O => \N__26487\,
            I => \N__26484\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__26484\,
            I => \pid_alt.error_p_regZ0Z_14\
        );

    \I__3301\ : InMux
    port map (
            O => \N__26481\,
            I => \N__26475\
        );

    \I__3300\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26475\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__26475\,
            I => \N__26472\
        );

    \I__3298\ : Span4Mux_v
    port map (
            O => \N__26472\,
            I => \N__26469\
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__26469\,
            I => \pid_alt.error_d_reg_prevZ0Z_14\
        );

    \I__3296\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__26463\,
            I => \N__26458\
        );

    \I__3294\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26455\
        );

    \I__3293\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26452\
        );

    \I__3292\ : Sp12to4
    port map (
            O => \N__26458\,
            I => \N__26445\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__26455\,
            I => \N__26445\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26445\
        );

    \I__3289\ : Span12Mux_v
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__3288\ : Odrv12
    port map (
            O => \N__26442\,
            I => \pid_alt.error_d_regZ0Z_14\
        );

    \I__3287\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26435\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__26438\,
            I => \N__26432\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__26435\,
            I => \N__26429\
        );

    \I__3284\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26426\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__26429\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__26426\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__26421\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\
        );

    \I__3280\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26415\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__26415\,
            I => \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\
        );

    \I__3278\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26409\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__26409\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\
        );

    \I__3276\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26400\
        );

    \I__3275\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26400\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__26400\,
            I => \N__26397\
        );

    \I__3273\ : Span4Mux_v
    port map (
            O => \N__26397\,
            I => \N__26394\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__26394\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\
        );

    \I__3271\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26388\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26383\
        );

    \I__3269\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26378\
        );

    \I__3268\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26378\
        );

    \I__3267\ : Span4Mux_v
    port map (
            O => \N__26383\,
            I => \N__26373\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__26378\,
            I => \N__26373\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__26373\,
            I => \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__26370\,
            I => \N__26367\
        );

    \I__3263\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26363\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__26366\,
            I => \N__26360\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__26363\,
            I => \N__26357\
        );

    \I__3260\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26354\
        );

    \I__3259\ : Span4Mux_h
    port map (
            O => \N__26357\,
            I => \N__26351\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__26354\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__26351\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\
        );

    \I__3256\ : InMux
    port map (
            O => \N__26346\,
            I => \N__26343\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__26343\,
            I => \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\
        );

    \I__3254\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__26337\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__26334\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\
        );

    \I__3251\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26327\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__26330\,
            I => \N__26324\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__26327\,
            I => \N__26321\
        );

    \I__3248\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26318\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__26321\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__26318\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\
        );

    \I__3245\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__26310\,
            I => \N__26306\
        );

    \I__3243\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26303\
        );

    \I__3242\ : Span4Mux_v
    port map (
            O => \N__26306\,
            I => \N__26300\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__26303\,
            I => \N__26297\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__26300\,
            I => \N__26294\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__26297\,
            I => \N__26291\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__26294\,
            I => \pid_alt.error_p_regZ0Z_10\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__26291\,
            I => \pid_alt.error_p_regZ0Z_10\
        );

    \I__3236\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26283\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__26283\,
            I => \N__26279\
        );

    \I__3234\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26276\
        );

    \I__3233\ : Odrv12
    port map (
            O => \N__26279\,
            I => \pid_alt.error_d_reg_prevZ0Z_10\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__26276\,
            I => \pid_alt.error_d_reg_prevZ0Z_10\
        );

    \I__3231\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26266\
        );

    \I__3230\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26261\
        );

    \I__3229\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26261\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__26266\,
            I => \N__26258\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26255\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__26258\,
            I => \N__26252\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__26255\,
            I => \N__26249\
        );

    \I__3224\ : Span4Mux_v
    port map (
            O => \N__26252\,
            I => \N__26246\
        );

    \I__3223\ : Span4Mux_v
    port map (
            O => \N__26249\,
            I => \N__26243\
        );

    \I__3222\ : Span4Mux_v
    port map (
            O => \N__26246\,
            I => \N__26240\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__26243\,
            I => \N__26237\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__26240\,
            I => \pid_alt.error_d_regZ0Z_10\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__26237\,
            I => \pid_alt.error_d_regZ0Z_10\
        );

    \I__3218\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26229\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__26226\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__26223\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_\
        );

    \I__3214\ : InMux
    port map (
            O => \N__26220\,
            I => \N__26217\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__26217\,
            I => \N__26214\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__26214\,
            I => \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\
        );

    \I__3211\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26207\
        );

    \I__3210\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26204\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__26207\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__26204\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\
        );

    \I__3207\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26196\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__26196\,
            I => \N__26193\
        );

    \I__3205\ : Span12Mux_s4_h
    port map (
            O => \N__26193\,
            I => \N__26190\
        );

    \I__3204\ : Odrv12
    port map (
            O => \N__26190\,
            I => drone_altitude_i_11
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__26187\,
            I => \N__26184\
        );

    \I__3202\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26180\
        );

    \I__3201\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26177\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26174\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__26177\,
            I => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__26174\,
            I => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\
        );

    \I__3197\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26164\
        );

    \I__3196\ : InMux
    port map (
            O => \N__26168\,
            I => \N__26159\
        );

    \I__3195\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26159\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__26164\,
            I => \N__26154\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__26159\,
            I => \N__26154\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__26154\,
            I => \N__26151\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__26151\,
            I => \pid_alt.error_d_regZ0Z_9\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__26148\,
            I => \N__26145\
        );

    \I__3189\ : InMux
    port map (
            O => \N__26145\,
            I => \N__26139\
        );

    \I__3188\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26139\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__26139\,
            I => \N__26136\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__26136\,
            I => \pid_alt.error_d_reg_prevZ0Z_9\
        );

    \I__3185\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26127\
        );

    \I__3184\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26127\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__26127\,
            I => \N__26124\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__26124\,
            I => \N__26121\
        );

    \I__3181\ : Span4Mux_v
    port map (
            O => \N__26121\,
            I => \N__26118\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__26118\,
            I => \pid_alt.error_p_regZ0Z_9\
        );

    \I__3179\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26112\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__26112\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\
        );

    \I__3177\ : InMux
    port map (
            O => \N__26109\,
            I => \N__26103\
        );

    \I__3176\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26103\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__26103\,
            I => \N__26100\
        );

    \I__3174\ : Span4Mux_v
    port map (
            O => \N__26100\,
            I => \N__26097\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__26097\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__26094\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\
        );

    \I__3171\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26088\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__26088\,
            I => \N__26085\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__26085\,
            I => \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\
        );

    \I__3168\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26079\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__3166\ : Span4Mux_v
    port map (
            O => \N__26076\,
            I => \N__26073\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__26073\,
            I => \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__26070\,
            I => \N__26067\
        );

    \I__3163\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26063\
        );

    \I__3162\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26060\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__26063\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__26060\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__26055\,
            I => \N__26052\
        );

    \I__3158\ : InMux
    port map (
            O => \N__26052\,
            I => \N__26048\
        );

    \I__3157\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26045\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__26048\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__26045\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__3154\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26036\
        );

    \I__3153\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26033\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__26036\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__26033\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__26028\,
            I => \N__26025\
        );

    \I__3149\ : InMux
    port map (
            O => \N__26025\,
            I => \N__26021\
        );

    \I__3148\ : InMux
    port map (
            O => \N__26024\,
            I => \N__26018\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__26021\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__26018\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__26013\,
            I => \N__26010\
        );

    \I__3144\ : InMux
    port map (
            O => \N__26010\,
            I => \N__26006\
        );

    \I__3143\ : InMux
    port map (
            O => \N__26009\,
            I => \N__26003\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__26006\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__26003\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__3140\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25994\
        );

    \I__3139\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25991\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__25994\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__25991\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__3136\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25983\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__25983\,
            I => \N__25980\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__25980\,
            I => \pid_alt.m35_e_2\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__25977\,
            I => \N__25974\
        );

    \I__3132\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25970\
        );

    \I__3131\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25967\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__25970\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__25967\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__3128\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25959\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__25959\,
            I => \N__25956\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__25956\,
            I => \N__25953\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__25953\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\
        );

    \I__3124\ : InMux
    port map (
            O => \N__25950\,
            I => \N__25947\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25943\
        );

    \I__3122\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25940\
        );

    \I__3121\ : Span4Mux_v
    port map (
            O => \N__25943\,
            I => \N__25937\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__25940\,
            I => \N__25934\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__25937\,
            I => \N__25931\
        );

    \I__3118\ : Span4Mux_v
    port map (
            O => \N__25934\,
            I => \N__25928\
        );

    \I__3117\ : Odrv4
    port map (
            O => \N__25931\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__25928\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11\
        );

    \I__3115\ : InMux
    port map (
            O => \N__25923\,
            I => \N__25919\
        );

    \I__3114\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25915\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25912\
        );

    \I__3112\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25909\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__25915\,
            I => \N__25906\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__25912\,
            I => \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__25909\,
            I => \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__25906\,
            I => \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__25899\,
            I => \N__25895\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__25898\,
            I => \N__25892\
        );

    \I__3105\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25889\
        );

    \I__3104\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25886\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__25889\,
            I => \N__25883\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__25886\,
            I => \N__25880\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__25883\,
            I => \N__25877\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__25880\,
            I => \N__25874\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__25877\,
            I => \pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__25874\,
            I => \pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11\
        );

    \I__3097\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25865\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__25868\,
            I => \N__25862\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__25865\,
            I => \N__25858\
        );

    \I__3094\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25855\
        );

    \I__3093\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25852\
        );

    \I__3092\ : Span12Mux_s3_h
    port map (
            O => \N__25858\,
            I => \N__25847\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25847\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__25852\,
            I => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\
        );

    \I__3089\ : Odrv12
    port map (
            O => \N__25847\,
            I => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\
        );

    \I__3088\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25839\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__25839\,
            I => \pid_alt.error_i_acummZ0Z_3\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__25836\,
            I => \N__25833\
        );

    \I__3085\ : InMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__25827\,
            I => \pid_alt.error_i_acummZ0Z_1\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__25824\,
            I => \pid_alt.N_9_0_cascade_\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__25821\,
            I => \pid_alt.N_62_mux_cascade_\
        );

    \I__3080\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__25815\,
            I => \N__25811\
        );

    \I__3078\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25808\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__25811\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__25808\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__3075\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__25800\,
            I => \pid_alt.error_i_acummZ0Z_4\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__25797\,
            I => \N__25793\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__25796\,
            I => \N__25789\
        );

    \I__3071\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25779\
        );

    \I__3070\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25779\
        );

    \I__3069\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25779\
        );

    \I__3068\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25779\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__25779\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3Z0Z_5\
        );

    \I__3066\ : InMux
    port map (
            O => \N__25776\,
            I => \N__25773\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__25773\,
            I => \pid_alt.error_i_acummZ0Z_2\
        );

    \I__3064\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25767\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__25767\,
            I => \pid_alt.error_i_acumm_preregZ0Z_16\
        );

    \I__3062\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25761\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__25761\,
            I => \pid_alt.error_i_acumm_preregZ0Z_17\
        );

    \I__3060\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25755\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__25755\,
            I => \pid_alt.error_i_acumm_preregZ0Z_14\
        );

    \I__3058\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25749\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__25749\,
            I => \pid_alt.error_i_acumm_preregZ0Z_15\
        );

    \I__3056\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25741\
        );

    \I__3055\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25736\
        );

    \I__3054\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25736\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__25741\,
            I => \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__25736\,
            I => \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__25731\,
            I => \N__25728\
        );

    \I__3050\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25723\
        );

    \I__3049\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25720\
        );

    \I__3048\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25717\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__25723\,
            I => \N__25714\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__25720\,
            I => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__25717\,
            I => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__25714\,
            I => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\
        );

    \I__3043\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25702\
        );

    \I__3042\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25697\
        );

    \I__3041\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25697\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__25702\,
            I => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__25697\,
            I => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\
        );

    \I__3038\ : InMux
    port map (
            O => \N__25692\,
            I => \N__25689\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__25689\,
            I => \N__25686\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__25686\,
            I => \N__25683\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__25683\,
            I => alt_kp_2
        );

    \I__3034\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__25677\,
            I => \N__25674\
        );

    \I__3032\ : Span4Mux_s3_h
    port map (
            O => \N__25674\,
            I => \N__25671\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__25671\,
            I => alt_kp_5
        );

    \I__3030\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25664\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__25667\,
            I => \N__25661\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__25664\,
            I => \N__25658\
        );

    \I__3027\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25655\
        );

    \I__3026\ : Span4Mux_h
    port map (
            O => \N__25658\,
            I => \N__25652\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__25655\,
            I => \Commands_frame_decoder.stateZ0Z_2\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__25652\,
            I => \Commands_frame_decoder.stateZ0Z_2\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__3022\ : InMux
    port map (
            O => \N__25644\,
            I => \N__25640\
        );

    \I__3021\ : InMux
    port map (
            O => \N__25643\,
            I => \N__25637\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__25640\,
            I => \N__25634\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__25637\,
            I => \N__25631\
        );

    \I__3018\ : Span4Mux_v
    port map (
            O => \N__25634\,
            I => \N__25628\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__25631\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__25628\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__3015\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__25620\,
            I => \pid_alt.error_i_acumm_preregZ0Z_18\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__3012\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__25611\,
            I => \pid_alt.error_i_acumm_preregZ0Z_19\
        );

    \I__3010\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25605\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__25605\,
            I => \pid_alt.error_i_acumm_preregZ0Z_20\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__25602\,
            I => \pid_alt.m7_e_4_cascade_\
        );

    \I__3007\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25595\
        );

    \I__3006\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25592\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__25592\,
            I => \N__25586\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__25589\,
            I => \N__25583\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__25586\,
            I => \N__25580\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__25583\,
            I => \pid_alt.error_p_regZ0Z_13\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__25580\,
            I => \pid_alt.error_p_regZ0Z_13\
        );

    \I__2999\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25569\
        );

    \I__2998\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25569\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__25569\,
            I => \N__25566\
        );

    \I__2996\ : Span4Mux_h
    port map (
            O => \N__25566\,
            I => \N__25562\
        );

    \I__2995\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25559\
        );

    \I__2994\ : Span4Mux_v
    port map (
            O => \N__25562\,
            I => \N__25556\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__25559\,
            I => \N__25553\
        );

    \I__2992\ : Sp12to4
    port map (
            O => \N__25556\,
            I => \N__25548\
        );

    \I__2991\ : Span12Mux_s5_h
    port map (
            O => \N__25553\,
            I => \N__25548\
        );

    \I__2990\ : Span12Mux_v
    port map (
            O => \N__25548\,
            I => \N__25545\
        );

    \I__2989\ : Odrv12
    port map (
            O => \N__25545\,
            I => \pid_alt.error_d_regZ0Z_13\
        );

    \I__2988\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25539\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__25539\,
            I => \N__25535\
        );

    \I__2986\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25532\
        );

    \I__2985\ : Span4Mux_s3_h
    port map (
            O => \N__25535\,
            I => \N__25529\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__25532\,
            I => \pid_alt.error_d_reg_prevZ0Z_13\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__25529\,
            I => \pid_alt.error_d_reg_prevZ0Z_13\
        );

    \I__2982\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__25521\,
            I => \N__25518\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__25518\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__2978\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25509\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__25509\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__25506\,
            I => \N__25503\
        );

    \I__2975\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25499\
        );

    \I__2974\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25496\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__25499\,
            I => \N__25493\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__25496\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\
        );

    \I__2971\ : Odrv4
    port map (
            O => \N__25493\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\
        );

    \I__2970\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25485\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__25485\,
            I => \dron_frame_decoder_1.drone_altitude_10\
        );

    \I__2968\ : InMux
    port map (
            O => \N__25482\,
            I => \pid_alt.un1_pid_prereg_0_cry_15\
        );

    \I__2967\ : InMux
    port map (
            O => \N__25479\,
            I => \pid_alt.un1_pid_prereg_0_cry_16\
        );

    \I__2966\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__25473\,
            I => \N__25470\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__25470\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\
        );

    \I__2963\ : InMux
    port map (
            O => \N__25467\,
            I => \pid_alt.un1_pid_prereg_0_cry_17\
        );

    \I__2962\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25461\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__25461\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__25458\,
            I => \N__25454\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__25457\,
            I => \N__25451\
        );

    \I__2958\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25448\
        );

    \I__2957\ : InMux
    port map (
            O => \N__25451\,
            I => \N__25445\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__25448\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__25445\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\
        );

    \I__2954\ : InMux
    port map (
            O => \N__25440\,
            I => \pid_alt.un1_pid_prereg_0_cry_18\
        );

    \I__2953\ : InMux
    port map (
            O => \N__25437\,
            I => \pid_alt.un1_pid_prereg_0_cry_19\
        );

    \I__2952\ : InMux
    port map (
            O => \N__25434\,
            I => \pid_alt.un1_pid_prereg_0_cry_20\
        );

    \I__2951\ : InMux
    port map (
            O => \N__25431\,
            I => \pid_alt.un1_pid_prereg_0_cry_21\
        );

    \I__2950\ : InMux
    port map (
            O => \N__25428\,
            I => \bfn_3_20_0_\
        );

    \I__2949\ : InMux
    port map (
            O => \N__25425\,
            I => \pid_alt.un1_pid_prereg_0_cry_23\
        );

    \I__2948\ : InMux
    port map (
            O => \N__25422\,
            I => \bfn_3_18_0_\
        );

    \I__2947\ : InMux
    port map (
            O => \N__25419\,
            I => \pid_alt.un1_pid_prereg_0_cry_7\
        );

    \I__2946\ : InMux
    port map (
            O => \N__25416\,
            I => \pid_alt.un1_pid_prereg_0_cry_8\
        );

    \I__2945\ : InMux
    port map (
            O => \N__25413\,
            I => \pid_alt.un1_pid_prereg_0_cry_9\
        );

    \I__2944\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__25407\,
            I => \N__25404\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__25404\,
            I => \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__25401\,
            I => \N__25397\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__25400\,
            I => \N__25394\
        );

    \I__2939\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25391\
        );

    \I__2938\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25388\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__25391\,
            I => \N__25385\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__25388\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__25385\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\
        );

    \I__2934\ : InMux
    port map (
            O => \N__25380\,
            I => \pid_alt.un1_pid_prereg_0_cry_10\
        );

    \I__2933\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__25374\,
            I => \pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__25371\,
            I => \N__25368\
        );

    \I__2930\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25364\
        );

    \I__2929\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25361\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__25364\,
            I => \N__25358\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__25361\,
            I => \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__25358\,
            I => \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\
        );

    \I__2925\ : InMux
    port map (
            O => \N__25353\,
            I => \pid_alt.un1_pid_prereg_0_cry_11\
        );

    \I__2924\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25347\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__25347\,
            I => \pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12\
        );

    \I__2922\ : InMux
    port map (
            O => \N__25344\,
            I => \pid_alt.un1_pid_prereg_0_cry_12\
        );

    \I__2921\ : InMux
    port map (
            O => \N__25341\,
            I => \pid_alt.un1_pid_prereg_0_cry_13\
        );

    \I__2920\ : InMux
    port map (
            O => \N__25338\,
            I => \bfn_3_19_0_\
        );

    \I__2919\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25332\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__25332\,
            I => \N__25329\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__25329\,
            I => \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__25326\,
            I => \N__25323\
        );

    \I__2915\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25320\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__25320\,
            I => \N__25316\
        );

    \I__2913\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25313\
        );

    \I__2912\ : Span4Mux_v
    port map (
            O => \N__25316\,
            I => \N__25310\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__25313\,
            I => \pid_alt.un1_pid_prereg_0\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__25310\,
            I => \pid_alt.un1_pid_prereg_0\
        );

    \I__2909\ : InMux
    port map (
            O => \N__25305\,
            I => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\
        );

    \I__2908\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25299\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__25299\,
            I => \N__25296\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__25296\,
            I => \N__25293\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__25293\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__25290\,
            I => \N__25286\
        );

    \I__2903\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25283\
        );

    \I__2902\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25280\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__25283\,
            I => \N__25275\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25275\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__25275\,
            I => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\
        );

    \I__2898\ : InMux
    port map (
            O => \N__25272\,
            I => \pid_alt.un1_pid_prereg_0_cry_0\
        );

    \I__2897\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25266\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__25266\,
            I => \N__25263\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__25263\,
            I => \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1\
        );

    \I__2894\ : InMux
    port map (
            O => \N__25260\,
            I => \pid_alt.un1_pid_prereg_0_cry_1\
        );

    \I__2893\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25254\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__25254\,
            I => \N__25251\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__25248\,
            I => \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\
        );

    \I__2889\ : InMux
    port map (
            O => \N__25245\,
            I => \pid_alt.un1_pid_prereg_0_cry_2\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__2887\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25235\
        );

    \I__2886\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25232\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__25235\,
            I => \N__25229\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__25232\,
            I => \N__25226\
        );

    \I__2883\ : Span4Mux_v
    port map (
            O => \N__25229\,
            I => \N__25221\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__25226\,
            I => \N__25221\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__25221\,
            I => \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__25218\,
            I => \N__25215\
        );

    \I__2879\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25212\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__25212\,
            I => \N__25209\
        );

    \I__2877\ : Odrv12
    port map (
            O => \N__25209\,
            I => \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3\
        );

    \I__2876\ : InMux
    port map (
            O => \N__25206\,
            I => \pid_alt.un1_pid_prereg_0_cry_3\
        );

    \I__2875\ : InMux
    port map (
            O => \N__25203\,
            I => \N__25200\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__25200\,
            I => \N__25197\
        );

    \I__2873\ : Odrv12
    port map (
            O => \N__25197\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__25194\,
            I => \N__25191\
        );

    \I__2871\ : InMux
    port map (
            O => \N__25191\,
            I => \N__25188\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__25188\,
            I => \N__25184\
        );

    \I__2869\ : InMux
    port map (
            O => \N__25187\,
            I => \N__25181\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__25184\,
            I => \N__25178\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__25181\,
            I => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\
        );

    \I__2866\ : Odrv4
    port map (
            O => \N__25178\,
            I => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\
        );

    \I__2865\ : InMux
    port map (
            O => \N__25173\,
            I => \pid_alt.un1_pid_prereg_0_cry_4\
        );

    \I__2864\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25167\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__25167\,
            I => \N__25164\
        );

    \I__2862\ : Span4Mux_v
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__25161\,
            I => \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__25158\,
            I => \N__25154\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__25157\,
            I => \N__25151\
        );

    \I__2858\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25148\
        );

    \I__2857\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25145\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__25148\,
            I => \N__25142\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__25145\,
            I => \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\
        );

    \I__2854\ : Odrv12
    port map (
            O => \N__25142\,
            I => \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\
        );

    \I__2853\ : InMux
    port map (
            O => \N__25137\,
            I => \pid_alt.un1_pid_prereg_0_cry_5\
        );

    \I__2852\ : InMux
    port map (
            O => \N__25134\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_14\
        );

    \I__2851\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__25128\,
            I => \N__25125\
        );

    \I__2849\ : Span4Mux_v
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__25122\,
            I => \N__25119\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__25119\,
            I => \pid_alt.error_i_regZ0Z_16\
        );

    \I__2846\ : InMux
    port map (
            O => \N__25116\,
            I => \bfn_3_16_0_\
        );

    \I__2845\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__25110\,
            I => \N__25107\
        );

    \I__2843\ : Span4Mux_v
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__25104\,
            I => \N__25101\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__25101\,
            I => \pid_alt.error_i_regZ0Z_17\
        );

    \I__2840\ : InMux
    port map (
            O => \N__25098\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_16\
        );

    \I__2839\ : InMux
    port map (
            O => \N__25095\,
            I => \N__25092\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__25092\,
            I => \N__25089\
        );

    \I__2837\ : Span4Mux_v
    port map (
            O => \N__25089\,
            I => \N__25086\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__25086\,
            I => \N__25083\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__25083\,
            I => \pid_alt.error_i_regZ0Z_18\
        );

    \I__2834\ : InMux
    port map (
            O => \N__25080\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_17\
        );

    \I__2833\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25074\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__25071\,
            I => \N__25068\
        );

    \I__2830\ : Span4Mux_v
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__25065\,
            I => \pid_alt.error_i_regZ0Z_19\
        );

    \I__2828\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25057\
        );

    \I__2827\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25052\
        );

    \I__2826\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25052\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__25057\,
            I => \N__25049\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25046\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__25049\,
            I => \N__25043\
        );

    \I__2822\ : Span4Mux_v
    port map (
            O => \N__25046\,
            I => \N__25040\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__25043\,
            I => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__25040\,
            I => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\
        );

    \I__2819\ : InMux
    port map (
            O => \N__25035\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_18\
        );

    \I__2818\ : InMux
    port map (
            O => \N__25032\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19\
        );

    \I__2817\ : InMux
    port map (
            O => \N__25029\,
            I => \N__25023\
        );

    \I__2816\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25023\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__2814\ : Span4Mux_h
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__25014\,
            I => \pid_alt.error_i_regZ0Z_20\
        );

    \I__2811\ : InMux
    port map (
            O => \N__25011\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20\
        );

    \I__2810\ : InMux
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__24999\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\
        );

    \I__2806\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24992\
        );

    \I__2805\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24989\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__24992\,
            I => \N__24986\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24982\
        );

    \I__2802\ : Span4Mux_v
    port map (
            O => \N__24986\,
            I => \N__24979\
        );

    \I__2801\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24976\
        );

    \I__2800\ : Odrv12
    port map (
            O => \N__24982\,
            I => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__24979\,
            I => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__24976\,
            I => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__2796\ : InMux
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__2794\ : Span4Mux_v
    port map (
            O => \N__24960\,
            I => \N__24957\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__24957\,
            I => \pid_alt.error_i_regZ0Z_7\
        );

    \I__2792\ : InMux
    port map (
            O => \N__24954\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__2790\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__24945\,
            I => \N__24942\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__24942\,
            I => \N__24939\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__24939\,
            I => \pid_alt.error_i_regZ0Z_8\
        );

    \I__2786\ : InMux
    port map (
            O => \N__24936\,
            I => \bfn_3_15_0_\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__24933\,
            I => \N__24930\
        );

    \I__2784\ : InMux
    port map (
            O => \N__24930\,
            I => \N__24927\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24924\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__24924\,
            I => \N__24921\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__24921\,
            I => \pid_alt.error_i_regZ0Z_9\
        );

    \I__2780\ : InMux
    port map (
            O => \N__24918\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__24915\,
            I => \N__24912\
        );

    \I__2778\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__2776\ : Span4Mux_v
    port map (
            O => \N__24906\,
            I => \N__24903\
        );

    \I__2775\ : Span4Mux_v
    port map (
            O => \N__24903\,
            I => \N__24900\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__24900\,
            I => \pid_alt.error_i_regZ0Z_10\
        );

    \I__2773\ : InMux
    port map (
            O => \N__24897\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__24894\,
            I => \N__24891\
        );

    \I__2771\ : InMux
    port map (
            O => \N__24891\,
            I => \N__24888\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__24888\,
            I => \N__24885\
        );

    \I__2769\ : Odrv12
    port map (
            O => \N__24885\,
            I => \pid_alt.error_i_regZ0Z_11\
        );

    \I__2768\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24873\
        );

    \I__2767\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24873\
        );

    \I__2766\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24873\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__24873\,
            I => \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\
        );

    \I__2764\ : InMux
    port map (
            O => \N__24870\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_10\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__2762\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__24858\,
            I => \N__24855\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__24855\,
            I => \pid_alt.error_i_regZ0Z_12\
        );

    \I__2758\ : InMux
    port map (
            O => \N__24852\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_11\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__24849\,
            I => \N__24846\
        );

    \I__2756\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__24843\,
            I => \N__24840\
        );

    \I__2754\ : Span4Mux_h
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__2753\ : Span4Mux_v
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__24834\,
            I => \pid_alt.error_i_regZ0Z_13\
        );

    \I__2751\ : InMux
    port map (
            O => \N__24831\,
            I => \N__24826\
        );

    \I__2750\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24821\
        );

    \I__2749\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24821\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24818\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__24821\,
            I => \N__24815\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__24818\,
            I => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__24815\,
            I => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\
        );

    \I__2744\ : InMux
    port map (
            O => \N__24810\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_12\
        );

    \I__2743\ : InMux
    port map (
            O => \N__24807\,
            I => \N__24804\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__2741\ : Span4Mux_v
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__24798\,
            I => \pid_alt.error_i_regZ0Z_14\
        );

    \I__2739\ : InMux
    port map (
            O => \N__24795\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_13\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__2737\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__24780\,
            I => \pid_alt.error_i_regZ0Z_15\
        );

    \I__2733\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24774\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__24774\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\
        );

    \I__2731\ : InMux
    port map (
            O => \N__24771\,
            I => \N__24765\
        );

    \I__2730\ : InMux
    port map (
            O => \N__24770\,
            I => \N__24765\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__24765\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\
        );

    \I__2728\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24759\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__24759\,
            I => \pid_alt.error_i_regZ0Z_1\
        );

    \I__2726\ : InMux
    port map (
            O => \N__24756\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_0\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__2724\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24744\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__24744\,
            I => \N__24741\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__24741\,
            I => \pid_alt.error_i_regZ0Z_2\
        );

    \I__2720\ : InMux
    port map (
            O => \N__24738\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_1\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__24735\,
            I => \N__24732\
        );

    \I__2718\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24729\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__24729\,
            I => \N__24726\
        );

    \I__2716\ : Odrv12
    port map (
            O => \N__24726\,
            I => \pid_alt.error_i_regZ0Z_3\
        );

    \I__2715\ : InMux
    port map (
            O => \N__24723\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_2\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__24720\,
            I => \N__24717\
        );

    \I__2713\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__2711\ : Span4Mux_h
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__2710\ : Span4Mux_v
    port map (
            O => \N__24708\,
            I => \N__24705\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__24705\,
            I => \pid_alt.error_i_regZ0Z_4\
        );

    \I__2708\ : InMux
    port map (
            O => \N__24702\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_3\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__24699\,
            I => \N__24696\
        );

    \I__2706\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24693\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__24693\,
            I => \N__24690\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__24690\,
            I => \N__24687\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__24687\,
            I => \pid_alt.error_i_regZ0Z_5\
        );

    \I__2702\ : InMux
    port map (
            O => \N__24684\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_4\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__24681\,
            I => \N__24678\
        );

    \I__2700\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24675\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__24675\,
            I => \N__24672\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__24672\,
            I => \N__24669\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__24669\,
            I => \pid_alt.error_i_regZ0Z_6\
        );

    \I__2696\ : InMux
    port map (
            O => \N__24666\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5\
        );

    \I__2695\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24658\
        );

    \I__2694\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24655\
        );

    \I__2693\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24652\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__24658\,
            I => \N__24649\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__24655\,
            I => \N__24646\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__24652\,
            I => \N__24641\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__24649\,
            I => \N__24641\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__24646\,
            I => \N__24638\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__24641\,
            I => \N__24635\
        );

    \I__2686\ : Span4Mux_v
    port map (
            O => \N__24638\,
            I => \N__24632\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__24635\,
            I => \pid_alt.error_p_regZ0Z_3\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__24632\,
            I => \pid_alt.error_p_regZ0Z_3\
        );

    \I__2683\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24622\
        );

    \I__2682\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24619\
        );

    \I__2681\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24616\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__24622\,
            I => \pid_alt.error_d_reg_prevZ0Z_3\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__24619\,
            I => \pid_alt.error_d_reg_prevZ0Z_3\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__24616\,
            I => \pid_alt.error_d_reg_prevZ0Z_3\
        );

    \I__2677\ : InMux
    port map (
            O => \N__24609\,
            I => \N__24605\
        );

    \I__2676\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24601\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__24605\,
            I => \N__24597\
        );

    \I__2674\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24594\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__24601\,
            I => \N__24591\
        );

    \I__2672\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24588\
        );

    \I__2671\ : Span4Mux_h
    port map (
            O => \N__24597\,
            I => \N__24585\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__24594\,
            I => \N__24578\
        );

    \I__2669\ : Span4Mux_h
    port map (
            O => \N__24591\,
            I => \N__24578\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24578\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__24585\,
            I => \N__24575\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__24578\,
            I => \N__24572\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__24575\,
            I => \pid_alt.error_d_regZ0Z_3\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__24572\,
            I => \pid_alt.error_d_regZ0Z_3\
        );

    \I__2663\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24564\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__24564\,
            I => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__24561\,
            I => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_\
        );

    \I__2660\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24552\
        );

    \I__2659\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24552\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__24552\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\
        );

    \I__2657\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24543\
        );

    \I__2656\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24543\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__24543\,
            I => \N__24540\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__24537\,
            I => \N__24534\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__24534\,
            I => \N__24531\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__24531\,
            I => \pid_alt.error_p_regZ0Z_4\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__24528\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_\
        );

    \I__2649\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24516\
        );

    \I__2648\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24516\
        );

    \I__2647\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24516\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__2645\ : Odrv12
    port map (
            O => \N__24513\,
            I => \pid_alt.error_d_regZ0Z_4\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__24510\,
            I => \N__24507\
        );

    \I__2643\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24501\
        );

    \I__2642\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24501\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__24501\,
            I => \pid_alt.error_d_reg_prevZ0Z_4\
        );

    \I__2640\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__24495\,
            I => \N__24492\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__24492\,
            I => \N__24489\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__24489\,
            I => \pid_alt.O_4_4\
        );

    \I__2636\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24483\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__24483\,
            I => \N__24480\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__24480\,
            I => \N__24477\
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__24477\,
            I => \pid_alt.O_4_7\
        );

    \I__2632\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24471\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__24471\,
            I => \N__24468\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__24468\,
            I => \N__24465\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__24465\,
            I => \pid_alt.O_4_15\
        );

    \I__2628\ : CEMux
    port map (
            O => \N__24462\,
            I => \N__24417\
        );

    \I__2627\ : CEMux
    port map (
            O => \N__24461\,
            I => \N__24417\
        );

    \I__2626\ : CEMux
    port map (
            O => \N__24460\,
            I => \N__24417\
        );

    \I__2625\ : CEMux
    port map (
            O => \N__24459\,
            I => \N__24417\
        );

    \I__2624\ : CEMux
    port map (
            O => \N__24458\,
            I => \N__24417\
        );

    \I__2623\ : CEMux
    port map (
            O => \N__24457\,
            I => \N__24417\
        );

    \I__2622\ : CEMux
    port map (
            O => \N__24456\,
            I => \N__24417\
        );

    \I__2621\ : CEMux
    port map (
            O => \N__24455\,
            I => \N__24417\
        );

    \I__2620\ : CEMux
    port map (
            O => \N__24454\,
            I => \N__24417\
        );

    \I__2619\ : CEMux
    port map (
            O => \N__24453\,
            I => \N__24417\
        );

    \I__2618\ : CEMux
    port map (
            O => \N__24452\,
            I => \N__24417\
        );

    \I__2617\ : CEMux
    port map (
            O => \N__24451\,
            I => \N__24417\
        );

    \I__2616\ : CEMux
    port map (
            O => \N__24450\,
            I => \N__24417\
        );

    \I__2615\ : CEMux
    port map (
            O => \N__24449\,
            I => \N__24417\
        );

    \I__2614\ : CEMux
    port map (
            O => \N__24448\,
            I => \N__24417\
        );

    \I__2613\ : GlobalMux
    port map (
            O => \N__24417\,
            I => \N__24414\
        );

    \I__2612\ : gio2CtrlBuf
    port map (
            O => \N__24414\,
            I => \pid_alt.N_664_0_g\
        );

    \I__2611\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24408\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__24408\,
            I => \N__24405\
        );

    \I__2609\ : Span4Mux_s3_h
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__24402\,
            I => \N__24399\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__24399\,
            I => \N__24396\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__24396\,
            I => \Commands_frame_decoder.source_CH1data8lt7_0\
        );

    \I__2605\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24384\
        );

    \I__2604\ : InMux
    port map (
            O => \N__24392\,
            I => \N__24384\
        );

    \I__2603\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24381\
        );

    \I__2602\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24378\
        );

    \I__2601\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24375\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__24384\,
            I => \N__24372\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__24381\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__24378\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__24375\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__24372\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2595\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24360\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__24360\,
            I => \N__24357\
        );

    \I__2593\ : Span4Mux_v
    port map (
            O => \N__24357\,
            I => \N__24354\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__24354\,
            I => \pid_alt.O_5_9\
        );

    \I__2591\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24345\
        );

    \I__2590\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24345\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24342\
        );

    \I__2588\ : Odrv12
    port map (
            O => \N__24342\,
            I => \pid_alt.error_p_regZ0Z_5\
        );

    \I__2587\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24336\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__24336\,
            I => \N__24333\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__24333\,
            I => \N__24330\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__24330\,
            I => \pid_alt.O_5_10\
        );

    \I__2583\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24321\
        );

    \I__2582\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24321\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__2580\ : Span12Mux_v
    port map (
            O => \N__24318\,
            I => \N__24315\
        );

    \I__2579\ : Odrv12
    port map (
            O => \N__24315\,
            I => \pid_alt.error_p_regZ0Z_6\
        );

    \I__2578\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24309\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__24309\,
            I => \N__24306\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__24306\,
            I => alt_kp_7
        );

    \I__2575\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24300\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24297\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__24297\,
            I => alt_kp_3
        );

    \I__2572\ : InMux
    port map (
            O => \N__24294\,
            I => \N__24291\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__24291\,
            I => \N__24288\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__24285\,
            I => \pid_alt.O_3_8\
        );

    \I__2568\ : CEMux
    port map (
            O => \N__24282\,
            I => \N__24279\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__24276\,
            I => \N__24272\
        );

    \I__2565\ : CEMux
    port map (
            O => \N__24275\,
            I => \N__24268\
        );

    \I__2564\ : Span4Mux_s0_h
    port map (
            O => \N__24272\,
            I => \N__24265\
        );

    \I__2563\ : CEMux
    port map (
            O => \N__24271\,
            I => \N__24262\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__24268\,
            I => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__24265\,
            I => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__24262\,
            I => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\
        );

    \I__2559\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24252\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__24252\,
            I => \N__24249\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__24249\,
            I => \N__24246\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__24246\,
            I => \pid_alt.O_3_11\
        );

    \I__2555\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24240\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24237\
        );

    \I__2553\ : Span4Mux_h
    port map (
            O => \N__24237\,
            I => \N__24234\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__24234\,
            I => \pid_alt.O_3_12\
        );

    \I__2551\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24228\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__24228\,
            I => \N__24225\
        );

    \I__2549\ : Span4Mux_h
    port map (
            O => \N__24225\,
            I => \N__24222\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__24222\,
            I => \pid_alt.O_3_13\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__24219\,
            I => \N__24216\
        );

    \I__2546\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24213\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__24213\,
            I => \N__24210\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__24210\,
            I => alt_command_7
        );

    \I__2543\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24202\
        );

    \I__2542\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24199\
        );

    \I__2541\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24196\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24193\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__24199\,
            I => \N__24190\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__24196\,
            I => \N__24187\
        );

    \I__2537\ : Span12Mux_s2_h
    port map (
            O => \N__24193\,
            I => \N__24184\
        );

    \I__2536\ : Span4Mux_s2_h
    port map (
            O => \N__24190\,
            I => \N__24181\
        );

    \I__2535\ : Span4Mux_s2_h
    port map (
            O => \N__24187\,
            I => \N__24178\
        );

    \I__2534\ : Span12Mux_v
    port map (
            O => \N__24184\,
            I => \N__24175\
        );

    \I__2533\ : Span4Mux_v
    port map (
            O => \N__24181\,
            I => \N__24172\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__24178\,
            I => \N__24169\
        );

    \I__2531\ : Odrv12
    port map (
            O => \N__24175\,
            I => \pid_alt.error_11\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__24172\,
            I => \pid_alt.error_11\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__24169\,
            I => \pid_alt.error_11\
        );

    \I__2528\ : InMux
    port map (
            O => \N__24162\,
            I => \pid_alt.error_cry_10\
        );

    \I__2527\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24156\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__24156\,
            I => \N__24153\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__24153\,
            I => \N__24148\
        );

    \I__2524\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24145\
        );

    \I__2523\ : InMux
    port map (
            O => \N__24151\,
            I => \N__24142\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__24148\,
            I => \N__24139\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__24145\,
            I => \N__24136\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__24142\,
            I => \N__24133\
        );

    \I__2519\ : Span4Mux_v
    port map (
            O => \N__24139\,
            I => \N__24130\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__24136\,
            I => \N__24127\
        );

    \I__2517\ : Span12Mux_s2_h
    port map (
            O => \N__24133\,
            I => \N__24124\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__24130\,
            I => \N__24119\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__24127\,
            I => \N__24119\
        );

    \I__2514\ : Odrv12
    port map (
            O => \N__24124\,
            I => \pid_alt.error_12\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__24119\,
            I => \pid_alt.error_12\
        );

    \I__2512\ : InMux
    port map (
            O => \N__24114\,
            I => \pid_alt.error_cry_11\
        );

    \I__2511\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24108\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24104\
        );

    \I__2509\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24101\
        );

    \I__2508\ : Span4Mux_s1_h
    port map (
            O => \N__24104\,
            I => \N__24097\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__24101\,
            I => \N__24094\
        );

    \I__2506\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24091\
        );

    \I__2505\ : Sp12to4
    port map (
            O => \N__24097\,
            I => \N__24088\
        );

    \I__2504\ : Span4Mux_s2_h
    port map (
            O => \N__24094\,
            I => \N__24085\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__24091\,
            I => \N__24082\
        );

    \I__2502\ : Span12Mux_v
    port map (
            O => \N__24088\,
            I => \N__24079\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__24085\,
            I => \N__24076\
        );

    \I__2500\ : Span12Mux_s2_h
    port map (
            O => \N__24082\,
            I => \N__24073\
        );

    \I__2499\ : Odrv12
    port map (
            O => \N__24079\,
            I => \pid_alt.error_13\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__24076\,
            I => \pid_alt.error_13\
        );

    \I__2497\ : Odrv12
    port map (
            O => \N__24073\,
            I => \pid_alt.error_13\
        );

    \I__2496\ : InMux
    port map (
            O => \N__24066\,
            I => \pid_alt.error_cry_12\
        );

    \I__2495\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24059\
        );

    \I__2494\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24055\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24052\
        );

    \I__2492\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24049\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__24055\,
            I => \N__24046\
        );

    \I__2490\ : Span12Mux_s7_v
    port map (
            O => \N__24052\,
            I => \N__24041\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24041\
        );

    \I__2488\ : Span4Mux_s2_h
    port map (
            O => \N__24046\,
            I => \N__24038\
        );

    \I__2487\ : Span12Mux_v
    port map (
            O => \N__24041\,
            I => \N__24035\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__24038\,
            I => \N__24032\
        );

    \I__2485\ : Odrv12
    port map (
            O => \N__24035\,
            I => \pid_alt.error_14\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__24032\,
            I => \pid_alt.error_14\
        );

    \I__2483\ : InMux
    port map (
            O => \N__24027\,
            I => \pid_alt.error_cry_13\
        );

    \I__2482\ : InMux
    port map (
            O => \N__24024\,
            I => \pid_alt.error_cry_14\
        );

    \I__2481\ : InMux
    port map (
            O => \N__24021\,
            I => \N__24018\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__24018\,
            I => \N__24014\
        );

    \I__2479\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24011\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__24014\,
            I => \N__24007\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24004\
        );

    \I__2476\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24001\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__24007\,
            I => \N__23996\
        );

    \I__2474\ : Span4Mux_s1_h
    port map (
            O => \N__24004\,
            I => \N__23996\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__24001\,
            I => \N__23993\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__23996\,
            I => \N__23990\
        );

    \I__2471\ : Span4Mux_s2_h
    port map (
            O => \N__23993\,
            I => \N__23987\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__23990\,
            I => \N__23984\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__23987\,
            I => \N__23981\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__23984\,
            I => \pid_alt.error_15\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__23981\,
            I => \pid_alt.error_15\
        );

    \I__2466\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23973\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__23973\,
            I => \N__23970\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__23970\,
            I => \N__23967\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__23967\,
            I => alt_kp_1
        );

    \I__2462\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23961\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__23961\,
            I => drone_altitude_i_10
        );

    \I__2460\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23955\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__23955\,
            I => \N__23952\
        );

    \I__2458\ : Span4Mux_s2_h
    port map (
            O => \N__23952\,
            I => \N__23949\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__23949\,
            I => alt_kp_0
        );

    \I__2456\ : InMux
    port map (
            O => \N__23946\,
            I => \N__23943\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__23943\,
            I => \N__23940\
        );

    \I__2454\ : Span4Mux_s2_h
    port map (
            O => \N__23940\,
            I => \N__23937\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__23937\,
            I => alt_kp_6
        );

    \I__2452\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23930\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__23933\,
            I => \N__23927\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23924\
        );

    \I__2449\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23921\
        );

    \I__2448\ : Odrv12
    port map (
            O => \N__23924\,
            I => alt_command_0
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__23921\,
            I => alt_command_0
        );

    \I__2446\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23913\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__23913\,
            I => \N__23910\
        );

    \I__2444\ : Span4Mux_h
    port map (
            O => \N__23910\,
            I => \N__23905\
        );

    \I__2443\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23902\
        );

    \I__2442\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23899\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__23905\,
            I => \N__23894\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__23902\,
            I => \N__23894\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__23899\,
            I => \N__23891\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__23894\,
            I => \N__23888\
        );

    \I__2437\ : Span4Mux_s3_h
    port map (
            O => \N__23891\,
            I => \N__23885\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__23888\,
            I => \N__23882\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__23885\,
            I => \N__23879\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__23882\,
            I => \pid_alt.error_4\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__23879\,
            I => \pid_alt.error_4\
        );

    \I__2432\ : InMux
    port map (
            O => \N__23874\,
            I => \pid_alt.error_cry_3\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__23871\,
            I => \N__23867\
        );

    \I__2430\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23864\
        );

    \I__2429\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23861\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__23864\,
            I => alt_command_1
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__23861\,
            I => alt_command_1
        );

    \I__2426\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23853\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__23853\,
            I => \N__23850\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__23850\,
            I => \N__23845\
        );

    \I__2423\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23842\
        );

    \I__2422\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23839\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__23845\,
            I => \N__23834\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__23842\,
            I => \N__23834\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23831\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__23834\,
            I => \N__23828\
        );

    \I__2417\ : Span4Mux_s2_h
    port map (
            O => \N__23831\,
            I => \N__23825\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__23828\,
            I => \N__23822\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__23825\,
            I => \N__23819\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__23822\,
            I => \pid_alt.error_5\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__23819\,
            I => \pid_alt.error_5\
        );

    \I__2412\ : InMux
    port map (
            O => \N__23814\,
            I => \pid_alt.error_cry_4\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__23811\,
            I => \N__23807\
        );

    \I__2410\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23804\
        );

    \I__2409\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23801\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__23804\,
            I => alt_command_2
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__23801\,
            I => alt_command_2
        );

    \I__2406\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23791\
        );

    \I__2405\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23788\
        );

    \I__2404\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23785\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__23791\,
            I => \N__23782\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__23788\,
            I => \N__23779\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__23785\,
            I => \N__23776\
        );

    \I__2400\ : Span12Mux_s4_h
    port map (
            O => \N__23782\,
            I => \N__23773\
        );

    \I__2399\ : Span4Mux_s2_h
    port map (
            O => \N__23779\,
            I => \N__23770\
        );

    \I__2398\ : Span4Mux_s2_h
    port map (
            O => \N__23776\,
            I => \N__23767\
        );

    \I__2397\ : Span12Mux_v
    port map (
            O => \N__23773\,
            I => \N__23764\
        );

    \I__2396\ : Span4Mux_v
    port map (
            O => \N__23770\,
            I => \N__23761\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__23767\,
            I => \N__23758\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__23764\,
            I => \pid_alt.error_6\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__23761\,
            I => \pid_alt.error_6\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__23758\,
            I => \pid_alt.error_6\
        );

    \I__2391\ : InMux
    port map (
            O => \N__23751\,
            I => \pid_alt.error_cry_5\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__23748\,
            I => \N__23744\
        );

    \I__2389\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23741\
        );

    \I__2388\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23738\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__23741\,
            I => alt_command_3
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__23738\,
            I => alt_command_3
        );

    \I__2385\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23728\
        );

    \I__2384\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23725\
        );

    \I__2383\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23722\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__23728\,
            I => \N__23719\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__23725\,
            I => \N__23716\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__23722\,
            I => \N__23713\
        );

    \I__2379\ : Span12Mux_s3_h
    port map (
            O => \N__23719\,
            I => \N__23710\
        );

    \I__2378\ : Span4Mux_s2_h
    port map (
            O => \N__23716\,
            I => \N__23707\
        );

    \I__2377\ : Span4Mux_s2_h
    port map (
            O => \N__23713\,
            I => \N__23704\
        );

    \I__2376\ : Span12Mux_v
    port map (
            O => \N__23710\,
            I => \N__23701\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__23707\,
            I => \N__23698\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__23704\,
            I => \N__23695\
        );

    \I__2373\ : Odrv12
    port map (
            O => \N__23701\,
            I => \pid_alt.error_7\
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__23698\,
            I => \pid_alt.error_7\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__23695\,
            I => \pid_alt.error_7\
        );

    \I__2370\ : InMux
    port map (
            O => \N__23688\,
            I => \pid_alt.error_cry_6\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__2368\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__23679\,
            I => alt_command_4
        );

    \I__2366\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__23670\,
            I => \N__23665\
        );

    \I__2363\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23662\
        );

    \I__2362\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23659\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__23665\,
            I => \N__23656\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__23662\,
            I => \N__23653\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__23659\,
            I => \N__23650\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__23656\,
            I => \N__23647\
        );

    \I__2357\ : Span4Mux_s2_h
    port map (
            O => \N__23653\,
            I => \N__23644\
        );

    \I__2356\ : Span4Mux_s3_h
    port map (
            O => \N__23650\,
            I => \N__23641\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__23647\,
            I => \N__23638\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__23644\,
            I => \N__23635\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__23641\,
            I => \N__23632\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__23638\,
            I => \pid_alt.error_8\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__23635\,
            I => \pid_alt.error_8\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__23632\,
            I => \pid_alt.error_8\
        );

    \I__2349\ : InMux
    port map (
            O => \N__23625\,
            I => \bfn_2_20_0_\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__23622\,
            I => \N__23619\
        );

    \I__2347\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23616\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__23613\,
            I => alt_command_5
        );

    \I__2344\ : InMux
    port map (
            O => \N__23610\,
            I => \N__23607\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__23607\,
            I => \N__23602\
        );

    \I__2342\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23599\
        );

    \I__2341\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23596\
        );

    \I__2340\ : Span4Mux_v
    port map (
            O => \N__23602\,
            I => \N__23593\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__23599\,
            I => \N__23590\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__23596\,
            I => \N__23587\
        );

    \I__2337\ : Sp12to4
    port map (
            O => \N__23593\,
            I => \N__23584\
        );

    \I__2336\ : Span4Mux_s2_h
    port map (
            O => \N__23590\,
            I => \N__23581\
        );

    \I__2335\ : Span4Mux_s2_h
    port map (
            O => \N__23587\,
            I => \N__23578\
        );

    \I__2334\ : Span12Mux_s2_h
    port map (
            O => \N__23584\,
            I => \N__23575\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__23581\,
            I => \N__23572\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__23578\,
            I => \N__23569\
        );

    \I__2331\ : Odrv12
    port map (
            O => \N__23575\,
            I => \pid_alt.error_9\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__23572\,
            I => \pid_alt.error_9\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__23569\,
            I => \pid_alt.error_9\
        );

    \I__2328\ : InMux
    port map (
            O => \N__23562\,
            I => \pid_alt.error_cry_8\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__23559\,
            I => \N__23556\
        );

    \I__2326\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23553\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__23553\,
            I => alt_command_6
        );

    \I__2324\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23547\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__2322\ : Span4Mux_s2_h
    port map (
            O => \N__23544\,
            I => \N__23539\
        );

    \I__2321\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23536\
        );

    \I__2320\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23533\
        );

    \I__2319\ : Span4Mux_v
    port map (
            O => \N__23539\,
            I => \N__23530\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__23536\,
            I => \N__23527\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__23533\,
            I => \N__23524\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__23530\,
            I => \N__23521\
        );

    \I__2315\ : Span4Mux_s2_h
    port map (
            O => \N__23527\,
            I => \N__23518\
        );

    \I__2314\ : Span4Mux_s3_h
    port map (
            O => \N__23524\,
            I => \N__23515\
        );

    \I__2313\ : Span4Mux_v
    port map (
            O => \N__23521\,
            I => \N__23512\
        );

    \I__2312\ : Span4Mux_v
    port map (
            O => \N__23518\,
            I => \N__23509\
        );

    \I__2311\ : Span4Mux_v
    port map (
            O => \N__23515\,
            I => \N__23506\
        );

    \I__2310\ : Odrv4
    port map (
            O => \N__23512\,
            I => \pid_alt.error_10\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__23509\,
            I => \pid_alt.error_10\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__23506\,
            I => \pid_alt.error_10\
        );

    \I__2307\ : InMux
    port map (
            O => \N__23499\,
            I => \pid_alt.error_cry_9\
        );

    \I__2306\ : CascadeMux
    port map (
            O => \N__23496\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\
        );

    \I__2305\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23487\
        );

    \I__2304\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23487\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__23487\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\
        );

    \I__2302\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23478\
        );

    \I__2301\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23478\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__23478\,
            I => \N__23475\
        );

    \I__2299\ : Span4Mux_h
    port map (
            O => \N__23475\,
            I => \N__23472\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__23472\,
            I => \pid_alt.error_p_regZ0Z_18\
        );

    \I__2297\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23463\
        );

    \I__2296\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23463\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__23463\,
            I => \pid_alt.error_d_reg_prevZ0Z_18\
        );

    \I__2294\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23451\
        );

    \I__2293\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23451\
        );

    \I__2292\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23451\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__23451\,
            I => \N__23448\
        );

    \I__2290\ : Span12Mux_s8_h
    port map (
            O => \N__23448\,
            I => \N__23445\
        );

    \I__2289\ : Span12Mux_v
    port map (
            O => \N__23445\,
            I => \N__23442\
        );

    \I__2288\ : Odrv12
    port map (
            O => \N__23442\,
            I => \pid_alt.error_d_regZ0Z_18\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__23439\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\
        );

    \I__2286\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23433\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__2284\ : Span4Mux_s1_h
    port map (
            O => \N__23430\,
            I => \N__23426\
        );

    \I__2283\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23423\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__23426\,
            I => \N__23417\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__23423\,
            I => \N__23417\
        );

    \I__2280\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23414\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__23417\,
            I => \N__23411\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23408\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__23411\,
            I => \N__23403\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__23408\,
            I => \N__23403\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__2274\ : Odrv4
    port map (
            O => \N__23400\,
            I => \pid_alt.error_1\
        );

    \I__2273\ : InMux
    port map (
            O => \N__23397\,
            I => \pid_alt.error_cry_0\
        );

    \I__2272\ : InMux
    port map (
            O => \N__23394\,
            I => \N__23391\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__2270\ : Span4Mux_s1_h
    port map (
            O => \N__23388\,
            I => \N__23383\
        );

    \I__2269\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23380\
        );

    \I__2268\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23377\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__23383\,
            I => \N__23372\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__23380\,
            I => \N__23372\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__23377\,
            I => \N__23369\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__23372\,
            I => \N__23366\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__23369\,
            I => \N__23363\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__23366\,
            I => \N__23358\
        );

    \I__2261\ : Span4Mux_v
    port map (
            O => \N__23363\,
            I => \N__23358\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__23358\,
            I => \pid_alt.error_2\
        );

    \I__2259\ : InMux
    port map (
            O => \N__23355\,
            I => \pid_alt.error_cry_1\
        );

    \I__2258\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23349\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23346\
        );

    \I__2256\ : Span4Mux_s1_h
    port map (
            O => \N__23346\,
            I => \N__23342\
        );

    \I__2255\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23339\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__23342\,
            I => \N__23333\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23333\
        );

    \I__2252\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23330\
        );

    \I__2251\ : Span4Mux_v
    port map (
            O => \N__23333\,
            I => \N__23327\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23324\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__23327\,
            I => \N__23321\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__23324\,
            I => \N__23318\
        );

    \I__2247\ : Span4Mux_s1_h
    port map (
            O => \N__23321\,
            I => \N__23313\
        );

    \I__2246\ : Span4Mux_v
    port map (
            O => \N__23318\,
            I => \N__23313\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__23313\,
            I => \pid_alt.error_3\
        );

    \I__2244\ : InMux
    port map (
            O => \N__23310\,
            I => \pid_alt.error_cry_2\
        );

    \I__2243\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__23304\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__23301\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\
        );

    \I__2240\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23292\
        );

    \I__2239\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23292\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__23292\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\
        );

    \I__2237\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23280\
        );

    \I__2236\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23280\
        );

    \I__2235\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23280\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__23280\,
            I => \N__23277\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__2232\ : Sp12to4
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__2231\ : Odrv12
    port map (
            O => \N__23271\,
            I => \pid_alt.error_d_regZ0Z_12\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__23268\,
            I => \N__23265\
        );

    \I__2229\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23259\
        );

    \I__2228\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23259\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__23259\,
            I => \pid_alt.error_d_reg_prevZ0Z_12\
        );

    \I__2226\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23250\
        );

    \I__2225\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23250\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23247\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__23247\,
            I => \N__23244\
        );

    \I__2222\ : Span4Mux_v
    port map (
            O => \N__23244\,
            I => \N__23241\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__23241\,
            I => \pid_alt.error_p_regZ0Z_12\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__23238\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\
        );

    \I__2219\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23232\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__23232\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\
        );

    \I__2217\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23225\
        );

    \I__2216\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23220\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__23225\,
            I => \N__23217\
        );

    \I__2214\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23212\
        );

    \I__2213\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23212\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__23220\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__23217\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__23212\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__23205\,
            I => \N__23202\
        );

    \I__2208\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__23199\,
            I => \pid_alt.N_1666_i\
        );

    \I__2206\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23186\
        );

    \I__2205\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23186\
        );

    \I__2204\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23181\
        );

    \I__2203\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23181\
        );

    \I__2202\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23176\
        );

    \I__2201\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23176\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__23186\,
            I => \N__23173\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__23181\,
            I => \N__23166\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23166\
        );

    \I__2197\ : Span4Mux_s2_h
    port map (
            O => \N__23173\,
            I => \N__23166\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__23166\,
            I => \pid_alt.error_p_regZ0Z_1\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__23163\,
            I => \N__23157\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__23162\,
            I => \N__23153\
        );

    \I__2193\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23147\
        );

    \I__2192\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23147\
        );

    \I__2191\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23142\
        );

    \I__2190\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23142\
        );

    \I__2189\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23137\
        );

    \I__2188\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23137\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__23147\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__23142\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__23137\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__23130\,
            I => \pid_alt.N_1666_i_cascade_\
        );

    \I__2183\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23121\
        );

    \I__2182\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23121\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__23121\,
            I => \N__23115\
        );

    \I__2180\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23108\
        );

    \I__2179\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23108\
        );

    \I__2178\ : InMux
    port map (
            O => \N__23118\,
            I => \N__23108\
        );

    \I__2177\ : Span4Mux_v
    port map (
            O => \N__23115\,
            I => \N__23103\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__23108\,
            I => \N__23100\
        );

    \I__2175\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23095\
        );

    \I__2174\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23095\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__23103\,
            I => \N__23092\
        );

    \I__2172\ : Span12Mux_v
    port map (
            O => \N__23100\,
            I => \N__23087\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__23095\,
            I => \N__23087\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__23092\,
            I => \pid_alt.error_d_regZ0Z_1\
        );

    \I__2169\ : Odrv12
    port map (
            O => \N__23087\,
            I => \pid_alt.error_d_regZ0Z_1\
        );

    \I__2168\ : InMux
    port map (
            O => \N__23082\,
            I => \N__23079\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__23079\,
            I => \pid_alt.un1_pid_prereg_0_axb_2_1\
        );

    \I__2166\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23073\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__23073\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__23070\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_\
        );

    \I__2163\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23064\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__23060\
        );

    \I__2161\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23057\
        );

    \I__2160\ : Span4Mux_v
    port map (
            O => \N__23060\,
            I => \N__23054\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23051\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__23054\,
            I => \N__23046\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__23051\,
            I => \N__23046\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__23046\,
            I => \pid_alt.error_p_regZ0Z_11\
        );

    \I__2155\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23037\
        );

    \I__2154\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23037\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__23037\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11\
        );

    \I__2152\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23027\
        );

    \I__2151\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23027\
        );

    \I__2150\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23024\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__23027\,
            I => \N__23021\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__23024\,
            I => \N__23016\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__23021\,
            I => \N__23016\
        );

    \I__2146\ : Span4Mux_v
    port map (
            O => \N__23016\,
            I => \N__23013\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__23013\,
            I => \pid_alt.error_d_regZ0Z_11\
        );

    \I__2144\ : InMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__23007\,
            I => \N__23004\
        );

    \I__2142\ : Span4Mux_s3_h
    port map (
            O => \N__23004\,
            I => \N__23000\
        );

    \I__2141\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22997\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__23000\,
            I => \pid_alt.error_d_reg_prevZ0Z_11\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__22997\,
            I => \pid_alt.error_d_reg_prevZ0Z_11\
        );

    \I__2138\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22986\
        );

    \I__2137\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22986\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__22986\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\
        );

    \I__2135\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22977\
        );

    \I__2134\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22977\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__22977\,
            I => \pid_alt.error_d_reg_prevZ0Z_5\
        );

    \I__2132\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22965\
        );

    \I__2131\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22965\
        );

    \I__2130\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22965\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22962\
        );

    \I__2128\ : Span12Mux_v
    port map (
            O => \N__22962\,
            I => \N__22959\
        );

    \I__2127\ : Odrv12
    port map (
            O => \N__22959\,
            I => \pid_alt.error_d_regZ0Z_5\
        );

    \I__2126\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22950\
        );

    \I__2125\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22950\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__2123\ : Odrv12
    port map (
            O => \N__22947\,
            I => \pid_alt.error_d_reg_prevZ0Z_6\
        );

    \I__2122\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22937\
        );

    \I__2121\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22937\
        );

    \I__2120\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22934\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__22937\,
            I => \N__22931\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22926\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__22931\,
            I => \N__22926\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__22926\,
            I => \N__22923\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__22923\,
            I => \pid_alt.error_d_regZ0Z_6\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__22920\,
            I => \N__22914\
        );

    \I__2113\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22908\
        );

    \I__2112\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22908\
        );

    \I__2111\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22903\
        );

    \I__2110\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22903\
        );

    \I__2109\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22900\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__22908\,
            I => \N__22897\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__22903\,
            I => \N__22894\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__22900\,
            I => \N__22889\
        );

    \I__2105\ : Span4Mux_s2_h
    port map (
            O => \N__22897\,
            I => \N__22889\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__22894\,
            I => \pid_alt.error_p_regZ0Z_2\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__22889\,
            I => \pid_alt.error_p_regZ0Z_2\
        );

    \I__2102\ : InMux
    port map (
            O => \N__22884\,
            I => \N__22880\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__22883\,
            I => \N__22875\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__22880\,
            I => \N__22871\
        );

    \I__2099\ : InMux
    port map (
            O => \N__22879\,
            I => \N__22866\
        );

    \I__2098\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22866\
        );

    \I__2097\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22861\
        );

    \I__2096\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22861\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__22871\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__22866\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__22861\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__2092\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__22851\,
            I => \N__22848\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__22848\,
            I => \N__22840\
        );

    \I__2089\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22835\
        );

    \I__2088\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22835\
        );

    \I__2087\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22828\
        );

    \I__2086\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22828\
        );

    \I__2085\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22828\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__22840\,
            I => \N__22825\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__22835\,
            I => \N__22820\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__22828\,
            I => \N__22820\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__22825\,
            I => \pid_alt.error_d_regZ0Z_2\
        );

    \I__2080\ : Odrv12
    port map (
            O => \N__22820\,
            I => \pid_alt.error_d_regZ0Z_2\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__22815\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_\
        );

    \I__2078\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22809\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__22809\,
            I => \N__22806\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__22803\,
            I => \N__22800\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__22800\,
            I => \pid_alt.O_5_4\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__22797\,
            I => \N__22794\
        );

    \I__2072\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22788\
        );

    \I__2071\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22788\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__22788\,
            I => \Commands_frame_decoder.stateZ0Z_3\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__22785\,
            I => \N__22780\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__22784\,
            I => \N__22777\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__22783\,
            I => \N__22774\
        );

    \I__2066\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22764\
        );

    \I__2065\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22764\
        );

    \I__2064\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22764\
        );

    \I__2063\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22764\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__2061\ : Span4Mux_s3_h
    port map (
            O => \N__22761\,
            I => \N__22758\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__22758\,
            I => \N__22754\
        );

    \I__2059\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22751\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__22754\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__22751\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__22746\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\
        );

    \I__2055\ : CEMux
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__22740\,
            I => \N__22737\
        );

    \I__2053\ : Span4Mux_v
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__22734\,
            I => \N__22731\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__22731\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\
        );

    \I__2050\ : InMux
    port map (
            O => \N__22728\,
            I => \N__22725\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__22725\,
            I => \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\
        );

    \I__2048\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22719\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__2046\ : Span4Mux_h
    port map (
            O => \N__22716\,
            I => \N__22713\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__22713\,
            I => \pid_alt.O_4_5\
        );

    \I__2044\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22707\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__22704\,
            I => \N__22701\
        );

    \I__2041\ : Span4Mux_v
    port map (
            O => \N__22701\,
            I => \N__22698\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__22698\,
            I => \pid_alt.O_3_4\
        );

    \I__2039\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22692\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__22692\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__22689\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_\
        );

    \I__2036\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22683\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__22680\,
            I => alt_kd_6
        );

    \I__2033\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22674\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22671\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__22671\,
            I => alt_kd_4
        );

    \I__2030\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22665\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__22665\,
            I => \N__22662\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__22662\,
            I => \N__22659\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__22659\,
            I => alt_kd_3
        );

    \I__2026\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22650\
        );

    \I__2024\ : Span4Mux_s2_h
    port map (
            O => \N__22650\,
            I => \N__22647\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__22647\,
            I => alt_kd_0
        );

    \I__2022\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22641\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__2020\ : Span4Mux_s3_h
    port map (
            O => \N__22638\,
            I => \N__22635\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__22635\,
            I => alt_ki_0
        );

    \I__2018\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22629\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__22629\,
            I => \N__22626\
        );

    \I__2016\ : Span4Mux_v
    port map (
            O => \N__22626\,
            I => \N__22623\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__22623\,
            I => alt_ki_2
        );

    \I__2014\ : CEMux
    port map (
            O => \N__22620\,
            I => \N__22617\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22612\
        );

    \I__2012\ : CEMux
    port map (
            O => \N__22616\,
            I => \N__22609\
        );

    \I__2011\ : CEMux
    port map (
            O => \N__22615\,
            I => \N__22606\
        );

    \I__2010\ : Span4Mux_s3_h
    port map (
            O => \N__22612\,
            I => \N__22603\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__22609\,
            I => \N__22598\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__22606\,
            I => \N__22598\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__22603\,
            I => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__22598\,
            I => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\
        );

    \I__2005\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22587\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__22584\,
            I => \pid_alt.g0_4_0\
        );

    \I__2001\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__22578\,
            I => \N__22575\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__22575\,
            I => \pid_alt.O_5_18\
        );

    \I__1998\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22569\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__22569\,
            I => \N__22566\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__22566\,
            I => \pid_alt.O_5_21\
        );

    \I__1995\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22560\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__22560\,
            I => \N__22557\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__22557\,
            I => \pid_alt.O_5_19\
        );

    \I__1992\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22551\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__22551\,
            I => \pid_alt.O_5_14\
        );

    \I__1990\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22545\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__22542\,
            I => \pid_alt.O_5_23\
        );

    \I__1987\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22536\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__22536\,
            I => \N__22533\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__22533\,
            I => \pid_alt.O_5_16\
        );

    \I__1984\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22527\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__22527\,
            I => \pid_alt.O_5_12\
        );

    \I__1982\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22521\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__22521\,
            I => \pid_alt.O_5_13\
        );

    \I__1980\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22515\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__22515\,
            I => \N__22512\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__22512\,
            I => \pid_alt.O_5_24\
        );

    \I__1977\ : InMux
    port map (
            O => \N__22509\,
            I => \N__22506\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__22506\,
            I => \N__22503\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__22503\,
            I => \pid_alt.O_5_7\
        );

    \I__1974\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22497\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__22497\,
            I => \N__22494\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__22494\,
            I => \pid_alt.O_5_8\
        );

    \I__1971\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22488\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__22488\,
            I => \N__22485\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__22485\,
            I => \N__22482\
        );

    \I__1968\ : Span4Mux_v
    port map (
            O => \N__22482\,
            I => \N__22479\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__22479\,
            I => \N__22476\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__22476\,
            I => \pid_alt.O_4_8\
        );

    \I__1965\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__22470\,
            I => \N__22467\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__22467\,
            I => \pid_alt.O_5_11\
        );

    \I__1962\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__1960\ : Span4Mux_h
    port map (
            O => \N__22458\,
            I => \N__22455\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__22455\,
            I => \pid_alt.O_5_22\
        );

    \I__1958\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__22449\,
            I => \N__22446\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__22446\,
            I => \pid_alt.O_5_15\
        );

    \I__1955\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22440\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__22440\,
            I => \N__22437\
        );

    \I__1953\ : Odrv4
    port map (
            O => \N__22437\,
            I => \pid_alt.O_5_17\
        );

    \I__1952\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22431\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__22428\,
            I => \pid_alt.O_5_20\
        );

    \I__1949\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22422\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__1947\ : Span4Mux_h
    port map (
            O => \N__22419\,
            I => \N__22416\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__22416\,
            I => \N__22413\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__22413\,
            I => \pid_alt.O_5_5\
        );

    \I__1944\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22407\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__22407\,
            I => \N__22404\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__22404\,
            I => \pid_front.O_0_8\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__22401\,
            I => \Commands_frame_decoder.source_CH1data8_cascade_\
        );

    \I__1940\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22389\
        );

    \I__1939\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22389\
        );

    \I__1938\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22389\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__22389\,
            I => \Commands_frame_decoder.source_CH1data8\
        );

    \I__1936\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22383\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22380\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__22380\,
            I => \pid_front.O_0_22\
        );

    \I__1933\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22374\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__22374\,
            I => \N__22371\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__22371\,
            I => \pid_front.O_0_23\
        );

    \I__1930\ : InMux
    port map (
            O => \N__22368\,
            I => \N__22365\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__22365\,
            I => \N__22362\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__22362\,
            I => \pid_front.O_0_24\
        );

    \I__1927\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__22356\,
            I => \pid_front.O_0_21\
        );

    \I__1925\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22350\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__22350\,
            I => \pid_front.O_0_20\
        );

    \I__1923\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22344\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__22344\,
            I => \pid_front.O_0_14\
        );

    \I__1921\ : InMux
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__22338\,
            I => \pid_front.O_0_10\
        );

    \I__1919\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__22332\,
            I => \pid_front.O_0_13\
        );

    \I__1917\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__22323\,
            I => \N__22320\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__22320\,
            I => \N__22317\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__22317\,
            I => \pid_alt.O_5_6\
        );

    \I__1912\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__22311\,
            I => \pid_alt.N_5\
        );

    \I__1910\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__22305\,
            I => \pid_alt.N_1672_0\
        );

    \I__1908\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22299\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__22299\,
            I => \N__22296\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__22296\,
            I => \pid_front.O_0_16\
        );

    \I__1905\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__22290\,
            I => \N__22287\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__22287\,
            I => \pid_front.O_0_17\
        );

    \I__1902\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22281\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__22281\,
            I => \N__22278\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__22278\,
            I => \pid_front.O_0_18\
        );

    \I__1899\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22272\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__22272\,
            I => \N__22269\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__22269\,
            I => \pid_front.O_0_19\
        );

    \I__1896\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22263\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__22263\,
            I => \pid_front.O_0_12\
        );

    \I__1894\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22257\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__22257\,
            I => \pid_front.O_0_7\
        );

    \I__1892\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22251\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__22251\,
            I => \pid_alt.N_3_1\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__22248\,
            I => \N__22245\
        );

    \I__1889\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__22242\,
            I => \pid_alt.N_1668_1\
        );

    \I__1887\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__22236\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2\
        );

    \I__1885\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22230\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__22230\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__22227\,
            I => \pid_alt.N_1674_0_cascade_\
        );

    \I__1882\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22221\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__22221\,
            I => \pid_alt.N_1666_i_0\
        );

    \I__1880\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22215\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__22215\,
            I => \pid_alt.N_3_0\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__1877\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22206\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__22206\,
            I => \pid_alt.N_1668_0\
        );

    \I__1875\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22200\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__22200\,
            I => \pid_alt.O_4_19\
        );

    \I__1873\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22194\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__22194\,
            I => \pid_alt.O_4_6\
        );

    \I__1871\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22188\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__22188\,
            I => \pid_alt.O_4_21\
        );

    \I__1869\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22182\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__22182\,
            I => \pid_alt.O_4_13\
        );

    \I__1867\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22176\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__22176\,
            I => \pid_alt.O_4_12\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__22173\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_\
        );

    \I__1864\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22167\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__22167\,
            I => \pid_alt.N_1666_i_1\
        );

    \I__1862\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22161\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__22161\,
            I => \N__22158\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__22158\,
            I => \pid_alt.O_4_23\
        );

    \I__1859\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22152\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__22149\,
            I => \pid_alt.O_4_22\
        );

    \I__1856\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22143\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__22143\,
            I => \pid_alt.O_4_10\
        );

    \I__1854\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__22137\,
            I => \pid_alt.O_4_14\
        );

    \I__1852\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22131\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__22131\,
            I => \pid_alt.O_4_11\
        );

    \I__1850\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__22122\,
            I => \pid_alt.O_4_17\
        );

    \I__1847\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__22116\,
            I => \pid_alt.O_4_16\
        );

    \I__1845\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22110\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__22110\,
            I => \pid_alt.O_4_20\
        );

    \I__1843\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22104\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__22104\,
            I => \pid_alt.O_4_18\
        );

    \I__1841\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22098\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__22098\,
            I => alt_kd_5
        );

    \I__1839\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22092\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__1837\ : Span4Mux_s2_h
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__22086\,
            I => alt_ki_6
        );

    \I__1835\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__22080\,
            I => \N__22077\
        );

    \I__1833\ : Span4Mux_s2_h
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__22074\,
            I => alt_ki_7
        );

    \I__1831\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22068\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__22068\,
            I => \N__22065\
        );

    \I__1829\ : Span4Mux_s2_h
    port map (
            O => \N__22065\,
            I => \N__22062\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__22062\,
            I => alt_ki_1
        );

    \I__1827\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22056\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__22056\,
            I => \N__22053\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__22053\,
            I => alt_ki_3
        );

    \I__1824\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22047\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__22047\,
            I => \N__22044\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__22044\,
            I => alt_ki_4
        );

    \I__1821\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22038\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__22035\
        );

    \I__1819\ : Span4Mux_s2_h
    port map (
            O => \N__22035\,
            I => \N__22032\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__22032\,
            I => alt_ki_5
        );

    \I__1817\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22026\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__22026\,
            I => \pid_alt.O_4_9\
        );

    \I__1815\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22020\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__22020\,
            I => \N__22017\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__22017\,
            I => \pid_alt.O_4_24\
        );

    \I__1812\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22011\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__22011\,
            I => \pid_alt.O_3_21\
        );

    \I__1810\ : InMux
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__22005\,
            I => \pid_alt.O_3_22\
        );

    \I__1808\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21999\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__21999\,
            I => \pid_alt.O_3_23\
        );

    \I__1806\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21993\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__21993\,
            I => \pid_alt.O_3_6\
        );

    \I__1804\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21984\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__21984\,
            I => \pid_alt.O_3_24\
        );

    \I__1801\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__21978\,
            I => \pid_alt.O_3_7\
        );

    \I__1799\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__21972\,
            I => \pid_alt.O_3_9\
        );

    \I__1797\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21966\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__21966\,
            I => alt_kd_7
        );

    \I__1795\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__21960\,
            I => alt_kd_2
        );

    \I__1793\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21954\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__21954\,
            I => alt_kd_1
        );

    \I__1791\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21945\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__21945\,
            I => \pid_alt.O_3_10\
        );

    \I__1788\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21939\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__21939\,
            I => \pid_alt.O_3_5\
        );

    \I__1786\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21933\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__21933\,
            I => \pid_alt.O_3_14\
        );

    \I__1784\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__21927\,
            I => \pid_alt.O_3_15\
        );

    \I__1782\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21921\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__21921\,
            I => \N__21918\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__21918\,
            I => \pid_alt.O_3_16\
        );

    \I__1779\ : InMux
    port map (
            O => \N__21915\,
            I => \N__21912\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__21912\,
            I => \N__21909\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__21909\,
            I => \pid_alt.O_3_17\
        );

    \I__1776\ : InMux
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__21900\,
            I => \pid_alt.O_3_18\
        );

    \I__1773\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__21894\,
            I => \N__21891\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__21891\,
            I => \pid_alt.O_3_19\
        );

    \I__1770\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21885\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__21885\,
            I => \N__21882\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__21882\,
            I => \pid_alt.O_3_20\
        );

    \I__1767\ : IoInMux
    port map (
            O => \N__21879\,
            I => \N__21876\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__1765\ : IoSpan4Mux
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__1764\ : Span4Mux_s2_v
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__1763\ : Sp12to4
    port map (
            O => \N__21867\,
            I => \N__21864\
        );

    \I__1762\ : Span12Mux_v
    port map (
            O => \N__21864\,
            I => \N__21861\
        );

    \I__1761\ : Span12Mux_v
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__1760\ : Odrv12
    port map (
            O => \N__21858\,
            I => \Pc2drone_pll_inst.clk_system_pll\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_6\,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_14\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_22\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un3_source_data_0_cry_7\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un2_source_data_0_cry_8\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_throttle_cry_7\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_rudder_cry_13\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_elevator_cry_7\,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_aileron_cry_7\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.counter24_0_data_tmp_7\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_2_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.error_cry_7\,
            carryinitout => \bfn_2_20_0_\
        );

    \IN_MUX_bfv_20_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_9_0_\
        );

    \IN_MUX_bfv_20_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_side.un1_pid_prereg_cry_5\,
            carryinitout => \bfn_20_10_0_\
        );

    \IN_MUX_bfv_20_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_side.un1_pid_prereg_cry_13\,
            carryinitout => \bfn_20_11_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_front.un1_pid_prereg_cry_5\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_12_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_front.un1_pid_prereg_cry_13\,
            carryinitout => \bfn_12_23_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_7\,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_15\,
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_21_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_17_0_\
        );

    \IN_MUX_bfv_21_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_side.error_cry_3_0\,
            carryinitout => \bfn_21_18_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_front.error_cry_3_0\,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \dron_frame_decoder_1.un1_WDT_cry_7\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Commands_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_8_6_0_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__41964\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_419_g\
        );

    \pid_alt.state_RNICP2N1_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__47781\,
            GLOBALBUFFEROUTPUT => \pid_alt.N_664_0_g\
        );

    \Pc2drone_pll_inst.PLLOUTCORE_derived_clock_RNI5FOA\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21879\,
            GLOBALBUFFEROUTPUT => clk_system_pll_g
        );

    \reset_module_System.reset_RNITC69_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__49272\,
            GLOBALBUFFEROUTPUT => \N_665_g\
        );

    \reset_module_System.reset_RNITC69\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__44971\,
            GLOBALBUFFEROUTPUT => reset_system_g
        );

    \pid_front.state_RNIPKTD_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__31203\,
            GLOBALBUFFEROUTPUT => \pid_front.state_0_g_0\
        );

    \pid_side.state_RNIL5IF_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__35586\,
            GLOBALBUFFEROUTPUT => \pid_side.state_0_g_0\
        );

    \pid_alt.state_RNIH1EN_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__39351\,
            GLOBALBUFFEROUTPUT => \pid_alt.state_0_g_0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_6_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21951\,
            lcout => \pid_alt.error_d_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59139\,
            ce => \N__24449\,
            sr => \N__58219\
        );

    \pid_alt.error_d_reg_esr_1_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21942\,
            lcout => \pid_alt.error_d_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_10_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21936\,
            lcout => \pid_alt.error_d_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_11_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21930\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_12_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_13_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21915\,
            lcout => \pid_alt.error_d_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_14_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21906\,
            lcout => \pid_alt.error_d_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_15_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21897\,
            lcout => \pid_alt.error_d_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_16_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21888\,
            lcout => \pid_alt.error_d_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59152\,
            ce => \N__24450\,
            sr => \N__58218\
        );

    \pid_alt.error_d_reg_esr_17_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22014\,
            lcout => \pid_alt.error_d_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59165\,
            ce => \N__24451\,
            sr => \N__58217\
        );

    \pid_alt.error_d_reg_esr_18_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22008\,
            lcout => \pid_alt.error_d_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59165\,
            ce => \N__24451\,
            sr => \N__58217\
        );

    \pid_alt.error_d_reg_esr_19_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22002\,
            lcout => \pid_alt.error_d_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59165\,
            ce => \N__24451\,
            sr => \N__58217\
        );

    \pid_alt.error_d_reg_esr_2_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21996\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59165\,
            ce => \N__24451\,
            sr => \N__58217\
        );

    \pid_alt.error_d_reg_esr_20_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21990\,
            lcout => \pid_alt.error_d_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59165\,
            ce => \N__24451\,
            sr => \N__58217\
        );

    \pid_alt.error_d_reg_esr_3_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21981\,
            lcout => \pid_alt.error_d_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59165\,
            ce => \N__24451\,
            sr => \N__58217\
        );

    \pid_alt.error_d_reg_esr_5_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21975\,
            lcout => \pid_alt.error_d_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59165\,
            ce => \N__24451\,
            sr => \N__58217\
        );

    \Commands_frame_decoder.source_alt_kd_7_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55566\,
            lcout => alt_kd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59179\,
            ce => \N__24282\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_2_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56111\,
            lcout => alt_kd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59179\,
            ce => \N__24282\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_1_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56278\,
            in2 => \_gnd_net_\,
            in3 => \N__58354\,
            lcout => alt_kd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59179\,
            ce => \N__24282\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_5_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55899\,
            lcout => alt_kd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59179\,
            ce => \N__24282\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_6_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55732\,
            in2 => \_gnd_net_\,
            in3 => \N__58352\,
            lcout => alt_ki_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59194\,
            ce => \N__22615\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58353\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55565\,
            lcout => alt_ki_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59194\,
            ce => \N__22615\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56242\,
            in2 => \_gnd_net_\,
            in3 => \N__58346\,
            lcout => alt_ki_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59206\,
            ce => \N__22620\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_3_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55354\,
            in2 => \_gnd_net_\,
            in3 => \N__58347\,
            lcout => alt_ki_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59206\,
            ce => \N__22620\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_4_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53360\,
            lcout => alt_ki_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59206\,
            ce => \N__22620\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_5_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55876\,
            in2 => \_gnd_net_\,
            in3 => \N__58349\,
            lcout => alt_ki_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59206\,
            ce => \N__22620\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_5_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22029\,
            lcout => \pid_alt.error_i_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_20_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22023\,
            lcout => \pid_alt.error_i_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_19_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22164\,
            lcout => \pid_alt.error_i_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_18_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22155\,
            lcout => \pid_alt.error_i_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_6_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22146\,
            lcout => \pid_alt.error_i_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_10_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22140\,
            lcout => \pid_alt.error_i_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_7_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22134\,
            lcout => \pid_alt.error_i_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_13_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22128\,
            lcout => \pid_alt.error_i_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59221\,
            ce => \N__24453\,
            sr => \N__58215\
        );

    \pid_alt.error_i_reg_esr_12_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22119\,
            lcout => \pid_alt.error_i_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_i_reg_esr_16_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22113\,
            lcout => \pid_alt.error_i_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_i_reg_esr_14_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22107\,
            lcout => \pid_alt.error_i_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_i_reg_esr_15_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22203\,
            lcout => \pid_alt.error_i_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_i_reg_esr_2_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22197\,
            lcout => \pid_alt.error_i_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_i_reg_esr_17_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22191\,
            lcout => \pid_alt.error_i_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_i_reg_esr_9_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22185\,
            lcout => \pid_alt.error_i_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_i_reg_esr_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22179\,
            lcout => \pid_alt.error_i_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59237\,
            ce => \N__24454\,
            sr => \N__58213\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__23067\,
            in1 => \N__23010\,
            in2 => \_gnd_net_\,
            in3 => \N__23032\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110001"
        )
    port map (
            in0 => \N__22170\,
            in1 => \N__22239\,
            in2 => \N__22248\,
            in3 => \N__22254\,
            lcout => OPEN,
            ltout => \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22728\,
            in1 => \N__25869\,
            in2 => \N__22173\,
            in3 => \N__22233\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23229\,
            in2 => \_gnd_net_\,
            in3 => \N__24389\,
            lcout => \pid_alt.N_1666_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23195\,
            in1 => \N__23152\,
            in2 => \_gnd_net_\,
            in3 => \N__23106\,
            lcout => \pid_alt.N_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__23107\,
            in1 => \_gnd_net_\,
            in2 => \N__23162\,
            in3 => \N__23196\,
            lcout => \pid_alt.N_1668_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22918\,
            in1 => \N__22874\,
            in2 => \_gnd_net_\,
            in3 => \N__22843\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__22844\,
            in1 => \_gnd_net_\,
            in2 => \N__22883\,
            in3 => \N__22919\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_2_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22845\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59270\,
            ce => \N__27612\,
            sr => \N__57531\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110001"
        )
    port map (
            in0 => \N__22224\,
            in1 => \N__22314\,
            in2 => \N__22212\,
            in3 => \N__22218\,
            lcout => OPEN,
            ltout => \pid_alt.N_1674_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011010100"
        )
    port map (
            in0 => \N__22593\,
            in1 => \N__22308\,
            in2 => \N__22227\,
            in3 => \N__24661\,
            lcout => \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23228\,
            in2 => \_gnd_net_\,
            in3 => \N__24390\,
            lcout => \pid_alt.N_1666_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23191\,
            in1 => \N__23156\,
            in2 => \_gnd_net_\,
            in3 => \N__23118\,
            lcout => \pid_alt.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__23119\,
            in1 => \_gnd_net_\,
            in2 => \N__23163\,
            in3 => \N__23192\,
            lcout => \pid_alt.N_1668_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22878\,
            in1 => \_gnd_net_\,
            in2 => \N__22920\,
            in3 => \N__22846\,
            lcout => \pid_alt.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__22847\,
            in1 => \N__22917\,
            in2 => \_gnd_net_\,
            in3 => \N__22879\,
            lcout => \pid_alt.N_1672_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_1_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23120\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59283\,
            ce => \N__27609\,
            sr => \N__57538\
        );

    \pid_front.error_p_reg_esr_12_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22302\,
            lcout => \pid_front.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_13_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22293\,
            lcout => \pid_front.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_14_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_15_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22275\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_8_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22266\,
            lcout => \pid_front.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_3_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22260\,
            lcout => \pid_front.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_18_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22386\,
            lcout => \pid_front.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_19_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22377\,
            lcout => \pid_front.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59293\,
            ce => \N__58537\,
            sr => \N__58211\
        );

    \pid_front.error_p_reg_esr_20_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22368\,
            lcout => \pid_front.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59303\,
            ce => \N__58539\,
            sr => \N__58209\
        );

    \pid_front.error_p_reg_esr_17_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22359\,
            lcout => \pid_front.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59303\,
            ce => \N__58539\,
            sr => \N__58209\
        );

    \pid_front.error_p_reg_esr_16_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22353\,
            lcout => \pid_front.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59303\,
            ce => \N__58539\,
            sr => \N__58209\
        );

    \pid_front.error_p_reg_esr_10_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22347\,
            lcout => \pid_front.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59303\,
            ce => \N__58539\,
            sr => \N__58209\
        );

    \pid_front.error_p_reg_esr_6_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22341\,
            lcout => \pid_front.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59303\,
            ce => \N__58539\,
            sr => \N__58209\
        );

    \pid_front.error_p_reg_esr_9_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22335\,
            lcout => \pid_front.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59303\,
            ce => \N__58539\,
            sr => \N__58209\
        );

    \pid_alt.error_p_reg_esr_2_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22329\,
            lcout => \pid_alt.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59310\,
            ce => \N__24457\,
            sr => \N__58208\
        );

    \pid_alt.error_p_reg_esr_1_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22425\,
            lcout => \pid_alt.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59310\,
            ce => \N__24457\,
            sr => \N__58208\
        );

    \pid_front.error_p_reg_esr_4_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22410\,
            lcout => \pid_front.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59314\,
            ce => \N__58538\,
            sr => \N__58207\
        );

    \Commands_frame_decoder.source_CH1data_3_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__22398\,
            in1 => \N__55373\,
            in2 => \N__22785\,
            in3 => \N__23747\,
            lcout => alt_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59318\,
            ce => 'H',
            sr => \N__57580\
        );

    \Commands_frame_decoder.source_CH1data_1_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__22396\,
            in1 => \N__56304\,
            in2 => \N__22783\,
            in3 => \N__23870\,
            lcout => alt_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59318\,
            ce => 'H',
            sr => \N__57580\
        );

    \Commands_frame_decoder.source_CH1data8lto7_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__29166\,
            in1 => \N__24411\,
            in2 => \N__53405\,
            in3 => \N__55716\,
            lcout => \Commands_frame_decoder.source_CH1data8\,
            ltout => \Commands_frame_decoder.source_CH1data8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_0_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__23934\,
            in1 => \N__56486\,
            in2 => \N__22401\,
            in3 => \N__22773\,
            lcout => alt_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59318\,
            ce => 'H',
            sr => \N__57580\
        );

    \Commands_frame_decoder.source_CH1data_2_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__22397\,
            in1 => \N__56139\,
            in2 => \N__22784\,
            in3 => \N__23810\,
            lcout => alt_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59318\,
            ce => 'H',
            sr => \N__57580\
        );

    \Commands_frame_decoder.source_CH1data_esr_4_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53401\,
            lcout => alt_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59321\,
            ce => \N__22743\,
            sr => \N__57589\
        );

    \Commands_frame_decoder.source_CH1data_esr_5_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55927\,
            lcout => alt_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59321\,
            ce => \N__22743\,
            sr => \N__57589\
        );

    \Commands_frame_decoder.source_CH1data_esr_6_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55750\,
            lcout => alt_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59321\,
            ce => \N__22743\,
            sr => \N__57589\
        );

    \Commands_frame_decoder.source_CH1data_esr_7_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55583\,
            lcout => alt_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59321\,
            ce => \N__22743\,
            sr => \N__57589\
        );

    \pid_alt.error_p_reg_esr_3_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22509\,
            lcout => \pid_alt.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59326\,
            ce => \N__24458\,
            sr => \N__58205\
        );

    \pid_alt.error_p_reg_esr_4_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22500\,
            lcout => \pid_alt.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59326\,
            ce => \N__24458\,
            sr => \N__58205\
        );

    \pid_alt.error_i_reg_esr_4_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22491\,
            lcout => \pid_alt.error_i_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59331\,
            ce => \N__24459\,
            sr => \N__58203\
        );

    \pid_alt.error_p_reg_esr_7_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59331\,
            ce => \N__24459\,
            sr => \N__58203\
        );

    \pid_alt.error_p_reg_esr_18_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22464\,
            lcout => \pid_alt.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59331\,
            ce => \N__24459\,
            sr => \N__58203\
        );

    \pid_alt.error_p_reg_esr_11_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22452\,
            lcout => \pid_alt.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59331\,
            ce => \N__24459\,
            sr => \N__58203\
        );

    \pid_alt.error_p_reg_esr_13_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22443\,
            lcout => \pid_alt.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59331\,
            ce => \N__24459\,
            sr => \N__58203\
        );

    \pid_alt.error_p_reg_esr_16_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22434\,
            lcout => \pid_alt.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59331\,
            ce => \N__24459\,
            sr => \N__58203\
        );

    \pid_alt.error_p_reg_esr_14_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22581\,
            lcout => \pid_alt.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59331\,
            ce => \N__24459\,
            sr => \N__58203\
        );

    \pid_alt.error_p_reg_esr_17_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22572\,
            lcout => \pid_alt.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59334\,
            ce => \N__24461\,
            sr => \N__58201\
        );

    \pid_alt.error_p_reg_esr_15_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22563\,
            lcout => \pid_alt.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59334\,
            ce => \N__24461\,
            sr => \N__58201\
        );

    \pid_alt.error_p_reg_esr_10_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22554\,
            lcout => \pid_alt.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59334\,
            ce => \N__24461\,
            sr => \N__58201\
        );

    \pid_alt.error_p_reg_esr_19_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22548\,
            lcout => \pid_alt.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59334\,
            ce => \N__24461\,
            sr => \N__58201\
        );

    \pid_alt.error_p_reg_esr_12_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22539\,
            lcout => \pid_alt.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59334\,
            ce => \N__24461\,
            sr => \N__58201\
        );

    \pid_alt.error_p_reg_esr_8_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22530\,
            lcout => \pid_alt.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59334\,
            ce => \N__24461\,
            sr => \N__58201\
        );

    \pid_alt.error_p_reg_esr_9_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22524\,
            lcout => \pid_alt.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59334\,
            ce => \N__24461\,
            sr => \N__58201\
        );

    \pid_alt.error_p_reg_esr_20_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22518\,
            lcout => \pid_alt.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59337\,
            ce => \N__24462\,
            sr => \N__58198\
        );

    \Commands_frame_decoder.source_alt_kd_6_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58359\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55731\,
            lcout => alt_kd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59154\,
            ce => \N__24275\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_4_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53386\,
            in2 => \_gnd_net_\,
            in3 => \N__58358\,
            lcout => alt_kd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59154\,
            ce => \N__24275\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_3_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55355\,
            lcout => alt_kd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59169\,
            ce => \N__24271\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_0_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56465\,
            in2 => \_gnd_net_\,
            in3 => \N__58350\,
            lcout => alt_kd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59169\,
            ce => \N__24271\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIQRI31_10_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__29352\,
            in1 => \N__31773\,
            in2 => \_gnd_net_\,
            in3 => \N__57866\,
            lcout => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_6_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22942\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59198\,
            ce => \N__27615\,
            sr => \N__57507\
        );

    \Commands_frame_decoder.source_alt_ki_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56464\,
            in2 => \_gnd_net_\,
            in3 => \N__58344\,
            lcout => alt_ki_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59210\,
            ce => \N__22616\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_2_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56125\,
            in2 => \_gnd_net_\,
            in3 => \N__58345\,
            lcout => alt_ki_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59210\,
            ce => \N__22616\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24627\,
            in2 => \_gnd_net_\,
            in3 => \N__24604\,
            lcout => \pid_alt.g0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_3_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__31741\,
            in1 => \N__22757\,
            in2 => \N__22797\,
            in3 => \N__31317\,
            lcout => \Commands_frame_decoder.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59242\,
            ce => 'H',
            sr => \N__57520\
        );

    \Commands_frame_decoder.state_RNIFJ1J_3_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22793\,
            in2 => \_gnd_net_\,
            in3 => \N__31739\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIEI1J_2_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25668\,
            in2 => \_gnd_net_\,
            in3 => \N__31740\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0\,
            ltout => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIBV7S_2_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22746\,
            in3 => \N__57854\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24662\,
            in1 => \N__24625\,
            in2 => \_gnd_net_\,
            in3 => \N__24600\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_1_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22722\,
            lcout => \pid_alt.error_i_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59259\,
            ce => \N__24455\,
            sr => \N__58212\
        );

    \pid_alt.error_d_reg_esr_0_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22710\,
            lcout => \pid_alt.error_d_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59259\,
            ce => \N__24455\,
            sr => \N__58212\
        );

    \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22695\,
            in1 => \N__22991\,
            in2 => \N__25157\,
            in3 => \N__27835\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24351\,
            in1 => \N__22983\,
            in2 => \_gnd_net_\,
            in3 => \N__22973\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22992\,
            in2 => \N__22689\,
            in3 => \N__27836\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24326\,
            in1 => \N__22955\,
            in2 => \_gnd_net_\,
            in3 => \N__22943\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_5_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59274\,
            ce => \N__27606\,
            sr => \N__57532\
        );

    \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24350\,
            in1 => \N__22982\,
            in2 => \_gnd_net_\,
            in3 => \N__22972\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24327\,
            in1 => \N__22956\,
            in2 => \_gnd_net_\,
            in3 => \N__22944\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__22913\,
            in1 => \N__22884\,
            in2 => \_gnd_net_\,
            in3 => \N__22854\,
            lcout => OPEN,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25727\,
            in2 => \N__22815\,
            in3 => \N__23082\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25319\,
            in1 => \N__23224\,
            in2 => \_gnd_net_\,
            in3 => \N__24393\,
            lcout => \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23194\,
            in1 => \N__23161\,
            in2 => \N__23205\,
            in3 => \N__23127\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_0_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22812\,
            lcout => \pid_alt.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59287\,
            ce => \N__24456\,
            sr => \N__58210\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23223\,
            in2 => \_gnd_net_\,
            in3 => \N__24392\,
            lcout => \pid_alt.N_1666_i\,
            ltout => \pid_alt.N_1666_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001011010100"
        )
    port map (
            in0 => \N__23193\,
            in1 => \N__23160\,
            in2 => \N__23130\,
            in3 => \N__23126\,
            lcout => \pid_alt.un1_pid_prereg_0_axb_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23042\,
            in1 => \N__23076\,
            in2 => \N__25400\,
            in3 => \N__24880\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__26309\,
            in1 => \N__26282\,
            in2 => \_gnd_net_\,
            in3 => \N__26269\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__23043\,
            in1 => \_gnd_net_\,
            in2 => \N__23070\,
            in3 => \N__24881\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__23063\,
            in1 => \N__23003\,
            in2 => \_gnd_net_\,
            in3 => \N__23033\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_10_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26270\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59297\,
            ce => \N__27604\,
            sr => \N__57546\
        );

    \pid_alt.error_d_reg_prev_esr_11_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23034\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59297\,
            ce => \N__27604\,
            sr => \N__57546\
        );

    \pid_alt.error_i_acumm_prereg_esr_11_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59297\,
            ce => \N__27604\,
            sr => \N__57546\
        );

    \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23297\,
            in1 => \N__23307\,
            in2 => \N__25899\,
            in3 => \N__24829\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__23255\,
            in1 => \N__23264\,
            in2 => \_gnd_net_\,
            in3 => \N__23287\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__23298\,
            in1 => \_gnd_net_\,
            in2 => \N__23301\,
            in3 => \N__24830\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__25542\,
            in1 => \N__25598\,
            in2 => \_gnd_net_\,
            in3 => \N__25565\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_12_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23289\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59305\,
            ce => \N__27602\,
            sr => \N__57556\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__23288\,
            in1 => \_gnd_net_\,
            in2 => \N__23268\,
            in3 => \N__23256\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__25922\,
            in1 => \N__25946\,
            in2 => \N__23238\,
            in3 => \N__25367\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23235\,
            in1 => \N__23492\,
            in2 => \N__25458\,
            in3 => \N__25060\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__23484\,
            in1 => \N__23469\,
            in2 => \_gnd_net_\,
            in3 => \N__23459\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23493\,
            in2 => \N__23496\,
            in3 => \N__25061\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__27305\,
            in1 => \N__27282\,
            in2 => \_gnd_net_\,
            in3 => \N__27251\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_18_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59311\,
            ce => \N__27600\,
            sr => \N__57566\
        );

    \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__23483\,
            in1 => \N__23468\,
            in2 => \_gnd_net_\,
            in3 => \N__23458\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28605\,
            in2 => \N__23439\,
            in3 => \N__24996\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => \pid_alt.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_RNI1N2F_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32319\,
            in2 => \_gnd_net_\,
            in3 => \N__23397\,
            lcout => \pid_alt.error_1\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_0\,
            carryout => \pid_alt.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34848\,
            in2 => \_gnd_net_\,
            in3 => \N__23355\,
            lcout => \pid_alt.error_2\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_1\,
            carryout => \pid_alt.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_2_c_RNI5T4F_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34830\,
            in2 => \_gnd_net_\,
            in3 => \N__23310\,
            lcout => \pid_alt.error_3\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_2\,
            carryout => \pid_alt.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_3_c_RNIKE1T_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29658\,
            in2 => \N__23933\,
            in3 => \N__23874\,
            lcout => \pid_alt.error_4\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_3\,
            carryout => \pid_alt.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_4_c_RNINI2T_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29643\,
            in2 => \N__23871\,
            in3 => \N__23814\,
            lcout => \pid_alt.error_5\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_4\,
            carryout => \pid_alt.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_5_c_RNIQM3T_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29628\,
            in2 => \N__23811\,
            in3 => \N__23751\,
            lcout => \pid_alt.error_6\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_5\,
            carryout => \pid_alt.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_6_c_RNITQ4T_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29754\,
            in2 => \N__23748\,
            in3 => \N__23688\,
            lcout => \pid_alt.error_7\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_6\,
            carryout => \pid_alt.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_7_c_RNI9LEM_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29592\,
            in2 => \N__23685\,
            in3 => \N__23625\,
            lcout => \pid_alt.error_8\,
            ltout => OPEN,
            carryin => \bfn_2_20_0_\,
            carryout => \pid_alt.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_8_c_RNICPFM_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29607\,
            in2 => \N__23622\,
            in3 => \N__23562\,
            lcout => \pid_alt.error_9\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_8\,
            carryout => \pid_alt.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23964\,
            in2 => \N__23559\,
            in3 => \N__23499\,
            lcout => \pid_alt.error_10\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_9\,
            carryout => \pid_alt.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_10_c_RNI0SDO_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26199\,
            in2 => \N__24219\,
            in3 => \N__24162\,
            lcout => \pid_alt.error_11\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_10\,
            carryout => \pid_alt.error_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_11_c_RNI5JAH_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29706\,
            in2 => \_gnd_net_\,
            in3 => \N__24114\,
            lcout => \pid_alt.error_12\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_11\,
            carryout => \pid_alt.error_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_12_c_RNI7MBH_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29724\,
            in2 => \_gnd_net_\,
            in3 => \N__24066\,
            lcout => \pid_alt.error_13\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_12\,
            carryout => \pid_alt.error_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_13_c_RNI9PCH_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29715\,
            in2 => \_gnd_net_\,
            in3 => \N__24027\,
            lcout => \pid_alt.error_14\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_13\,
            carryout => \pid_alt.error_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_14_c_RNIBSDH_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29673\,
            in2 => \_gnd_net_\,
            in3 => \N__24024\,
            lcout => \pid_alt.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56312\,
            in2 => \_gnd_net_\,
            in3 => \N__58336\,
            lcout => alt_kp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59324\,
            ce => \N__27483\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25488\,
            lcout => drone_altitude_i_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_0_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56487\,
            in2 => \_gnd_net_\,
            in3 => \N__58334\,
            lcout => alt_kp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59329\,
            ce => \N__27484\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55723\,
            lcout => alt_kp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59329\,
            ce => \N__27484\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_5_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24363\,
            lcout => \pid_alt.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59333\,
            ce => \N__24460\,
            sr => \N__58200\
        );

    \pid_alt.error_p_reg_esr_6_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24339\,
            lcout => \pid_alt.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59333\,
            ce => \N__24460\,
            sr => \N__58200\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58333\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55581\,
            lcout => alt_kp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59336\,
            ce => \N__27489\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55377\,
            in2 => \_gnd_net_\,
            in3 => \N__58332\,
            lcout => alt_kp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59336\,
            ce => \N__27489\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_4_LC_3_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24294\,
            lcout => \pid_alt.error_d_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59127\,
            ce => \N__24448\,
            sr => \N__58216\
        );

    \Commands_frame_decoder.state_RNIRSI31_11_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__27004\,
            in1 => \N__31772\,
            in2 => \_gnd_net_\,
            in3 => \N__57860\,
            lcout => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_7_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24255\,
            lcout => \pid_alt.error_d_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59182\,
            ce => \N__24452\,
            sr => \N__58214\
        );

    \pid_alt.error_d_reg_esr_8_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24243\,
            lcout => \pid_alt.error_d_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59182\,
            ce => \N__24452\,
            sr => \N__58214\
        );

    \pid_alt.error_d_reg_esr_9_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24231\,
            lcout => \pid_alt.error_d_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59182\,
            ce => \N__24452\,
            sr => \N__58214\
        );

    \pid_alt.error_i_reg_esr_0_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24498\,
            lcout => \pid_alt.error_i_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59182\,
            ce => \N__24452\,
            sr => \N__58214\
        );

    \pid_alt.error_i_reg_esr_3_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24486\,
            lcout => \pid_alt.error_i_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59182\,
            ce => \N__24452\,
            sr => \N__58214\
        );

    \pid_alt.error_i_reg_esr_11_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24474\,
            lcout => \pid_alt.error_i_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59182\,
            ce => \N__24452\,
            sr => \N__58214\
        );

    \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__55284\,
            in1 => \N__56074\,
            in2 => \_gnd_net_\,
            in3 => \N__56266\,
            lcout => \Commands_frame_decoder.source_CH1data8lt7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_14_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59211\,
            ce => \N__27613\,
            sr => \N__57511\
        );

    \pid_alt.error_d_reg_prev_esr_0_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24391\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59226\,
            ce => \N__27610\,
            sr => \N__57515\
        );

    \pid_alt.error_i_acumm_prereg_esr_20_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27199\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59226\,
            ce => \N__27610\,
            sr => \N__57515\
        );

    \pid_alt.error_d_reg_prev_esr_3_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24609\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59226\,
            ce => \N__27610\,
            sr => \N__57515\
        );

    \pid_alt.error_i_acumm_prereg_esr_18_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24995\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59226\,
            ce => \N__27610\,
            sr => \N__57515\
        );

    \pid_alt.error_i_acumm_prereg_esr_19_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25062\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59226\,
            ce => \N__27610\,
            sr => \N__57515\
        );

    \pid_alt.error_i_acumm_prereg_esr_13_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24831\,
            lcout => \pid_alt.error_i_acumm7lto13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59226\,
            ce => \N__27610\,
            sr => \N__57515\
        );

    \pid_alt.error_i_acumm_prereg_esr_1_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25289\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59226\,
            ce => \N__27610\,
            sr => \N__57515\
        );

    \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24557\,
            in1 => \N__24567\,
            in2 => \N__25242\,
            in3 => \N__25705\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24663\,
            in1 => \N__24626\,
            in2 => \_gnd_net_\,
            in3 => \N__24608\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__24558\,
            in1 => \_gnd_net_\,
            in2 => \N__24561\,
            in3 => \N__25706\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24548\,
            in1 => \N__24506\,
            in2 => \_gnd_net_\,
            in3 => \N__24523\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__24524\,
            in1 => \_gnd_net_\,
            in2 => \N__24510\,
            in3 => \N__24549\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__25187\,
            in1 => \N__24770\,
            in2 => \N__24528\,
            in3 => \N__25744\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_4_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59243\,
            ce => \N__27607\,
            sr => \N__57521\
        );

    \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__24777\,
            in1 => \N__24771\,
            in2 => \_gnd_net_\,
            in3 => \N__25745\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25814\,
            in2 => \N__25647\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.un1_pid_prereg_0\,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24762\,
            in2 => \N__25836\,
            in3 => \N__24756\,
            lcout => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25776\,
            in2 => \N__24753\,
            in3 => \N__24738\,
            lcout => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25842\,
            in2 => \N__24735\,
            in3 => \N__24723\,
            lcout => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25803\,
            in2 => \N__24720\,
            in3 => \N__24702\,
            lcout => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33366\,
            in2 => \N__24699\,
            in3 => \N__24684\,
            lcout => \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26039\,
            in2 => \N__24681\,
            in3 => \N__24666\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26024\,
            in2 => \N__24969\,
            in3 => \N__24954\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26009\,
            in2 => \N__24951\,
            in3 => \N__24936\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25997\,
            in2 => \N__24933\,
            in3 => \N__24918\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26066\,
            in2 => \N__24915\,
            in3 => \N__24897\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26051\,
            in2 => \N__24894\,
            in3 => \N__24870\,
            lcout => \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25973\,
            in2 => \N__24867\,
            in3 => \N__24852\,
            lcout => \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27960\,
            in2 => \N__24849\,
            in3 => \N__24810\,
            lcout => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24807\,
            in2 => \_gnd_net_\,
            in3 => \N__24795\,
            lcout => \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24792\,
            in3 => \N__25134\,
            lcout => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25131\,
            in2 => \_gnd_net_\,
            in3 => \N__25116\,
            lcout => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25113\,
            in2 => \_gnd_net_\,
            in3 => \N__25098\,
            lcout => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25095\,
            in2 => \_gnd_net_\,
            in3 => \N__25080\,
            lcout => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25077\,
            in2 => \_gnd_net_\,
            in3 => \N__25035\,
            lcout => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25028\,
            in2 => \_gnd_net_\,
            in3 => \N__25032\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25029\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25011\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25008\,
            in1 => \N__28604\,
            in2 => \N__26562\,
            in3 => \N__24985\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26232\,
            in1 => \N__26211\,
            in2 => \_gnd_net_\,
            in3 => \N__27647\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34904\,
            in2 => \N__34911\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_0_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25335\,
            in2 => \N__25326\,
            in3 => \N__25305\,
            lcout => \pid_alt.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_0\,
            clk => \N__59298\,
            ce => \N__27601\,
            sr => \N__57547\
        );

    \pid_alt.pid_prereg_esr_1_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25302\,
            in2 => \N__25290\,
            in3 => \N__25272\,
            lcout => \pid_alt.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_0\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_1\,
            clk => \N__59298\,
            ce => \N__27601\,
            sr => \N__57547\
        );

    \pid_alt.pid_prereg_esr_2_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25269\,
            in2 => \N__25731\,
            in3 => \N__25260\,
            lcout => \pid_alt.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_1\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_2\,
            clk => \N__59298\,
            ce => \N__27601\,
            sr => \N__57547\
        );

    \pid_alt.pid_prereg_esr_3_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25257\,
            in2 => \N__25868\,
            in3 => \N__25245\,
            lcout => \pid_alt.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_2\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_3\,
            clk => \N__59298\,
            ce => \N__27601\,
            sr => \N__57547\
        );

    \pid_alt.pid_prereg_esr_4_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25238\,
            in2 => \N__25218\,
            in3 => \N__25206\,
            lcout => \pid_alt.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_3\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_4\,
            clk => \N__59298\,
            ce => \N__27601\,
            sr => \N__57547\
        );

    \pid_alt.pid_prereg_esr_5_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25203\,
            in2 => \N__25194\,
            in3 => \N__25173\,
            lcout => \pid_alt.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_4\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_5\,
            clk => \N__59298\,
            ce => \N__27601\,
            sr => \N__57547\
        );

    \pid_alt.pid_prereg_esr_6_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25170\,
            in2 => \N__25158\,
            in3 => \N__25137\,
            lcout => \pid_alt.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_5\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_6\,
            clk => \N__59298\,
            ce => \N__27601\,
            sr => \N__57547\
        );

    \pid_alt.pid_prereg_esr_7_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26610\,
            in2 => \N__26663\,
            in3 => \N__25422\,
            lcout => \pid_alt.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_7\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_8_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26346\,
            in2 => \N__26750\,
            in3 => \N__25419\,
            lcout => \pid_alt.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_7\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_8\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_9_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26091\,
            in2 => \N__26330\,
            in3 => \N__25416\,
            lcout => \pid_alt.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_8\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_9\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_10_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26220\,
            in2 => \N__26187\,
            in3 => \N__25413\,
            lcout => \pid_alt.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_9\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_10\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_11_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25410\,
            in2 => \N__25401\,
            in3 => \N__25380\,
            lcout => \pid_alt.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_10\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_11\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_12_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25377\,
            in2 => \N__25371\,
            in3 => \N__25353\,
            lcout => \pid_alt.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_11\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_12\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_13_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25350\,
            in2 => \N__25898\,
            in3 => \N__25344\,
            lcout => \pid_alt.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_12\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_13\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_14_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26418\,
            in2 => \N__26438\,
            in3 => \N__25341\,
            lcout => \pid_alt.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_13\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_14\,
            clk => \N__59306\,
            ce => \N__27599\,
            sr => \N__57557\
        );

    \pid_alt.pid_prereg_esr_15_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26082\,
            in2 => \N__26370\,
            in3 => \N__25338\,
            lcout => \pid_alt.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_15\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_16_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26838\,
            in2 => \N__26889\,
            in3 => \N__25482\,
            lcout => \pid_alt.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_15\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_16\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_17_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26963\,
            in2 => \N__26604\,
            in3 => \N__25479\,
            lcout => \pid_alt.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_16\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_17\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_18_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25476\,
            in2 => \N__26561\,
            in3 => \N__25467\,
            lcout => \pid_alt.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_17\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_18\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_19_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25464\,
            in2 => \N__25457\,
            in3 => \N__25440\,
            lcout => \pid_alt.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_18\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_19\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_20_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27177\,
            in2 => \N__27221\,
            in3 => \N__25437\,
            lcout => \pid_alt.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_19\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_20\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_21_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27018\,
            in2 => \N__27102\,
            in3 => \N__25434\,
            lcout => \pid_alt.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_20\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_21\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_22_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25524\,
            in2 => \N__25506\,
            in3 => \N__25431\,
            lcout => \pid_alt.pid_preregZ0Z_22\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_21\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_22\,
            clk => \N__59312\,
            ce => \N__27597\,
            sr => \N__57567\
        );

    \pid_alt.pid_prereg_esr_23_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25502\,
            in2 => \N__25515\,
            in3 => \N__25428\,
            lcout => \pid_alt.pid_preregZ0Z_23\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_23\,
            clk => \N__59317\,
            ce => \N__27595\,
            sr => \N__57575\
        );

    \pid_alt.pid_prereg_esr_24_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000101111110"
        )
    port map (
            in0 => \N__27086\,
            in1 => \N__27053\,
            in2 => \N__27123\,
            in3 => \N__25425\,
            lcout => \pid_alt.pid_preregZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59317\,
            ce => \N__27595\,
            sr => \N__57575\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__26813\,
            in1 => \N__26828\,
            in2 => \_gnd_net_\,
            in3 => \N__26786\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_8_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26787\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59320\,
            ce => \N__27593\,
            sr => \N__57582\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__25599\,
            in1 => \N__25538\,
            in2 => \_gnd_net_\,
            in3 => \N__25574\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_13_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25575\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59320\,
            ce => \N__27593\,
            sr => \N__57582\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27117\,
            in1 => \N__27081\,
            in2 => \_gnd_net_\,
            in3 => \N__27049\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__27051\,
            in1 => \_gnd_net_\,
            in2 => \N__27087\,
            in3 => \N__27119\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__27118\,
            in1 => \N__27082\,
            in2 => \_gnd_net_\,
            in3 => \N__27050\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_21_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59320\,
            ce => \N__27593\,
            sr => \N__57582\
        );

    \dron_frame_decoder_1.source_Altitude_esr_10_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50394\,
            lcout => \dron_frame_decoder_1.drone_altitude_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59325\,
            ce => \N__30861\,
            sr => \N__57593\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_2_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56141\,
            in2 => \_gnd_net_\,
            in3 => \N__58331\,
            lcout => alt_kp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59330\,
            ce => \N__27488\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55922\,
            in2 => \_gnd_net_\,
            in3 => \N__58330\,
            lcout => alt_kp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59330\,
            ce => \N__27488\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_11_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__31674\,
            in1 => \N__29351\,
            in2 => \N__27012\,
            in3 => \N__31315\,
            lcout => \Commands_frame_decoder.stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59141\,
            ce => 'H',
            sr => \N__57497\
        );

    \Commands_frame_decoder.state_2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__31316\,
            in1 => \N__31679\,
            in2 => \N__25667\,
            in3 => \N__27345\,
            lcout => \Commands_frame_decoder.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59170\,
            ce => 'H',
            sr => \N__57501\
        );

    \pid_alt.error_d_reg_prev_esr_15_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38527\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59183\,
            ce => \N__27614\,
            sr => \N__57503\
        );

    \pid_alt.error_d_reg_prev_esr_17_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59199\,
            ce => \N__27611\,
            sr => \N__57508\
        );

    \pid_alt.error_i_acumm_prereg_esr_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25643\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59199\,
            ce => \N__27611\,
            sr => \N__57508\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25623\,
            in1 => \N__25764\,
            in2 => \N__25617\,
            in3 => \N__25770\,
            lcout => OPEN,
            ltout => \pid_alt.m7_e_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__25608\,
            in1 => \N__25752\,
            in2 => \N__25602\,
            in3 => \N__25758\,
            lcout => \pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_16_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26865\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59212\,
            ce => \N__27608\,
            sr => \N__57512\
        );

    \pid_alt.error_i_acumm_prereg_esr_17_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26586\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59212\,
            ce => \N__27608\,
            sr => \N__57512\
        );

    \pid_alt.error_i_acumm_prereg_esr_14_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26391\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59212\,
            ce => \N__27608\,
            sr => \N__57512\
        );

    \pid_alt.error_i_acumm_prereg_esr_15_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26529\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_i_acumm_prereg_esr_12_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25923\,
            lcout => \pid_alt.error_i_acumm7lto12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_i_acumm_prereg_esr_5_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25746\,
            lcout => \pid_alt.error_i_acumm7lto5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_d_reg_prev_esr_9_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26169\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_i_acumm_prereg_esr_7_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26624\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_i_acumm_prereg_esr_2_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25726\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_i_acumm_prereg_esr_4_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25707\,
            lcout => \pid_alt.error_i_acumm7lto4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_i_acumm_prereg_esr_3_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25861\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59227\,
            ce => \N__27605\,
            sr => \N__57516\
        );

    \pid_alt.error_i_acumm_esr_3_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__33388\,
            in1 => \N__27900\,
            in2 => \N__25797\,
            in3 => \N__27378\,
            lcout => \pid_alt.error_i_acummZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59244\,
            ce => \N__27951\,
            sr => \N__33338\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27394\,
            in1 => \_gnd_net_\,
            in2 => \N__33428\,
            in3 => \N__33385\,
            lcout => \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_1_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__33386\,
            in1 => \N__27720\,
            in2 => \N__25796\,
            in3 => \N__27904\,
            lcout => \pid_alt.error_i_acummZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59244\,
            ce => \N__27951\,
            sr => \N__33338\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__28039\,
            in1 => \N__28006\,
            in2 => \_gnd_net_\,
            in3 => \N__27983\,
            lcout => \pid_alt.N_9_0\,
            ltout => \pid_alt.N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27873\,
            in1 => \N__25986\,
            in2 => \N__25824\,
            in3 => \N__27393\,
            lcout => \pid_alt.N_62_mux\,
            ltout => \pid_alt.N_62_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_0_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__27702\,
            in1 => \N__27896\,
            in2 => \N__25821\,
            in3 => \N__25788\,
            lcout => \pid_alt.error_i_acummZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59244\,
            ce => \N__27951\,
            sr => \N__33338\
        );

    \pid_alt.error_i_acumm_esr_4_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110111"
        )
    port map (
            in0 => \N__33389\,
            in1 => \N__33424\,
            in2 => \N__27905\,
            in3 => \N__27395\,
            lcout => \pid_alt.error_i_acummZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59244\,
            ce => \N__27951\,
            sr => \N__33338\
        );

    \pid_alt.error_i_acumm_esr_2_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__27366\,
            in1 => \N__25792\,
            in2 => \N__27906\,
            in3 => \N__33387\,
            lcout => \pid_alt.error_i_acummZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59244\,
            ce => \N__27951\,
            sr => \N__33338\
        );

    \pid_alt.error_i_acumm_10_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111010"
        )
    port map (
            in0 => \N__39731\,
            in1 => \N__27630\,
            in2 => \N__26070\,
            in3 => \N__27409\,
            lcout => \pid_alt.error_i_acummZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59260\,
            ce => 'H',
            sr => \N__33331\
        );

    \pid_alt.error_i_acumm_11_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__27410\,
            in1 => \N__27766\,
            in2 => \N__26055\,
            in3 => \N__39735\,
            lcout => \pid_alt.error_i_acummZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59260\,
            ce => 'H',
            sr => \N__33331\
        );

    \pid_alt.error_i_acumm_6_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__26040\,
            in1 => \N__27735\,
            in2 => \N__39738\,
            in3 => \N__27411\,
            lcout => \pid_alt.error_i_acummZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59260\,
            ce => 'H',
            sr => \N__33331\
        );

    \pid_alt.error_i_acumm_7_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__27412\,
            in1 => \N__27933\,
            in2 => \N__26028\,
            in3 => \N__39736\,
            lcout => \pid_alt.error_i_acummZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59260\,
            ce => 'H',
            sr => \N__33331\
        );

    \pid_alt.error_i_acumm_8_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011111100"
        )
    port map (
            in0 => \N__27783\,
            in1 => \N__39730\,
            in2 => \N__26013\,
            in3 => \N__27413\,
            lcout => \pid_alt.error_i_acummZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59260\,
            ce => 'H',
            sr => \N__33331\
        );

    \pid_alt.error_i_acumm_9_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__27414\,
            in1 => \N__25998\,
            in2 => \N__27801\,
            in3 => \N__39737\,
            lcout => \pid_alt.error_i_acummZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59260\,
            ce => 'H',
            sr => \N__33331\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27932\,
            in2 => \_gnd_net_\,
            in3 => \N__27734\,
            lcout => \pid_alt.m35_e_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_12_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__39729\,
            in1 => \N__27681\,
            in2 => \N__25977\,
            in3 => \N__28077\,
            lcout => \pid_alt.error_i_acummZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59260\,
            ce => 'H',
            sr => \N__33331\
        );

    \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__25962\,
            in1 => \N__25950\,
            in2 => \_gnd_net_\,
            in3 => \N__25918\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__26313\,
            in1 => \N__26286\,
            in2 => \_gnd_net_\,
            in3 => \N__26271\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__26183\,
            in1 => \N__26210\,
            in2 => \N__26223\,
            in3 => \N__27646\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__26132\,
            in1 => \N__26144\,
            in2 => \_gnd_net_\,
            in3 => \N__26167\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29445\,
            lcout => drone_altitude_i_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26109\,
            in1 => \N__26115\,
            in2 => \_gnd_net_\,
            in3 => \N__27815\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__26168\,
            in1 => \_gnd_net_\,
            in2 => \N__26148\,
            in3 => \N__26133\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__26108\,
            in1 => \N__26331\,
            in2 => \N__26094\,
            in3 => \N__27814\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26507\,
            in1 => \N__26538\,
            in2 => \N__26366\,
            in3 => \N__26524\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__26481\,
            in1 => \N__26499\,
            in2 => \_gnd_net_\,
            in3 => \N__26462\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__26508\,
            in1 => \_gnd_net_\,
            in2 => \N__26532\,
            in3 => \N__26525\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__38486\,
            in1 => \N__38453\,
            in2 => \_gnd_net_\,
            in3 => \N__38529\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__26498\,
            in1 => \N__26480\,
            in2 => \_gnd_net_\,
            in3 => \N__26461\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__26439\,
            in1 => \N__26405\,
            in2 => \N__26421\,
            in3 => \N__26386\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26412\,
            in1 => \N__26406\,
            in2 => \_gnd_net_\,
            in3 => \N__26387\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26759\,
            in1 => \N__26340\,
            in2 => \N__26751\,
            in3 => \N__27865\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__26699\,
            in1 => \N__26708\,
            in2 => \_gnd_net_\,
            in3 => \N__26731\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__26760\,
            in1 => \_gnd_net_\,
            in2 => \N__26334\,
            in3 => \N__27866\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__26829\,
            in1 => \N__26814\,
            in2 => \_gnd_net_\,
            in3 => \N__26780\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_7_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26733\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59299\,
            ce => \N__27598\,
            sr => \N__57548\
        );

    \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26679\,
            in1 => \N__26685\,
            in2 => \_gnd_net_\,
            in3 => \N__26631\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__26732\,
            in1 => \_gnd_net_\,
            in2 => \N__26712\,
            in3 => \N__26700\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__26678\,
            in1 => \N__26664\,
            in2 => \N__26634\,
            in3 => \N__26630\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26595\,
            in1 => \N__26975\,
            in2 => \N__26967\,
            in3 => \N__26584\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__28661\,
            in1 => \N__28685\,
            in2 => \_gnd_net_\,
            in3 => \N__28640\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26976\,
            in2 => \N__26589\,
            in3 => \N__26585\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__26912\,
            in1 => \N__26921\,
            in2 => \_gnd_net_\,
            in3 => \N__26950\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_16_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59307\,
            ce => \N__27596\,
            sr => \N__57558\
        );

    \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26895\,
            in1 => \N__38430\,
            in2 => \_gnd_net_\,
            in3 => \N__26864\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__26951\,
            in1 => \_gnd_net_\,
            in2 => \N__26925\,
            in3 => \N__26913\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__26888\,
            in1 => \N__38429\,
            in2 => \N__26868\,
            in3 => \N__26863\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__27170\,
            in1 => \N__27155\,
            in2 => \_gnd_net_\,
            in3 => \N__27145\,
            lcout => \pid_alt.un1_pid_prereg_236_1\,
            ltout => \pid_alt.un1_pid_prereg_236_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27231\,
            in2 => \N__26832\,
            in3 => \N__27201\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_20_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27147\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59313\,
            ce => \N__27594\,
            sr => \N__57568\
        );

    \pid_alt.error_d_reg_prev_esr_19_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59313\,
            ce => \N__27594\,
            sr => \N__57568\
        );

    \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__27306\,
            in1 => \N__27275\,
            in2 => \_gnd_net_\,
            in3 => \N__27260\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__27225\,
            in1 => \N__27079\,
            in2 => \N__27204\,
            in3 => \N__27200\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__27171\,
            in1 => \N__27156\,
            in2 => \_gnd_net_\,
            in3 => \N__27146\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__27101\,
            in1 => \N__27080\,
            in2 => \N__27057\,
            in3 => \N__27054\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_12_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__27011\,
            in1 => \N__26987\,
            in2 => \N__31738\,
            in3 => \N__31290\,
            lcout => \Commands_frame_decoder.stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59128\,
            ce => 'H',
            sr => \N__57496\
        );

    \Commands_frame_decoder.state_13_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__31291\,
            in1 => \N__31804\,
            in2 => \N__26988\,
            in3 => \N__31678\,
            lcout => \Commands_frame_decoder.stateZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59128\,
            ce => 'H',
            sr => \N__57496\
        );

    \uart_pc.data_rdy_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30344\,
            in2 => \_gnd_net_\,
            in3 => \N__29292\,
            lcout => uart_pc_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59142\,
            ce => 'H',
            sr => \N__57498\
        );

    \Commands_frame_decoder.state_RNO_1_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__27332\,
            in1 => \N__27539\,
            in2 => \N__29067\,
            in3 => \N__27507\,
            lcout => \Commands_frame_decoder.N_377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56224\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_0_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__55705\,
            in1 => \N__31655\,
            in2 => \N__27351\,
            in3 => \N__55332\,
            lcout => \Commands_frame_decoder.N_416\,
            ltout => \Commands_frame_decoder.N_416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_2_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__27339\,
            in1 => \N__55846\,
            in2 => \N__27348\,
            in3 => \N__56046\,
            lcout => \Commands_frame_decoder.N_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNI6QPK_1_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31831\,
            in2 => \_gnd_net_\,
            in3 => \N__27523\,
            lcout => \Commands_frame_decoder.N_376_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_1_2_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__56433\,
            in1 => \N__27522\,
            in2 => \_gnd_net_\,
            in3 => \N__55521\,
            lcout => \Commands_frame_decoder.state_ns_0_a3_0_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__31304\,
            in1 => \N__31726\,
            in2 => \N__29198\,
            in3 => \N__27333\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.N_376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29268\,
            in1 => \N__27321\,
            in2 => \N__27315\,
            in3 => \N__27312\,
            lcout => \Commands_frame_decoder.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59171\,
            ce => 'H',
            sr => \N__57502\
        );

    \Commands_frame_decoder.state_14_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__31808\,
            in1 => \N__29267\,
            in2 => \_gnd_net_\,
            in3 => \N__31727\,
            lcout => \Commands_frame_decoder.stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59171\,
            ce => 'H',
            sr => \N__57502\
        );

    \Commands_frame_decoder.state_RNIOMNA5_1_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__31725\,
            in1 => \N__27525\,
            in2 => \_gnd_net_\,
            in3 => \N__31303\,
            lcout => \Commands_frame_decoder.N_379\,
            ltout => \Commands_frame_decoder.N_379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__29178\,
            in1 => \N__27540\,
            in2 => \N__27528\,
            in3 => \N__55549\,
            lcout => \Commands_frame_decoder.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59171\,
            ce => 'H',
            sr => \N__57502\
        );

    \Commands_frame_decoder.state_RNO_2_0_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__27524\,
            in1 => \N__56440\,
            in2 => \N__56106\,
            in3 => \N__29159\,
            lcout => \Commands_frame_decoder.N_412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_9_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__31314\,
            in1 => \N__27497\,
            in2 => \N__31774\,
            in3 => \N__27426\,
            lcout => \Commands_frame_decoder.stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59184\,
            ce => 'H',
            sr => \N__57504\
        );

    \Commands_frame_decoder.state_8_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__29391\,
            in1 => \N__31728\,
            in2 => \N__27501\,
            in3 => \N__31313\,
            lcout => \Commands_frame_decoder.stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59184\,
            ce => 'H',
            sr => \N__57504\
        );

    \Commands_frame_decoder.state_RNIF38S_6_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__29550\,
            in1 => \N__31778\,
            in2 => \_gnd_net_\,
            in3 => \N__57837\,
            lcout => \Commands_frame_decoder.state_RNIF38SZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNILP1J_9_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27425\,
            in2 => \_gnd_net_\,
            in3 => \N__31777\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__28013\,
            in1 => \N__27677\,
            in2 => \N__28059\,
            in3 => \N__27979\,
            lcout => \pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27377\,
            in2 => \_gnd_net_\,
            in3 => \N__27362\,
            lcout => OPEN,
            ltout => \pid_alt.m21_e_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27925\,
            in1 => \N__33420\,
            in2 => \N__27909\,
            in3 => \N__27895\,
            lcout => \pid_alt.m21_e_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27797\,
            in1 => \N__27782\,
            in2 => \N__27768\,
            in3 => \N__27629\,
            lcout => \pid_alt.m35_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_8_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27867\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59228\,
            ce => \N__27603\,
            sr => \N__57517\
        );

    \pid_alt.error_i_acumm_prereg_esr_6_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27840\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59228\,
            ce => \N__27603\,
            sr => \N__57517\
        );

    \pid_alt.error_i_acumm_prereg_esr_9_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27822\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59228\,
            ce => \N__27603\,
            sr => \N__57517\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27796\,
            in1 => \N__27781\,
            in2 => \N__27767\,
            in3 => \N__27733\,
            lcout => OPEN,
            ltout => \pid_alt.m21_e_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIEK7C2_0_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27719\,
            in1 => \N__27701\,
            in2 => \N__27684\,
            in3 => \N__27660\,
            lcout => \pid_alt.m21_e_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27628\,
            in2 => \_gnd_net_\,
            in3 => \N__27676\,
            lcout => \pid_alt.m21_e_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_10_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27654\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59228\,
            ce => \N__27603\,
            sr => \N__57517\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28092\,
            in1 => \N__28083\,
            in2 => \N__28058\,
            in3 => \N__28076\,
            lcout => OPEN,
            ltout => \pid_alt.error_i_acumm_prereg_esr_RNIO7B05Z0Z_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIAAPN5_1_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__39720\,
            in1 => \_gnd_net_\,
            in2 => \N__28065\,
            in3 => \N__44979\,
            lcout => \pid_alt.un1_reset_1_0_i\,
            ltout => \pid_alt.un1_reset_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIVV066_1_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28062\,
            in3 => \N__39721\,
            lcout => \pid_alt.N_72_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_13_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__28054\,
            in1 => \N__28014\,
            in2 => \_gnd_net_\,
            in3 => \N__27987\,
            lcout => \pid_alt.error_i_acummZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59245\,
            ce => \N__27950\,
            sr => \N__33330\
        );

    \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__39719\,
            in1 => \N__44978\,
            in2 => \N__28910\,
            in3 => \N__28545\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__28320\,
            in1 => \N__28960\,
            in2 => \N__27939\,
            in3 => \N__28832\,
            lcout => \pid_alt.un1_reset_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__28961\,
            in1 => \N__28899\,
            in2 => \N__28779\,
            in3 => \N__28833\,
            lcout => \pid_alt.source_pid_9_0_tz_6\,
            ltout => \pid_alt.source_pid_9_0_tz_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_10_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001001110"
        )
    port map (
            in0 => \N__39723\,
            in1 => \N__34717\,
            in2 => \N__27936\,
            in3 => \N__28257\,
            lcout => throttle_order_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59261\,
            ce => 'H',
            sr => \N__28708\
        );

    \pid_alt.source_pid_1_11_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__28148\,
            in1 => \N__39726\,
            in2 => \N__40045\,
            in3 => \N__28305\,
            lcout => throttle_order_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59261\,
            ce => 'H',
            sr => \N__28708\
        );

    \pid_alt.source_pid_1_6_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__39724\,
            in1 => \N__28149\,
            in2 => \N__36124\,
            in3 => \N__28179\,
            lcout => throttle_order_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59261\,
            ce => 'H',
            sr => \N__28708\
        );

    \pid_alt.source_pid_1_7_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__28150\,
            in1 => \N__39727\,
            in2 => \N__36215\,
            in3 => \N__28206\,
            lcout => throttle_order_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59261\,
            ce => 'H',
            sr => \N__28708\
        );

    \pid_alt.source_pid_1_8_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__39725\,
            in1 => \N__28151\,
            in2 => \N__35971\,
            in3 => \N__28230\,
            lcout => throttle_order_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59261\,
            ce => 'H',
            sr => \N__28708\
        );

    \pid_alt.source_pid_1_9_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__28152\,
            in1 => \N__39728\,
            in2 => \N__36058\,
            in3 => \N__28281\,
            lcout => throttle_order_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59261\,
            ce => 'H',
            sr => \N__28708\
        );

    \pid_alt.state_RNIOVDUE_1_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__39722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28699\,
            lcout => \pid_alt.N_72_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28103\,
            in1 => \N__28130\,
            in2 => \N__28119\,
            in3 => \N__28337\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_2_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__28835\,
            in1 => \N__28349\,
            in2 => \N__28134\,
            in3 => \N__28901\,
            lcout => throttle_order_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59275\,
            ce => \N__28730\,
            sr => \N__28715\
        );

    \pid_alt.source_pid_1_esr_3_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__28118\,
            in1 => \N__28906\,
            in2 => \N__28353\,
            in3 => \N__28837\,
            lcout => throttle_order_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59275\,
            ce => \N__28730\,
            sr => \N__28715\
        );

    \pid_alt.source_pid_1_esr_1_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__28834\,
            in1 => \N__28348\,
            in2 => \N__28911\,
            in3 => \N__28104\,
            lcout => throttle_order_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59275\,
            ce => \N__28730\,
            sr => \N__28715\
        );

    \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__28959\,
            in1 => \N__28774\,
            in2 => \_gnd_net_\,
            in3 => \N__28557\,
            lcout => \pid_alt.N_44\,
            ltout => \pid_alt.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__28415\,
            in1 => \_gnd_net_\,
            in2 => \N__28356\,
            in3 => \N__28388\,
            lcout => \pid_alt.N_46\,
            ltout => \pid_alt.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_0_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__28900\,
            in1 => \N__28338\,
            in2 => \N__28326\,
            in3 => \N__28836\,
            lcout => throttle_order_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59275\,
            ce => \N__28730\,
            sr => \N__28715\
        );

    \pid_front.error_d_reg_esr_RNI1VUF_9_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__30774\,
            in1 => \N__32304\,
            in2 => \N__56775\,
            in3 => \N__32271\,
            lcout => \pid_front.error_d_reg_esr_RNI1VUFZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__28252\,
            in1 => \N__28311\,
            in2 => \N__28205\,
            in3 => \N__39678\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__28390\,
            in1 => \N__28569\,
            in2 => \N__28323\,
            in3 => \N__28414\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28226\,
            in1 => \N__28178\,
            in2 => \N__28280\,
            in3 => \N__28301\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI8H141_10_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__28300\,
            in1 => \N__28273\,
            in2 => \N__28256\,
            in3 => \N__28225\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__28198\,
            in1 => \_gnd_net_\,
            in2 => \N__28182\,
            in3 => \N__28177\,
            lcout => \pid_alt.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__28764\,
            in1 => \N__28991\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.N_90\,
            ltout => \pid_alt.N_90_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39677\,
            in1 => \N__28389\,
            in2 => \N__28572\,
            in3 => \N__28941\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__28808\,
            in1 => \N__28568\,
            in2 => \N__28560\,
            in3 => \N__28556\,
            lcout => \pid_alt.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28536\,
            in1 => \N__28527\,
            in2 => \N__28515\,
            in3 => \N__28500\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28491\,
            in1 => \N__28479\,
            in2 => \N__28470\,
            in3 => \N__28458\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__28449\,
            in1 => \N__28443\,
            in2 => \N__28431\,
            in3 => \N__28428\,
            lcout => \pid_alt.N_305\,
            ltout => \pid_alt.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__28391\,
            in1 => \N__28419\,
            in2 => \N__28398\,
            in3 => \N__28902\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_9_0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_4_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__29004\,
            in1 => \N__28825\,
            in2 => \N__28395\,
            in3 => \N__28392\,
            lcout => throttle_order_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59300\,
            ce => \N__28731\,
            sr => \N__28716\
        );

    \pid_alt.source_pid_1_esr_5_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__28905\,
            in1 => \N__29003\,
            in2 => \N__28839\,
            in3 => \N__28992\,
            lcout => throttle_order_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59300\,
            ce => \N__28731\,
            sr => \N__28716\
        );

    \pid_alt.source_pid_1_esr_13_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__28904\,
            in1 => \N__28824\,
            in2 => \_gnd_net_\,
            in3 => \N__28967\,
            lcout => throttle_order_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59300\,
            ce => \N__28731\,
            sr => \N__28716\
        );

    \pid_alt.source_pid_1_esr_12_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__28968\,
            in1 => \N__28903\,
            in2 => \N__28838\,
            in3 => \N__28778\,
            lcout => throttle_order_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59300\,
            ce => \N__28731\,
            sr => \N__28716\
        );

    \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__28686\,
            in1 => \N__28665\,
            in2 => \_gnd_net_\,
            in3 => \N__28644\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.un1_state57_i_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31771\,
            in2 => \_gnd_net_\,
            in3 => \N__57851\,
            lcout => \Commands_frame_decoder.un1_state57_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIRP8S_1_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__29085\,
            in1 => \N__29036\,
            in2 => \N__29088\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \uart_pc.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29136\,
            in2 => \_gnd_net_\,
            in3 => \N__28581\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_1\,
            carryout => \uart_pc.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29881\,
            in2 => \_gnd_net_\,
            in3 => \N__28578\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_2\,
            carryout => \uart_pc.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_4_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29919\,
            in2 => \_gnd_net_\,
            in3 => \N__28575\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29037\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_4_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__57881\,
            in1 => \N__29992\,
            in2 => \N__29118\,
            in3 => \N__29049\,
            lcout => \uart_pc.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__29043\,
            in1 => \N__29110\,
            in2 => \N__29998\,
            in3 => \N__57882\,
            lcout => \uart_pc.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_3_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__57880\,
            in1 => \N__29991\,
            in2 => \N__29117\,
            in3 => \N__29028\,
            lcout => \uart_pc.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNI5UFA2_3_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30620\,
            in1 => \N__29930\,
            in2 => \_gnd_net_\,
            in3 => \N__29878\,
            lcout => \uart_pc.N_144_1\,
            ltout => \uart_pc.N_144_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_4_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__30237\,
            in1 => \N__29108\,
            in2 => \N__29022\,
            in3 => \N__44951\,
            lcout => \uart_pc.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIBLRB2_4_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__29967\,
            in1 => \N__30029\,
            in2 => \N__29019\,
            in3 => \N__30236\,
            lcout => \uart_pc.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__29876\,
            in1 => \N__29134\,
            in2 => \N__29937\,
            in3 => \N__29965\,
            lcout => \uart_pc.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_2_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__29109\,
            in1 => \N__29010\,
            in2 => \N__30003\,
            in3 => \N__57869\,
            lcout => \uart_pc.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIVT8S_2_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29135\,
            lcout => \uart_pc.N_126_li\,
            ltout => \uart_pc.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIMQ8T1_4_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__29966\,
            in1 => \N__29931\,
            in2 => \N__29121\,
            in3 => \N__57867\,
            lcout => \uart_pc.N_143\,
            ltout => \uart_pc.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__57868\,
            in1 => \N__29999\,
            in2 => \N__29091\,
            in3 => \N__29087\,
            lcout => \uart_pc.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__29251\,
            in1 => \N__30411\,
            in2 => \N__29228\,
            in3 => \N__55818\,
            lcout => uart_pc_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__56388\,
            in1 => \N__29218\,
            in2 => \N__30108\,
            in3 => \N__29250\,
            lcout => uart_pc_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_3_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__56001\,
            in1 => \N__55446\,
            in2 => \N__56441\,
            in3 => \N__55817\,
            lcout => \Commands_frame_decoder.state_ns_i_a2_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNILR1B2_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__29287\,
            in1 => \N__30326\,
            in2 => \_gnd_net_\,
            in3 => \N__57861\,
            lcout => \uart_pc.timer_Count_RNILR1B2Z0Z_2\,
            ltout => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_4_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__30422\,
            in1 => \N__29288\,
            in2 => \N__29052\,
            in3 => \N__53324\,
            lcout => uart_pc_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__30074\,
            in1 => \N__29222\,
            in2 => \N__56073\,
            in3 => \N__29253\,
            lcout => uart_pc_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29286\,
            in2 => \_gnd_net_\,
            in3 => \N__44970\,
            lcout => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\,
            ltout => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__30089\,
            in1 => \N__29252\,
            in2 => \N__29271\,
            in3 => \N__56220\,
            lcout => uart_pc_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNISEFT5_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001001100"
        )
    port map (
            in0 => \N__31763\,
            in1 => \N__31840\,
            in2 => \N__31866\,
            in3 => \N__31269\,
            lcout => \Commands_frame_decoder.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_5_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__29255\,
            in1 => \N__30392\,
            in2 => \N__29229\,
            in3 => \N__55666\,
            lcout => uart_pc_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_3_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__55280\,
            in1 => \N__29223\,
            in2 => \N__30060\,
            in3 => \N__29254\,
            lcout => uart_pc_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_6_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__30278\,
            in1 => \N__29256\,
            in2 => \N__55534\,
            in3 => \N__29227\,
            lcout => uart_pc_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__31841\,
            in1 => \N__31864\,
            in2 => \N__31785\,
            in3 => \N__57853\,
            lcout => \Commands_frame_decoder.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__56384\,
            in1 => \N__56016\,
            in2 => \N__29199\,
            in3 => \N__55835\,
            lcout => \Commands_frame_decoder.state_ns_0_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIEAGS_4_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__30249\,
            in1 => \N__29973\,
            in2 => \_gnd_net_\,
            in3 => \N__57852\,
            lcout => \uart_pc.state_RNIEAGSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55445\,
            in2 => \_gnd_net_\,
            in3 => \N__55845\,
            lcout => \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIHL1J_5_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29574\,
            in2 => \_gnd_net_\,
            in3 => \N__31762\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIE28S_5_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29436\,
            in3 => \N__57864\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__29410\,
            in1 => \N__31767\,
            in2 => \N__29387\,
            in3 => \N__53349\,
            lcout => xy_kp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59172\,
            ce => 'H',
            sr => \N__57509\
        );

    \Commands_frame_decoder.state_7_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__31766\,
            in1 => \N__29383\,
            in2 => \N__29549\,
            in3 => \N__31306\,
            lcout => \Commands_frame_decoder.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59172\,
            ce => 'H',
            sr => \N__57509\
        );

    \Commands_frame_decoder.state_RNIG48S_7_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__29379\,
            in1 => \N__31764\,
            in2 => \_gnd_net_\,
            in3 => \N__57862\,
            lcout => \Commands_frame_decoder.state_RNIG48SZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNII68S_9_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__57863\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29363\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_10_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__31765\,
            in1 => \N__29364\,
            in2 => \N__29347\,
            in3 => \N__31305\,
            lcout => \Commands_frame_decoder.stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59172\,
            ce => 'H',
            sr => \N__57509\
        );

    \Commands_frame_decoder.source_alt_kp_4_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31780\,
            in1 => \N__29306\,
            in2 => \N__29547\,
            in3 => \N__53350\,
            lcout => alt_kp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59185\,
            ce => 'H',
            sr => \N__57513\
        );

    \Commands_frame_decoder.state_RNIGK1J_4_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29513\,
            in2 => \_gnd_net_\,
            in3 => \N__31779\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_5_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__31308\,
            in1 => \N__29573\,
            in2 => \N__29577\,
            in3 => \N__31782\,
            lcout => \Commands_frame_decoder.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59185\,
            ce => 'H',
            sr => \N__57513\
        );

    \Commands_frame_decoder.state_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__31309\,
            in1 => \N__29559\,
            in2 => \N__29548\,
            in3 => \N__31783\,
            lcout => \Commands_frame_decoder.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59185\,
            ce => 'H',
            sr => \N__57513\
        );

    \Commands_frame_decoder.state_4_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__29514\,
            in1 => \N__31781\,
            in2 => \N__47946\,
            in3 => \N__31307\,
            lcout => \Commands_frame_decoder.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59185\,
            ce => 'H',
            sr => \N__57513\
        );

    \Commands_frame_decoder.state_RNID18S_4_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29502\,
            in2 => \_gnd_net_\,
            in3 => \N__57846\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_2_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29496\,
            lcout => \pid_front.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59213\,
            ce => \N__58507\,
            sr => \N__58206\
        );

    \pid_front.error_p_reg_esr_0_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29487\,
            lcout => \pid_front.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59213\,
            ce => \N__58507\,
            sr => \N__58206\
        );

    \pid_front.error_p_reg_esr_5_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29475\,
            lcout => \pid_front.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59213\,
            ce => \N__58507\,
            sr => \N__58206\
        );

    \pid_front.error_p_reg_esr_11_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29460\,
            lcout => \pid_front.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59213\,
            ce => \N__58507\,
            sr => \N__58206\
        );

    \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52679\,
            lcout => \dron_frame_decoder_1.drone_altitude_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59229\,
            ce => \N__30854\,
            sr => \N__57526\
        );

    \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52361\,
            lcout => drone_altitude_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59229\,
            ce => \N__30854\,
            sr => \N__57526\
        );

    \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50767\,
            lcout => \dron_frame_decoder_1.drone_altitude_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59229\,
            ce => \N__30854\,
            sr => \N__57526\
        );

    \dron_frame_decoder_1.state_7_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__32142\,
            in1 => \N__32170\,
            in2 => \_gnd_net_\,
            in3 => \N__34698\,
            lcout => \dron_frame_decoder_1.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59246\,
            ce => 'H',
            sr => \N__57533\
        );

    \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35810\,
            in2 => \_gnd_net_\,
            in3 => \N__35787\,
            lcout => \scaler_4.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30642\,
            lcout => drone_altitude_i_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30903\,
            lcout => drone_altitude_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30897\,
            lcout => drone_altitude_i_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29613\,
            lcout => drone_altitude_i_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30885\,
            lcout => drone_altitude_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30891\,
            lcout => drone_altitude_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_inv_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__42299\,
            in1 => \N__30655\,
            in2 => \_gnd_net_\,
            in3 => \N__29738\,
            lcout => \pid_alt.drone_altitude_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_13_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30873\,
            lcout => \pid_alt.error_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_14_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30879\,
            lcout => \pid_alt.error_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_12_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30867\,
            lcout => \pid_alt.error_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIM6G7_9_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30825\,
            in2 => \_gnd_net_\,
            in3 => \N__30787\,
            lcout => \pid_front.error_p_reg_esr_RNIM6G7Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_0__0__0_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29697\,
            lcout => \uart_drone_sync.aux_0__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_3__0__0_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29679\,
            lcout => \uart_drone_sync.aux_3__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_1__0__0_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29691\,
            lcout => \uart_drone_sync.aux_1__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_2__0__0_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29685\,
            lcout => \uart_drone_sync.aux_2__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29799\,
            in2 => \N__31164\,
            in3 => \N__31163\,
            lcout => \Commands_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_0\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29793\,
            in2 => \_gnd_net_\,
            in3 => \N__29787\,
            lcout => \Commands_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_0\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_1\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_2_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29784\,
            in2 => \_gnd_net_\,
            in3 => \N__29778\,
            lcout => \Commands_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_1\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_2\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29775\,
            in2 => \_gnd_net_\,
            in3 => \N__29769\,
            lcout => \Commands_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_2\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_3\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_4_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31053\,
            in2 => \_gnd_net_\,
            in3 => \N__29766\,
            lcout => \Commands_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_3\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_4\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_5_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31080\,
            in2 => \_gnd_net_\,
            in3 => \N__29763\,
            lcout => \Commands_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_4\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_5\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_6_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31104\,
            in2 => \_gnd_net_\,
            in3 => \N__29760\,
            lcout => \Commands_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_5\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_6\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_7_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31131\,
            in2 => \_gnd_net_\,
            in3 => \N__29757\,
            lcout => \Commands_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_6\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_7\,
            clk => \N__59086\,
            ce => 'H',
            sr => \N__29823\
        );

    \Commands_frame_decoder.WDT_8_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31092\,
            in2 => \_gnd_net_\,
            in3 => \N__29847\,
            lcout => \Commands_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_8\,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \Commands_frame_decoder.WDT_9_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31067\,
            in2 => \_gnd_net_\,
            in3 => \N__29844\,
            lcout => \Commands_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_8\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_9\,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \Commands_frame_decoder.WDT_10_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31407\,
            in2 => \_gnd_net_\,
            in3 => \N__29841\,
            lcout => \Commands_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_9\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_10\,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \Commands_frame_decoder.WDT_11_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31118\,
            in2 => \_gnd_net_\,
            in3 => \N__29838\,
            lcout => \Commands_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_10\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_11\,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \Commands_frame_decoder.WDT_12_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31419\,
            in2 => \_gnd_net_\,
            in3 => \N__29835\,
            lcout => \Commands_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_11\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_12\,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \Commands_frame_decoder.WDT_13_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31335\,
            in2 => \_gnd_net_\,
            in3 => \N__29832\,
            lcout => \Commands_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_12\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_13\,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \Commands_frame_decoder.WDT_14_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31359\,
            in2 => \_gnd_net_\,
            in3 => \N__29829\,
            lcout => \Commands_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_13\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_14\,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \Commands_frame_decoder.WDT_15_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31377\,
            in2 => \_gnd_net_\,
            in3 => \N__29826\,
            lcout => \Commands_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59092\,
            ce => 'H',
            sr => \N__29819\
        );

    \uart_pc.state_RNO_0_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__30144\,
            in1 => \N__30327\,
            in2 => \N__30045\,
            in3 => \N__57878\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__29936\,
            in1 => \N__30043\,
            in2 => \N__29802\,
            in3 => \N__29883\,
            lcout => \uart_pc.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__30044\,
            in1 => \N__30329\,
            in2 => \N__30015\,
            in3 => \N__57879\,
            lcout => \uart_pc.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_3__0__0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_3_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__31509\,
            in1 => \N__31484\,
            in2 => \N__57901\,
            in3 => \N__32500\,
            lcout => \uart_drone.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__30328\,
            in1 => \N__57871\,
            in2 => \_gnd_net_\,
            in3 => \N__30011\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001111"
        )
    port map (
            in0 => \N__29972\,
            in1 => \N__30030\,
            in2 => \N__30018\,
            in3 => \N__29935\,
            lcout => \uart_pc.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIGRIF1_2_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111100"
        )
    port map (
            in0 => \N__29934\,
            in1 => \N__30238\,
            in2 => \N__30148\,
            in3 => \N__29882\,
            lcout => \uart_pc.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIITIF1_4_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100010001"
        )
    port map (
            in0 => \N__30233\,
            in1 => \N__29968\,
            in2 => \N__29932\,
            in3 => \N__29879\,
            lcout => \uart_pc.un1_state_4_0\,
            ltout => \uart_pc.un1_state_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIUPE73_3_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30234\,
            in2 => \N__29940\,
            in3 => \N__30619\,
            lcout => \uart_pc.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_3_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__30235\,
            in1 => \N__30149\,
            in2 => \N__29933\,
            in3 => \N__29880\,
            lcout => OPEN,
            ltout => \uart_pc.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__30159\,
            in1 => \N__44950\,
            in2 => \N__30153\,
            in3 => \N__30150\,
            lcout => \uart_pc.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.Q_0__0_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30117\,
            lcout => \debug_CH2_18A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31543\,
            in2 => \_gnd_net_\,
            in3 => \N__31557\,
            lcout => OPEN,
            ltout => \uart_drone.timer_Count_RNO_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__31482\,
            in1 => \N__57883\,
            in2 => \N__30111\,
            in3 => \N__32504\,
            lcout => \uart_drone.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__57884\,
            in1 => \N__31544\,
            in2 => \N__32505\,
            in3 => \N__31481\,
            lcout => \uart_drone.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__30591\,
            in1 => \N__30333\,
            in2 => \N__30107\,
            in3 => \N__30378\,
            lcout => \uart_pc.data_AuxZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.data_Aux_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__30374\,
            in1 => \N__30582\,
            in2 => \N__30090\,
            in3 => \N__30338\,
            lcout => \uart_pc.data_AuxZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.data_Aux_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__30573\,
            in1 => \N__30334\,
            in2 => \N__30075\,
            in3 => \N__30379\,
            lcout => \uart_pc.data_AuxZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.data_Aux_3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__30375\,
            in1 => \N__30056\,
            in2 => \N__30441\,
            in3 => \N__30339\,
            lcout => \uart_pc.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.data_Aux_4_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__30168\,
            in1 => \N__30335\,
            in2 => \N__30429\,
            in3 => \N__30380\,
            lcout => \uart_pc.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.data_Aux_5_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__30376\,
            in1 => \N__30407\,
            in2 => \N__30636\,
            in3 => \N__30340\,
            lcout => \uart_pc.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.data_Aux_6_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__30627\,
            in1 => \N__30336\,
            in2 => \N__30396\,
            in3 => \N__30381\,
            lcout => \uart_pc.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.data_Aux_7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__30377\,
            in1 => \N__30337\,
            in2 => \N__30279\,
            in3 => \N__30621\,
            lcout => \uart_pc.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59117\,
            ce => 'H',
            sr => \N__30264\
        );

    \uart_pc.bit_Count_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000101100"
        )
    port map (
            in0 => \N__30248\,
            in1 => \N__30527\,
            in2 => \N__30198\,
            in3 => \N__30618\,
            lcout => \uart_pc.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59130\,
            ce => 'H',
            sr => \N__57505\
        );

    \uart_pc.bit_Count_RNO_0_2_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__30526\,
            in1 => \N__30193\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \uart_pc.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__30180\,
            in1 => \N__30564\,
            in2 => \N__30201\,
            in3 => \N__30485\,
            lcout => \uart_pc.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59130\,
            ce => 'H',
            sr => \N__57505\
        );

    \uart_pc.bit_Count_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__30528\,
            in1 => \N__30197\,
            in2 => \N__30489\,
            in3 => \N__30179\,
            lcout => \uart_pc.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59130\,
            ce => 'H',
            sr => \N__57505\
        );

    \uart_pc.data_Aux_RNO_0_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__30561\,
            in1 => \N__30477\,
            in2 => \_gnd_net_\,
            in3 => \N__30523\,
            lcout => \uart_pc.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_5_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__30524\,
            in1 => \_gnd_net_\,
            in2 => \N__30488\,
            in3 => \N__30563\,
            lcout => \uart_pc.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_6_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30562\,
            in1 => \N__30481\,
            in2 => \_gnd_net_\,
            in3 => \N__30525\,
            lcout => \uart_pc.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_5_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41258\,
            in1 => \N__41197\,
            in2 => \_gnd_net_\,
            in3 => \N__41174\,
            lcout => scaler_4_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59144\,
            ce => \N__37453\,
            sr => \N__57510\
        );

    \uart_drone.data_Aux_RNO_0_5_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__35577\,
            in1 => \N__35502\,
            in2 => \N__35430\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNI4U6E1_2_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30556\,
            in1 => \N__30518\,
            in2 => \_gnd_net_\,
            in3 => \N__30468\,
            lcout => \uart_pc.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__30519\,
            in1 => \_gnd_net_\,
            in2 => \N__30486\,
            in3 => \N__30557\,
            lcout => \uart_pc.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30559\,
            in1 => \N__30520\,
            in2 => \_gnd_net_\,
            in3 => \N__30472\,
            lcout => \uart_pc.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_2_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__30521\,
            in1 => \_gnd_net_\,
            in2 => \N__30487\,
            in3 => \N__30558\,
            lcout => \uart_pc.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__30560\,
            in1 => \N__30522\,
            in2 => \_gnd_net_\,
            in3 => \N__30476\,
            lcout => \uart_pc.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56454\,
            lcout => \frame_decoder_OFF4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59155\,
            ce => \N__33077\,
            sr => \N__57514\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_5_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55709\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58343\,
            lcout => xy_kp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59173\,
            ce => \N__31925\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55875\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58342\,
            lcout => xy_kp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59173\,
            ce => \N__31925\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_data_valid_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__32213\,
            in1 => \N__40979\,
            in2 => \_gnd_net_\,
            in3 => \N__47661\,
            lcout => \debug_CH1_0A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59186\,
            ce => 'H',
            sr => \N__57522\
        );

    \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32148\,
            in2 => \_gnd_net_\,
            in3 => \N__57847\,
            lcout => \dron_frame_decoder_1.N_513_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.state_0_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__50480\,
            in1 => \N__50611\,
            in2 => \_gnd_net_\,
            in3 => \N__47677\,
            lcout => \pid_front.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59230\,
            ce => 'H',
            sr => \N__57539\
        );

    \dron_frame_decoder_1.source_Altitude_esr_0_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52259\,
            lcout => drone_altitude_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59247\,
            ce => \N__34946\,
            sr => \N__57549\
        );

    \dron_frame_decoder_1.source_Altitude_esr_1_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50772\,
            lcout => drone_altitude_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59247\,
            ce => \N__34946\,
            sr => \N__57549\
        );

    \dron_frame_decoder_1.source_Altitude_esr_4_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52576\,
            lcout => \dron_frame_decoder_1.drone_altitude_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59247\,
            ce => \N__34946\,
            sr => \N__57549\
        );

    \dron_frame_decoder_1.source_Altitude_esr_5_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52457\,
            lcout => \dron_frame_decoder_1.drone_altitude_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59247\,
            ce => \N__34946\,
            sr => \N__57549\
        );

    \dron_frame_decoder_1.source_Altitude_esr_6_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53204\,
            lcout => \dron_frame_decoder_1.drone_altitude_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59247\,
            ce => \N__34946\,
            sr => \N__57549\
        );

    \dron_frame_decoder_1.source_Altitude_esr_7_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52378\,
            lcout => \dron_frame_decoder_1.drone_altitude_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59247\,
            ce => \N__34946\,
            sr => \N__57549\
        );

    \dron_frame_decoder_1.source_Altitude_esr_8_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52273\,
            lcout => \dron_frame_decoder_1.drone_altitude_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59262\,
            ce => \N__30850\,
            sr => \N__57559\
        );

    \dron_frame_decoder_1.source_Altitude_esr_14_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53205\,
            lcout => drone_altitude_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59262\,
            ce => \N__30850\,
            sr => \N__57559\
        );

    \dron_frame_decoder_1.source_Altitude_esr_13_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52468\,
            lcout => drone_altitude_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59262\,
            ce => \N__30850\,
            sr => \N__57559\
        );

    \dron_frame_decoder_1.source_Altitude_esr_12_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52590\,
            lcout => drone_altitude_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59262\,
            ce => \N__30850\,
            sr => \N__57559\
        );

    \pid_front.error_d_reg_esr_RNIDQE8_9_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56773\,
            in1 => \N__30824\,
            in2 => \_gnd_net_\,
            in3 => \N__30789\,
            lcout => \pid_front.un1_pid_prereg_80_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_9_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56774\,
            lcout => \pid_front.error_d_reg_prevZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59276\,
            ce => \N__49364\,
            sr => \N__57569\
        );

    \pid_front.error_p_reg_esr_RNIM6G7_0_9_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30823\,
            in2 => \_gnd_net_\,
            in3 => \N__30788\,
            lcout => \pid_front.N_1459_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30918\,
            in2 => \_gnd_net_\,
            in3 => \N__33245\,
            lcout => \pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_7_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30948\,
            lcout => \pid_front.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59288\,
            ce => \N__58449\,
            sr => \N__58193\
        );

    \pid_front.error_p_reg_esr_RNII2G7_7_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__35128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35037\,
            lcout => OPEN,
            ltout => \pid_front.N_1451_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNINKUF_7_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100101011"
        )
    port map (
            in0 => \N__59397\,
            in1 => \N__34983\,
            in2 => \N__30930\,
            in3 => \N__35010\,
            lcout => \pid_front.error_d_reg_esr_RNINKUFZ0Z_7\,
            ltout => \pid_front.error_d_reg_esr_RNINKUFZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIJETV_7_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110011001"
        )
    port map (
            in0 => \N__35129\,
            in1 => \N__30924\,
            in2 => \N__30927\,
            in3 => \N__35038\,
            lcout => \pid_front.error_p_reg_esr_RNIJETVZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNIANE8_8_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__32267\,
            in1 => \_gnd_net_\,
            in2 => \N__32310\,
            in3 => \N__53911\,
            lcout => \pid_front.un1_pid_prereg_70_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIK4G7_8_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32305\,
            in2 => \_gnd_net_\,
            in3 => \N__32266\,
            lcout => \pid_front.N_1455_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI42GP4_13_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__30961\,
            in1 => \N__30917\,
            in2 => \N__33246\,
            in3 => \N__31001\,
            lcout => \pid_front.error_p_reg_esr_RNI42GP4Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__30987\,
            in1 => \N__45057\,
            in2 => \_gnd_net_\,
            in3 => \N__59466\,
            lcout => \pid_front.un1_pid_prereg_23\,
            ltout => \pid_front.un1_pid_prereg_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIN47A4_12_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__33241\,
            in1 => \N__33189\,
            in2 => \N__31041\,
            in3 => \N__32379\,
            lcout => \pid_front.error_p_reg_esr_RNIN47A4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIO6FT1_12_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33188\,
            in2 => \_gnd_net_\,
            in3 => \N__32378\,
            lcout => \pid_front.error_p_reg_esr_RNIO6FT1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIBAOC2_15_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33537\,
            in2 => \_gnd_net_\,
            in3 => \N__33509\,
            lcout => \pid_front.error_p_reg_esr_RNIBAOC2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIK3C61_15_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__59360\,
            in1 => \_gnd_net_\,
            in2 => \N__31014\,
            in3 => \N__31035\,
            lcout => \pid_front.un1_pid_prereg_30\,
            ltout => \pid_front.un1_pid_prereg_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIGEGP4_14_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__30963\,
            in1 => \N__33536\,
            in2 => \N__31038\,
            in3 => \N__31002\,
            lcout => \pid_front.error_p_reg_esr_RNIGEGP4Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_15_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__59361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59308\,
            ce => \N__49358\,
            sr => \N__57594\
        );

    \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31034\,
            in1 => \N__31010\,
            in2 => \_gnd_net_\,
            in3 => \N__59359\,
            lcout => \pid_front.un1_pid_prereg_29\,
            ltout => \pid_front.un1_pid_prereg_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI54OC2_14_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30990\,
            in3 => \N__30962\,
            lcout => \pid_front.error_p_reg_esr_RNI54OC2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIH0C61_14_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__30986\,
            in1 => \N__45056\,
            in2 => \_gnd_net_\,
            in3 => \N__59459\,
            lcout => \pid_front.un1_pid_prereg_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.state_RNIPKTD_0_LC_8_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50493\,
            in2 => \_gnd_net_\,
            in3 => \N__57833\,
            lcout => \pid_front.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_0__0__0_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31191\,
            lcout => \uart_pc_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_1__0__0_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31185\,
            lcout => \uart_pc_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.Q_0__0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31176\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \debug_CH0_16A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNI1NQ51_15_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__31375\,
            in1 => \N__31356\,
            in2 => \_gnd_net_\,
            in3 => \N__31333\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_RNIGA2K5_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__31357\,
            in1 => \N__31435\,
            in2 => \N__31167\,
            in3 => \N__31383\,
            lcout => \Commands_frame_decoder.state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_2__0__0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31149\,
            lcout => \uart_pc_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNI8EBE1_6_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__31405\,
            in1 => \N__31130\,
            in2 => \N__31119\,
            in3 => \N__31103\,
            lcout => \Commands_frame_decoder.WDT8lto15_N_5L7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNII19A1_4_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31091\,
            in1 => \N__31079\,
            in2 => \N__31068\,
            in3 => \N__31052\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIAERH3_12_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011111111"
        )
    port map (
            in0 => \N__31418\,
            in1 => \N__31406\,
            in2 => \N__31392\,
            in3 => \N__31389\,
            lcout => \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12\,
            ltout => \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIB5MN4_15_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__31376\,
            in1 => \N__31358\,
            in2 => \N__31338\,
            in3 => \N__31334\,
            lcout => \Commands_frame_decoder.WDT8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31775\,
            in2 => \_gnd_net_\,
            in3 => \N__31436\,
            lcout => \Commands_frame_decoder.preinitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59087\,
            ce => 'H',
            sr => \N__57499\
        );

    \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33825\,
            in2 => \_gnd_net_\,
            in3 => \N__31457\,
            lcout => \uart_drone.N_126_li\,
            ltout => \uart_drone.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIAT1D1_4_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__33788\,
            in1 => \N__32606\,
            in2 => \N__31209\,
            in3 => \N__57856\,
            lcout => \uart_drone.N_143\,
            ltout => \uart_drone.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_4_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__33741\,
            in1 => \N__33930\,
            in2 => \N__31206\,
            in3 => \N__44928\,
            lcout => \uart_drone.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI9ADK1_4_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__32624\,
            in1 => \N__33928\,
            in2 => \N__31524\,
            in3 => \N__32607\,
            lcout => \uart_drone.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_4_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__57857\,
            in1 => \N__31497\,
            in2 => \N__32490\,
            in3 => \N__31485\,
            lcout => \uart_drone.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIOU0N_4_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__33929\,
            in1 => \N__32608\,
            in2 => \_gnd_net_\,
            in3 => \N__57855\,
            lcout => \uart_drone.state_RNIOU0NZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI5A9J_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__31539\,
            in1 => \N__31556\,
            in2 => \N__31545\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \uart_drone.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31458\,
            in3 => \N__31512\,
            lcout => \uart_drone.timer_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_1\,
            carryout => \uart_drone.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33836\,
            in3 => \N__31503\,
            lcout => \uart_drone.timer_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_2\,
            carryout => \uart_drone.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_4_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33776\,
            in2 => \_gnd_net_\,
            in3 => \N__31500\,
            lcout => \uart_drone.timer_Count_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_2_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__31491\,
            in1 => \N__31483\,
            in2 => \N__57903\,
            in3 => \N__32491\,
            lcout => \uart_drone.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59101\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIDGR31_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__33821\,
            in1 => \N__31453\,
            in2 => \N__33789\,
            in3 => \N__32602\,
            lcout => \uart_drone.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_rdy_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32897\,
            in2 => \_gnd_net_\,
            in3 => \N__31885\,
            lcout => uart_drone_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59110\,
            ce => 'H',
            sr => \N__57506\
        );

    \Commands_frame_decoder.source_data_valid_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__31818\,
            in1 => \N__31776\,
            in2 => \N__41009\,
            in3 => \N__31440\,
            lcout => \debug_CH3_20A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59110\,
            ce => 'H',
            sr => \N__57506\
        );

    \uart_drone.timer_Count_RNIES9Q1_2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__32864\,
            in1 => \N__31886\,
            in2 => \_gnd_net_\,
            in3 => \N__57859\,
            lcout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\,
            ltout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIRC5U2_2_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__31887\,
            in1 => \_gnd_net_\,
            in2 => \N__31869\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.data_rdyc_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31865\,
            in2 => \_gnd_net_\,
            in3 => \N__31845\,
            lcout => \Commands_frame_decoder.count_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_esr_3_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32643\,
            lcout => uart_drone_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59131\,
            ce => \N__32997\,
            sr => \N__32985\
        );

    \Commands_frame_decoder.state_RNITUI31_13_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__31812\,
            in1 => \N__31784\,
            in2 => \_gnd_net_\,
            in3 => \N__57832\,
            lcout => \Commands_frame_decoder.state_RNITUI31Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40943\,
            lcout => \dron_frame_decoder_1.N_224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__34678\,
            in1 => \N__32945\,
            in2 => \N__31569\,
            in3 => \N__31578\,
            lcout => \dron_frame_decoder_1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59156\,
            ce => 'H',
            sr => \N__57523\
        );

    \dron_frame_decoder_1.state_ns_0_a3_0_1_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53184\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52541\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_a3_0_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52649\,
            in1 => \N__31909\,
            in2 => \N__31581\,
            in3 => \N__50749\,
            lcout => \dron_frame_decoder_1.N_220\,
            ltout => \dron_frame_decoder_1.N_220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__33060\,
            in1 => \N__31893\,
            in2 => \N__31572\,
            in3 => \N__31565\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.N_198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_0_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__34679\,
            in1 => \N__32121\,
            in2 => \N__32124\,
            in3 => \N__31913\,
            lcout => \dron_frame_decoder_1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59156\,
            ce => 'H',
            sr => \N__57523\
        );

    \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__40968\,
            in1 => \N__32941\,
            in2 => \N__31914\,
            in3 => \N__32214\,
            lcout => \dron_frame_decoder_1.N_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__56466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58337\,
            lcout => xy_kp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59174\,
            ce => \N__31932\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56271\,
            lcout => xy_kp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59174\,
            ce => \N__31932\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56110\,
            in2 => \_gnd_net_\,
            in3 => \N__58339\,
            lcout => xy_kp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59174\,
            ce => \N__31932\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55342\,
            lcout => xy_kp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59174\,
            ce => \N__31932\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55548\,
            in2 => \_gnd_net_\,
            in3 => \N__58341\,
            lcout => xy_kp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59174\,
            ce => \N__31932\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_2_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__32206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31908\,
            lcout => \dron_frame_decoder_1.state_ns_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_6_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__32212\,
            in1 => \N__40980\,
            in2 => \N__32178\,
            in3 => \N__34694\,
            lcout => \dron_frame_decoder_1.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59187\,
            ce => 'H',
            sr => \N__57534\
        );

    \dron_frame_decoder_1.state_RNI0TLI1_4_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__32208\,
            in1 => \N__33144\,
            in2 => \N__57900\,
            in3 => \N__33108\,
            lcout => \dron_frame_decoder_1.N_521_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__32207\,
            in1 => \N__33107\,
            in2 => \N__32177\,
            in3 => \N__33143\,
            lcout => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33109\,
            in2 => \_gnd_net_\,
            in3 => \N__40981\,
            lcout => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4\,
            ltout => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI36DT_4_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32133\,
            in3 => \N__57850\,
            lcout => \dron_frame_decoder_1.N_505_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI4KF7_0_0_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38386\,
            in2 => \_gnd_net_\,
            in3 => \N__38352\,
            lcout => \pid_front.un1_pid_prereg_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_8_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53915\,
            lcout => \pid_front.error_d_reg_prevZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59231\,
            ce => \N__49370\,
            sr => \N__57560\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32130\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \drone_H_disp_side_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50768\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59248\,
            ce => \N__53117\,
            sr => \N__57570\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50384\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59248\,
            ce => \N__53117\,
            sr => \N__57570\
        );

    \pid_alt.error_axb_1_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32325\,
            lcout => \pid_alt.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNITOTV_8_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101001011"
        )
    port map (
            in0 => \N__32309\,
            in1 => \N__32262\,
            in2 => \N__32235\,
            in3 => \N__36488\,
            lcout => \pid_front.error_p_reg_esr_RNITOTVZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNISPUF_8_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__32226\,
            in1 => \N__35039\,
            in2 => \N__53916\,
            in3 => \N__35130\,
            lcout => \pid_front.error_d_reg_esr_RNISPUFZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI57KP4_18_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__32403\,
            in1 => \N__32421\,
            in2 => \N__42636\,
            in3 => \N__33293\,
            lcout => \pid_front.error_p_reg_esr_RNI57KP4Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIO6FT1_0_12_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33182\,
            in2 => \_gnd_net_\,
            in3 => \N__32377\,
            lcout => \pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__33968\,
            in1 => \N__46850\,
            in2 => \_gnd_net_\,
            in3 => \N__56815\,
            lcout => \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11\,
            ltout => \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNIBO6A4_12_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010110010"
        )
    port map (
            in0 => \N__53853\,
            in1 => \N__32388\,
            in2 => \N__32220\,
            in3 => \N__36983\,
            lcout => \pid_front.error_d_reg_esr_RNIBO6A4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI0GC61_19_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__32441\,
            in1 => \N__32450\,
            in2 => \_gnd_net_\,
            in3 => \N__59527\,
            lcout => \pid_front.un1_pid_prereg_57\,
            ltout => \pid_front.un1_pid_prereg_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI8ARC2_19_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32217\,
            in3 => \N__42628\,
            lcout => \pid_front.error_p_reg_esr_RNI8ARC2Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_19_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59529\,
            lcout => \pid_front.error_d_reg_prevZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59301\,
            ce => \N__49360\,
            sr => \N__57601\
        );

    \pid_front.error_p_reg_esr_RNITCC61_18_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__33276\,
            in1 => \_gnd_net_\,
            in2 => \N__49404\,
            in3 => \N__59572\,
            lcout => \pid_front.un1_pid_prereg_48\,
            ltout => \pid_front.un1_pid_prereg_48_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIKJHP4_17_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__33621\,
            in1 => \N__33609\,
            in2 => \N__32457\,
            in3 => \N__32417\,
            lcout => \pid_front.error_p_reg_esr_RNIKJHP4Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__59528\,
            in1 => \_gnd_net_\,
            in2 => \N__32454\,
            in3 => \N__32442\,
            lcout => \pid_front.un1_pid_prereg_56\,
            ltout => \pid_front.un1_pid_prereg_56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNITSOC2_18_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32406\,
            in3 => \N__32399\,
            lcout => \pid_front.error_p_reg_esr_RNITSOC2Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIA93N_0_12_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32347\,
            in2 => \_gnd_net_\,
            in3 => \N__32359\,
            lcout => \pid_front.N_1471_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_12_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53849\,
            lcout => \pid_front.error_d_reg_prevZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59309\,
            ce => \N__49359\,
            sr => \N__57609\
        );

    \pid_front.error_p_reg_esr_RNIA93N_12_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32348\,
            in2 => \_gnd_net_\,
            in3 => \N__32360\,
            lcout => \pid_front.error_p_reg_esr_RNIA93NZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIBQB61_12_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32361\,
            in1 => \N__53848\,
            in2 => \_gnd_net_\,
            in3 => \N__32349\,
            lcout => OPEN,
            ltout => \pid_front.un1_pid_prereg_107_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI1E6A4_12_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__35676\,
            in1 => \N__35661\,
            in2 => \N__32328\,
            in3 => \N__32544\,
            lcout => \pid_front.error_p_reg_esr_RNI1E6A4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_3_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__33852\,
            in1 => \N__33911\,
            in2 => \N__33797\,
            in3 => \N__32525\,
            lcout => OPEN,
            ltout => \uart_drone.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_3_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__32526\,
            in1 => \N__33734\,
            in2 => \N__32535\,
            in3 => \N__44966\,
            lcout => \uart_drone.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59078\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI62411_4_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000101"
        )
    port map (
            in0 => \N__32610\,
            in1 => \N__33790\,
            in2 => \N__33919\,
            in3 => \N__33851\,
            lcout => \uart_drone.un1_state_4_0\,
            ltout => \uart_drone.un1_state_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI63LK2_3_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33910\,
            in2 => \N__32532\,
            in3 => \N__35615\,
            lcout => \uart_drone.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_2_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__32519\,
            in1 => \N__32860\,
            in2 => \N__32568\,
            in3 => \N__57876\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_2_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__32567\,
            in1 => \N__33787\,
            in2 => \N__32529\,
            in3 => \N__33859\,
            lcout => \uart_drone.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI40411_2_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101010"
        )
    port map (
            in0 => \N__33912\,
            in1 => \N__33785\,
            in2 => \N__33861\,
            in3 => \N__32518\,
            lcout => \uart_drone.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNO_0_2_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33874\,
            in2 => \_gnd_net_\,
            in3 => \N__35407\,
            lcout => \uart_drone.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_0_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__57875\,
            in1 => \N__32576\,
            in2 => \_gnd_net_\,
            in3 => \N__32859\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_0_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__33786\,
            in1 => \N__32625\,
            in2 => \N__32613\,
            in3 => \N__32609\,
            lcout => \uart_drone.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_1_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__57877\,
            in1 => \N__32566\,
            in2 => \N__32888\,
            in3 => \N__32577\,
            lcout => \uart_drone.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__32688\,
            in1 => \N__32676\,
            in2 => \N__34266\,
            in3 => \N__33669\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_6_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__35538\,
            in1 => \N__35465\,
            in2 => \_gnd_net_\,
            in3 => \N__35406\,
            lcout => \uart_drone.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34022\,
            in1 => \N__34037\,
            in2 => \N__34008\,
            in3 => \N__34067\,
            lcout => \reset_module_System.reset6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__34053\,
            in1 => \N__33660\,
            in2 => \N__34092\,
            in3 => \N__33681\,
            lcout => \reset_module_System.reset6_15\,
            ltout => \reset_module_System.reset6_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__33704\,
            in1 => \N__34261\,
            in2 => \N__32550\,
            in3 => \N__32686\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33703\,
            in2 => \_gnd_net_\,
            in3 => \N__33723\,
            lcout => OPEN,
            ltout => \reset_module_System.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__32675\,
            in1 => \N__34262\,
            in2 => \N__32547\,
            in3 => \N__32687\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35486\,
            in1 => \N__35560\,
            in2 => \_gnd_net_\,
            in3 => \N__35421\,
            lcout => \uart_drone.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIR9N6_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33644\,
            in2 => \_gnd_net_\,
            in3 => \N__33721\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIA72I1_16_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__34109\,
            in1 => \N__34127\,
            in2 => \N__32700\,
            in3 => \N__32697\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIMJ304_12_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__33984\,
            in1 => \N__33702\,
            in2 => \N__32691\,
            in3 => \N__34194\,
            lcout => \reset_module_System.reset6_19\,
            ltout => \reset_module_System.reset6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32674\,
            in2 => \N__32661\,
            in3 => \N__34250\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_2_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__35420\,
            in1 => \_gnd_net_\,
            in2 => \N__35572\,
            in3 => \N__35487\,
            lcout => \uart_drone.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__32658\,
            in1 => \N__32889\,
            in2 => \N__32778\,
            in3 => \N__32820\,
            lcout => \uart_drone.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_Aux_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__32894\,
            in1 => \N__34320\,
            in2 => \N__32763\,
            in3 => \N__32816\,
            lcout => \uart_drone.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_Aux_2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__32652\,
            in1 => \N__32890\,
            in2 => \N__32748\,
            in3 => \N__32821\,
            lcout => \uart_drone.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_Aux_3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__32895\,
            in1 => \N__35349\,
            in2 => \N__32642\,
            in3 => \N__32817\,
            lcout => \uart_drone.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_Aux_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__32964\,
            in1 => \N__32891\,
            in2 => \N__32718\,
            in3 => \N__32822\,
            lcout => \uart_drone.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_Aux_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__32896\,
            in1 => \N__32925\,
            in2 => \N__32733\,
            in3 => \N__32818\,
            lcout => \uart_drone.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_Aux_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__32913\,
            in1 => \N__32892\,
            in2 => \N__33027\,
            in3 => \N__32823\,
            lcout => \uart_drone.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_Aux_7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__32893\,
            in1 => \N__32819\,
            in2 => \N__33012\,
            in3 => \N__35616\,
            lcout => \uart_drone.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59095\,
            ce => 'H',
            sr => \N__32790\
        );

    \uart_drone.data_esr_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32777\,
            lcout => uart_drone_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59103\,
            ce => \N__32996\,
            sr => \N__32981\
        );

    \uart_drone.data_esr_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32762\,
            lcout => uart_drone_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59103\,
            ce => \N__32996\,
            sr => \N__32981\
        );

    \uart_drone.data_esr_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32747\,
            lcout => uart_drone_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59103\,
            ce => \N__32996\,
            sr => \N__32981\
        );

    \uart_drone.data_esr_5_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32732\,
            lcout => uart_drone_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59103\,
            ce => \N__32996\,
            sr => \N__32981\
        );

    \uart_drone.data_esr_4_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32714\,
            lcout => uart_drone_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59103\,
            ce => \N__32996\,
            sr => \N__32981\
        );

    \uart_drone.data_esr_6_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33026\,
            lcout => uart_drone_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59103\,
            ce => \N__32996\,
            sr => \N__32981\
        );

    \uart_drone.data_esr_7_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33011\,
            lcout => uart_drone_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59103\,
            ce => \N__32996\,
            sr => \N__32981\
        );

    \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010011"
        )
    port map (
            in0 => \N__34464\,
            in1 => \N__40944\,
            in2 => \N__34560\,
            in3 => \N__34580\,
            lcout => \dron_frame_decoder_1.N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__34579\,
            in1 => \N__34555\,
            in2 => \_gnd_net_\,
            in3 => \N__34463\,
            lcout => \dron_frame_decoder_1.WDT10_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_4_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__35422\,
            in1 => \N__35576\,
            in2 => \_gnd_net_\,
            in3 => \N__35498\,
            lcout => \uart_drone.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52426\,
            in1 => \N__52247\,
            in2 => \N__52347\,
            in3 => \N__50336\,
            lcout => \dron_frame_decoder_1.N_263_5\,
            ltout => \dron_frame_decoder_1.N_263_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_3_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40945\,
            in2 => \N__32949\,
            in3 => \N__32946\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_ctle_14_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41008\,
            in2 => \_gnd_net_\,
            in3 => \N__57849\,
            lcout => \scaler_4.debug_CH3_20A_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset4data_esr_2_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59119\,
            ce => \N__33081\,
            sr => \N__57518\
        );

    \Commands_frame_decoder.source_offset4data_esr_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56270\,
            lcout => \frame_decoder_OFF4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59119\,
            ce => \N__33081\,
            sr => \N__57518\
        );

    \Commands_frame_decoder.source_offset4data_esr_6_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55730\,
            lcout => \frame_decoder_OFF4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59119\,
            ce => \N__33081\,
            sr => \N__57518\
        );

    \Commands_frame_decoder.source_offset4data_esr_3_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__55343\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59119\,
            ce => \N__33081\,
            sr => \N__57518\
        );

    \Commands_frame_decoder.source_offset4data_esr_4_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53370\,
            lcout => \frame_decoder_OFF4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59119\,
            ce => \N__33081\,
            sr => \N__57518\
        );

    \Commands_frame_decoder.source_offset4data_esr_5_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55898\,
            lcout => \frame_decoder_OFF4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59119\,
            ce => \N__33081\,
            sr => \N__57518\
        );

    \Commands_frame_decoder.source_offset4data_ess_7_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55541\,
            lcout => \frame_decoder_OFF4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59119\,
            ce => \N__33081\,
            sr => \N__57518\
        );

    \dron_frame_decoder_1.state_ns_i_a2_0_4_0_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50731\,
            in1 => \N__53185\,
            in2 => \N__52663\,
            in3 => \N__52542\,
            lcout => \dron_frame_decoder_1.N_219_4\,
            ltout => \dron_frame_decoder_1.N_219_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_3_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__34366\,
            in1 => \N__34677\,
            in2 => \N__33051\,
            in3 => \N__33048\,
            lcout => \dron_frame_decoder_1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59132\,
            ce => 'H',
            sr => \N__57524\
        );

    \ppm_encoder_1.rudder_esr_5_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33039\,
            lcout => \ppm_encoder_1.rudderZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59146\,
            ce => \N__46763\,
            sr => \N__57527\
        );

    \pid_front.error_p_reg_esr_1_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33153\,
            lcout => \pid_front.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59158\,
            ce => \N__58503\,
            sr => \N__58197\
        );

    \dron_frame_decoder_1.state_RNI7Q6K_5_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40964\,
            in2 => \_gnd_net_\,
            in3 => \N__33129\,
            lcout => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_5_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__34693\,
            in1 => \_gnd_net_\,
            in2 => \N__33135\,
            in3 => \N__36174\,
            lcout => \dron_frame_decoder_1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59175\,
            ce => 'H',
            sr => \N__57540\
        );

    \dron_frame_decoder_1.state_4_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__40970\,
            in1 => \N__33131\,
            in2 => \N__33117\,
            in3 => \N__34692\,
            lcout => \dron_frame_decoder_1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59175\,
            ce => 'H',
            sr => \N__57540\
        );

    \dron_frame_decoder_1.state_RNI1H181_5_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__40969\,
            in1 => \N__33130\,
            in2 => \N__33116\,
            in3 => \N__57848\,
            lcout => \dron_frame_decoder_1.N_497_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_16_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56727\,
            lcout => \pid_front.error_d_reg_prevZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59189\,
            ce => \N__49371\,
            sr => \N__57550\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33087\,
            lcout => \drone_H_disp_side_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_10_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__50605\,
            in1 => \N__35271\,
            in2 => \N__37915\,
            in3 => \N__36378\,
            lcout => front_order_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59214\,
            ce => 'H',
            sr => \N__35189\
        );

    \pid_front.source_pid_1_11_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__35272\,
            in1 => \N__50608\,
            in2 => \N__37873\,
            in3 => \N__37062\,
            lcout => front_order_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59214\,
            ce => 'H',
            sr => \N__35189\
        );

    \pid_front.source_pid_1_6_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__50606\,
            in1 => \N__35273\,
            in2 => \N__37681\,
            in3 => \N__36633\,
            lcout => front_order_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59214\,
            ce => 'H',
            sr => \N__35189\
        );

    \pid_front.source_pid_1_7_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__35274\,
            in1 => \N__50609\,
            in2 => \N__40291\,
            in3 => \N__36585\,
            lcout => front_order_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59214\,
            ce => 'H',
            sr => \N__35189\
        );

    \pid_front.source_pid_1_8_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__50607\,
            in1 => \N__35275\,
            in2 => \N__37993\,
            in3 => \N__36525\,
            lcout => front_order_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59214\,
            ce => 'H',
            sr => \N__35189\
        );

    \pid_front.source_pid_1_9_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__35276\,
            in1 => \N__50610\,
            in2 => \N__37954\,
            in3 => \N__36459\,
            lcout => front_order_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59214\,
            ce => 'H',
            sr => \N__35189\
        );

    \pid_front.pid_prereg_esr_RNI6DCJ3_13_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111010"
        )
    port map (
            in0 => \N__37141\,
            in1 => \_gnd_net_\,
            in2 => \N__35331\,
            in3 => \N__36956\,
            lcout => \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13\,
            ltout => \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNICUKFA_6_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35085\,
            in1 => \N__35076\,
            in2 => \N__33171\,
            in3 => \N__33630\,
            lcout => OPEN,
            ltout => \pid_front.pid_prereg_esr_RNICUKFAZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIC8N8C_5_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33441\,
            in2 => \N__33168\,
            in3 => \N__33162\,
            lcout => \pid_front.un1_reset_0_i\,
            ltout => \pid_front.un1_reset_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.state_RNI9HEDC_1_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__50624\,
            in1 => \_gnd_net_\,
            in2 => \N__33165\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIKVDO_23_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__37142\,
            in1 => \N__50622\,
            in2 => \_gnd_net_\,
            in3 => \N__57831\,
            lcout => \pid_front.un1_reset_0_i_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNI86GE_2_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36336\,
            in1 => \N__49427\,
            in2 => \N__36780\,
            in3 => \N__50441\,
            lcout => OPEN,
            ltout => \pid_front.m32_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNICAK01_5_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__36678\,
            in1 => \N__50623\,
            in2 => \N__33156\,
            in3 => \N__44984\,
            lcout => \pid_front.un1_reset_0_i_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_5_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__33356\,
            in1 => \N__39675\,
            in2 => \N__33435\,
            in3 => \N__33402\,
            lcout => \pid_alt.error_i_acummZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59249\,
            ce => 'H',
            sr => \N__33342\
        );

    \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33581\,
            in1 => \N__33554\,
            in2 => \_gnd_net_\,
            in3 => \N__56723\,
            lcout => \pid_front.un1_pid_prereg_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIOUOP4_19_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42562\,
            in1 => \N__42635\,
            in2 => \N__33300\,
            in3 => \N__42634\,
            lcout => \pid_front.error_p_reg_esr_RNIOUOP4Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI09RP4_20_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__42566\,
            in1 => \N__42633\,
            in2 => \N__42567\,
            in3 => \N__42632\,
            lcout => \pid_front.error_p_reg_esr_RNI09RP4Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33272\,
            in1 => \N__49400\,
            in2 => \_gnd_net_\,
            in3 => \N__59574\,
            lcout => \pid_front.un1_pid_prereg_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIETB61_13_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__33219\,
            in1 => \N__56849\,
            in2 => \_gnd_net_\,
            in3 => \N__33198\,
            lcout => \pid_front.un1_pid_prereg_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_13_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56850\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59264\,
            ce => \N__49363\,
            sr => \N__57595\
        );

    \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33218\,
            in1 => \N__56848\,
            in2 => \_gnd_net_\,
            in3 => \N__33197\,
            lcout => \pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNI6FQ75_23_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__37140\,
            in1 => \N__36732\,
            in2 => \N__35094\,
            in3 => \N__35318\,
            lcout => \pid_front.pid_prereg_esr_RNI6FQ75Z0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNINMOC2_17_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33620\,
            lcout => \pid_front.error_p_reg_esr_RNINMOC2Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__56672\,
            in1 => \_gnd_net_\,
            in2 => \N__33477\,
            in3 => \N__33498\,
            lcout => \pid_front.un1_pid_prereg_42\,
            ltout => \pid_front.un1_pid_prereg_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI87HP4_16_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__33605\,
            in1 => \N__33453\,
            in2 => \N__33585\,
            in3 => \N__33465\,
            lcout => \pid_front.error_p_reg_esr_RNI87HP4Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_17_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59277\,
            ce => \N__49361\,
            sr => \N__57602\
        );

    \pid_front.error_p_reg_esr_RNIN6C61_16_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__33582\,
            in1 => \N__33558\,
            in2 => \_gnd_net_\,
            in3 => \N__56710\,
            lcout => \pid_front.un1_pid_prereg_36\,
            ltout => \pid_front.un1_pid_prereg_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNISQGP4_15_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__33464\,
            in1 => \N__33535\,
            in2 => \N__33516\,
            in3 => \N__33513\,
            lcout => \pid_front.error_p_reg_esr_RNISQGP4Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33497\,
            in1 => \N__33473\,
            in2 => \_gnd_net_\,
            in3 => \N__56671\,
            lcout => \pid_front.un1_pid_prereg_41\,
            ltout => \pid_front.un1_pid_prereg_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIHGOC2_16_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33456\,
            in3 => \N__33452\,
            lcout => \pid_front.error_p_reg_esr_RNIHGOC2Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33969\,
            in1 => \N__46851\,
            in2 => \_gnd_net_\,
            in3 => \N__56823\,
            lcout => \pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__35483\,
            in1 => \N__35408\,
            in2 => \N__33882\,
            in3 => \N__33944\,
            lcout => \uart_drone.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59079\,
            ce => 'H',
            sr => \N__57500\
        );

    \uart_drone.bit_Count_2_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__33945\,
            in1 => \N__33936\,
            in2 => \N__35571\,
            in3 => \N__35484\,
            lcout => \uart_drone.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59079\,
            ce => 'H',
            sr => \N__57500\
        );

    \uart_drone.bit_Count_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101000000"
        )
    port map (
            in0 => \N__35608\,
            in1 => \N__33918\,
            in2 => \N__33881\,
            in3 => \N__35409\,
            lcout => \uart_drone.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59079\,
            ce => 'H',
            sr => \N__57500\
        );

    \uart_drone.timer_Count_RNIU8TV1_3_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33860\,
            in1 => \N__35607\,
            in2 => \_gnd_net_\,
            in3 => \N__33798\,
            lcout => \uart_drone.N_144_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33722\,
            in2 => \N__33705\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33680\,
            in2 => \_gnd_net_\,
            in3 => \N__33663\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33659\,
            in2 => \_gnd_net_\,
            in3 => \N__33648\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__59082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33645\,
            in2 => \_gnd_net_\,
            in3 => \N__33633\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__59082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34068\,
            in2 => \_gnd_net_\,
            in3 => \N__34056\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__59082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34052\,
            in2 => \_gnd_net_\,
            in3 => \N__34041\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__59082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34038\,
            in2 => \_gnd_net_\,
            in3 => \N__34026\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__59082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34023\,
            in2 => \_gnd_net_\,
            in3 => \N__34011\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__59082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34007\,
            in2 => \_gnd_net_\,
            in3 => \N__33993\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34286\,
            in2 => \_gnd_net_\,
            in3 => \N__33990\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34301\,
            in2 => \_gnd_net_\,
            in3 => \N__33987\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33983\,
            in2 => \_gnd_net_\,
            in3 => \N__33972\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34206\,
            in2 => \_gnd_net_\,
            in3 => \N__34137\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34313\,
            in2 => \_gnd_net_\,
            in3 => \N__34134\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34230\,
            in2 => \_gnd_net_\,
            in3 => \N__34131\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34128\,
            in2 => \_gnd_net_\,
            in3 => \N__34116\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__59085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34274\,
            in2 => \_gnd_net_\,
            in3 => \N__34113\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__59090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34110\,
            in2 => \_gnd_net_\,
            in3 => \N__34098\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__59090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34239\,
            in2 => \_gnd_net_\,
            in3 => \N__34095\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__59090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34088\,
            in2 => \_gnd_net_\,
            in3 => \N__34074\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__59090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34217\,
            in2 => \_gnd_net_\,
            in3 => \N__34071\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__35485\,
            in1 => \N__35559\,
            in2 => \_gnd_net_\,
            in3 => \N__35419\,
            lcout => \uart_drone.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNISRMR1_10_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34314\,
            in1 => \N__34302\,
            in2 => \N__34290\,
            in3 => \N__34275\,
            lcout => \reset_module_System.reset6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34238\,
            in1 => \N__34229\,
            in2 => \N__34218\,
            in3 => \N__34205\,
            lcout => \reset_module_System.reset6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34173\,
            in2 => \N__34188\,
            in3 => \N__34187\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_0\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34167\,
            in2 => \_gnd_net_\,
            in3 => \N__34161\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_0\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_1\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34158\,
            in2 => \_gnd_net_\,
            in3 => \N__34152\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_1\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_2\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34149\,
            in2 => \_gnd_net_\,
            in3 => \N__34143\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_2\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_3\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34493\,
            in2 => \_gnd_net_\,
            in3 => \N__34140\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_3\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_4\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34541\,
            in2 => \_gnd_net_\,
            in3 => \N__34347\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_4\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_5\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34508\,
            in2 => \_gnd_net_\,
            in3 => \N__34344\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_5\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_6\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34526\,
            in2 => \_gnd_net_\,
            in3 => \N__34341\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_6\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_7\,
            clk => \N__59096\,
            ce => 'H',
            sr => \N__40875\
        );

    \dron_frame_decoder_1.WDT_8_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34407\,
            in2 => \_gnd_net_\,
            in3 => \N__34338\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_8\,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_9_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34479\,
            in2 => \_gnd_net_\,
            in3 => \N__34335\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_8\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_9\,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_10_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34442\,
            in2 => \_gnd_net_\,
            in3 => \N__34332\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_9\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_10\,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_11_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34422\,
            in2 => \_gnd_net_\,
            in3 => \N__34329\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_10\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_11\,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_12_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34394\,
            in2 => \_gnd_net_\,
            in3 => \N__34326\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_11\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_12\,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_13_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34455\,
            in2 => \_gnd_net_\,
            in3 => \N__34323\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_12\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_13\,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_14_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34581\,
            in2 => \_gnd_net_\,
            in3 => \N__34566\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_13\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_14\,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_15_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34559\,
            in2 => \_gnd_net_\,
            in3 => \N__34563\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59104\,
            ce => 'H',
            sr => \N__40871\
        );

    \dron_frame_decoder_1.WDT_RNIIVJ1_4_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34542\,
            in1 => \N__34527\,
            in2 => \N__34512\,
            in3 => \N__34494\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.WDT_RNIIVJ1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIATMH2_9_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__34478\,
            in1 => \N__34428\,
            in2 => \N__34467\,
            in3 => \N__34377\,
            lcout => \dron_frame_decoder_1.WDT10lt14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__34454\,
            in1 => \N__34393\,
            in2 => \N__34443\,
            in3 => \N__34421\,
            lcout => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI2LQQ_8_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__34420\,
            in1 => \N__34406\,
            in2 => \N__34395\,
            in3 => \_gnd_net_\,
            lcout => \dron_frame_decoder_1.WDT10lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNITC181_2_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__36153\,
            in1 => \N__40974\,
            in2 => \N__34370\,
            in3 => \N__57841\,
            lcout => \dron_frame_decoder_1.N_481_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_5_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__34596\,
            in1 => \N__34632\,
            in2 => \N__45314\,
            in3 => \N__43216\,
            lcout => \ppm_encoder_1.throttleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59120\,
            ce => 'H',
            sr => \N__57528\
        );

    \dron_frame_decoder_1.state_2_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__36152\,
            in1 => \N__40983\,
            in2 => \N__34371\,
            in3 => \N__34691\,
            lcout => \dron_frame_decoder_1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59120\,
            ce => 'H',
            sr => \N__57528\
        );

    \ppm_encoder_1.un1_throttle_cry_0_c_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36248\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41435\,
            in2 => \N__42295\,
            in3 => \N__34644\,
            lcout => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_0\,
            carryout => \ppm_encoder_1.un1_throttle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37613\,
            in2 => \_gnd_net_\,
            in3 => \N__34641\,
            lcout => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_1\,
            carryout => \ppm_encoder_1.un1_throttle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36086\,
            in2 => \N__42296\,
            in3 => \N__34638\,
            lcout => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_2\,
            carryout => \ppm_encoder_1.un1_throttle_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36020\,
            in2 => \_gnd_net_\,
            in3 => \N__34635\,
            lcout => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_3\,
            carryout => \ppm_encoder_1.un1_throttle_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34631\,
            in2 => \_gnd_net_\,
            in3 => \N__34590\,
            lcout => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_4\,
            carryout => \ppm_encoder_1.un1_throttle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36125\,
            in2 => \N__42297\,
            in3 => \N__34587\,
            lcout => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_5\,
            carryout => \ppm_encoder_1.un1_throttle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36219\,
            in2 => \_gnd_net_\,
            in3 => \N__34584\,
            lcout => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_6\,
            carryout => \ppm_encoder_1.un1_throttle_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35978\,
            in2 => \_gnd_net_\,
            in3 => \N__34785\,
            lcout => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36065\,
            in2 => \_gnd_net_\,
            in3 => \N__34782\,
            lcout => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_8\,
            carryout => \ppm_encoder_1.un1_throttle_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34728\,
            in2 => \_gnd_net_\,
            in3 => \N__34779\,
            lcout => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_9\,
            carryout => \ppm_encoder_1.un1_throttle_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40046\,
            in2 => \_gnd_net_\,
            in3 => \N__34776\,
            lcout => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_10\,
            carryout => \ppm_encoder_1.un1_throttle_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35939\,
            in2 => \_gnd_net_\,
            in3 => \N__34773\,
            lcout => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_11\,
            carryout => \ppm_encoder_1.un1_throttle_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42258\,
            in2 => \N__34764\,
            in3 => \N__34770\,
            lcout => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_12\,
            carryout => \ppm_encoder_1.un1_throttle_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_14_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34767\,
            lcout => \ppm_encoder_1.throttleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59147\,
            ce => \N__46762\,
            sr => \N__57541\
        );

    \ppm_encoder_1.throttle_13_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__34760\,
            in1 => \N__34734\,
            in2 => \N__45387\,
            in3 => \N__37813\,
            lcout => \ppm_encoder_1.throttleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59159\,
            ce => 'H',
            sr => \N__57551\
        );

    \ppm_encoder_1.aileron_9_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__42849\,
            in1 => \N__34875\,
            in2 => \N__45386\,
            in3 => \N__39974\,
            lcout => \ppm_encoder_1.aileronZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59159\,
            ce => 'H',
            sr => \N__57551\
        );

    \ppm_encoder_1.throttle_10_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__34727\,
            in1 => \N__34815\,
            in2 => \N__40552\,
            in3 => \N__45321\,
            lcout => \ppm_encoder_1.throttleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59159\,
            ce => 'H',
            sr => \N__57551\
        );

    \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43293\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41547\,
            in2 => \N__42364\,
            in3 => \N__34809\,
            lcout => \ppm_encoder_1.un1_aileron_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_0\,
            carryout => \ppm_encoder_1.un1_aileron_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41124\,
            in2 => \_gnd_net_\,
            in3 => \N__34806\,
            lcout => \ppm_encoder_1.un1_aileron_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_1\,
            carryout => \ppm_encoder_1.un1_aileron_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43952\,
            in2 => \N__42365\,
            in3 => \N__34803\,
            lcout => \ppm_encoder_1.un1_aileron_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_2\,
            carryout => \ppm_encoder_1.un1_aileron_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43247\,
            in2 => \_gnd_net_\,
            in3 => \N__34800\,
            lcout => \ppm_encoder_1.un1_aileron_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_3\,
            carryout => \ppm_encoder_1.un1_aileron_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43275\,
            in2 => \_gnd_net_\,
            in3 => \N__34797\,
            lcout => \ppm_encoder_1.un1_aileron_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_4\,
            carryout => \ppm_encoder_1.un1_aileron_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42336\,
            in2 => \N__42974\,
            in3 => \N__34794\,
            lcout => \ppm_encoder_1.un1_aileron_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_5\,
            carryout => \ppm_encoder_1.un1_aileron_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42929\,
            in3 => \N__34791\,
            lcout => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_6\,
            carryout => \ppm_encoder_1.un1_aileron_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42884\,
            in2 => \_gnd_net_\,
            in3 => \N__34788\,
            lcout => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42848\,
            in2 => \_gnd_net_\,
            in3 => \N__34866\,
            lcout => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_8\,
            carryout => \ppm_encoder_1.un1_aileron_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43044\,
            in2 => \_gnd_net_\,
            in3 => \N__34863\,
            lcout => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_9\,
            carryout => \ppm_encoder_1.un1_aileron_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43011\,
            in2 => \_gnd_net_\,
            in3 => \N__34860\,
            lcout => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_10\,
            carryout => \ppm_encoder_1.un1_aileron_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45597\,
            in2 => \_gnd_net_\,
            in3 => \N__34857\,
            lcout => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_11\,
            carryout => \ppm_encoder_1.un1_aileron_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48066\,
            in2 => \N__42366\,
            in3 => \N__34854\,
            lcout => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_12\,
            carryout => \ppm_encoder_1.un1_aileron_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_14_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34851\,
            lcout => \ppm_encoder_1.aileronZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59190\,
            ce => \N__46782\,
            sr => \N__57571\
        );

    \pid_alt.error_axb_2_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34836\,
            lcout => \pid_alt.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_2_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50383\,
            lcout => drone_altitude_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59200\,
            ce => \N__34953\,
            sr => \N__57576\
        );

    \pid_alt.error_axb_3_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34959\,
            lcout => \pid_alt.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_3_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52683\,
            lcout => drone_altitude_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59200\,
            ce => \N__34953\,
            sr => \N__57576\
        );

    \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34923\,
            lcout => \pid_alt.error_d_reg_prev_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_1_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36255\,
            lcout => \pid_front.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIUJRT3_12_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__36957\,
            in1 => \N__37008\,
            in2 => \N__37146\,
            in3 => \N__35330\,
            lcout => \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12\,
            ltout => \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNI3F0N8_10_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__35297\,
            in1 => \N__35233\,
            in2 => \N__34884\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10\,
            ltout => \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_esr_1_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__50442\,
            in1 => \N__36725\,
            in2 => \N__34881\,
            in3 => \N__35065\,
            lcout => front_order_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59215\,
            ce => \N__35209\,
            sr => \N__35187\
        );

    \pid_front.source_pid_1_esr_2_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__35066\,
            in1 => \N__36726\,
            in2 => \N__36335\,
            in3 => \N__35053\,
            lcout => front_order_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59215\,
            ce => \N__35209\,
            sr => \N__35187\
        );

    \pid_front.pid_prereg_esr_RNIDT6R8_5_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__35234\,
            in1 => \N__35298\,
            in2 => \N__36686\,
            in3 => \N__35269\,
            lcout => \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5\,
            ltout => \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_esr_0_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__36724\,
            in1 => \N__49431\,
            in2 => \N__34878\,
            in3 => \N__35052\,
            lcout => front_order_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59215\,
            ce => \N__35209\,
            sr => \N__35187\
        );

    \pid_front.source_pid_1_esr_4_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__35055\,
            in1 => \N__36723\,
            in2 => \N__36687\,
            in3 => \N__35270\,
            lcout => front_order_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59215\,
            ce => \N__35209\,
            sr => \N__35187\
        );

    \pid_front.source_pid_1_esr_3_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__35067\,
            in1 => \N__36727\,
            in2 => \N__36776\,
            in3 => \N__35054\,
            lcout => front_order_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59215\,
            ce => \N__35209\,
            sr => \N__35187\
        );

    \pid_front.error_d_reg_esr_RNI7KE8_7_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35040\,
            in1 => \N__35119\,
            in2 => \_gnd_net_\,
            in3 => \N__59395\,
            lcout => OPEN,
            ltout => \pid_front.un1_pid_prereg_60_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI94TV_6_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101001011"
        )
    port map (
            in0 => \N__35009\,
            in1 => \N__34979\,
            in2 => \N__35016\,
            in3 => \N__36606\,
            lcout => \pid_front.error_p_reg_esr_RNI94TVZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_6_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52217\,
            lcout => \pid_front.error_d_reg_prevZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59232\,
            ce => \N__49366\,
            sr => \N__57596\
        );

    \pid_front.error_p_reg_esr_RNIG0G7_6_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35007\,
            in2 => \_gnd_net_\,
            in3 => \N__34977\,
            lcout => OPEN,
            ltout => \pid_front.N_1447_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNIIFUF_6_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__52218\,
            in1 => \N__38049\,
            in2 => \N__35013\,
            in3 => \N__38304\,
            lcout => \pid_front.error_d_reg_esr_RNIIFUFZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNI4HE8_6_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52216\,
            in1 => \N__35008\,
            in2 => \_gnd_net_\,
            in3 => \N__34978\,
            lcout => OPEN,
            ltout => \pid_front.un1_pid_prereg_50_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIH8R01_5_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000001111"
        )
    port map (
            in0 => \N__38013\,
            in1 => \N__38048\,
            in2 => \N__34962\,
            in3 => \N__38303\,
            lcout => \pid_front.error_p_reg_esr_RNIH8R01Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_7_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__59396\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59232\,
            ce => \N__49366\,
            sr => \N__57596\
        );

    \pid_front.pid_prereg_esr_RNII3QG_6_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36524\,
            in1 => \N__36625\,
            in2 => \N__36580\,
            in3 => \N__36451\,
            lcout => \pid_front.m26_e_5\,
            ltout => \pid_front.m26_e_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIVDO51_10_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__37055\,
            in1 => \_gnd_net_\,
            in2 => \N__35106\,
            in3 => \N__36371\,
            lcout => \pid_front.pid_prereg_esr_RNIVDO51Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIHEUK_12_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37002\,
            in2 => \_gnd_net_\,
            in3 => \N__36942\,
            lcout => OPEN,
            ltout => \pid_front.m26_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIGSMQ1_10_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37053\,
            in1 => \N__36369\,
            in2 => \N__35103\,
            in3 => \N__35100\,
            lcout => \pid_front.pid_prereg_esr_RNIGSMQ1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIEUJ31_10_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36370\,
            in1 => \N__37054\,
            in2 => \N__36731\,
            in3 => \N__37003\,
            lcout => \pid_front.m18_s_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNII3QG_0_6_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36514\,
            in1 => \N__36626\,
            in2 => \N__36581\,
            in3 => \N__36452\,
            lcout => \pid_front.m18_s_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_esr_12_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__36949\,
            in1 => \N__37004\,
            in2 => \N__37139\,
            in3 => \N__35325\,
            lcout => front_order_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59250\,
            ce => \N__35220\,
            sr => \N__35188\
        );

    \pid_front.source_pid_1_esr_13_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__35326\,
            in1 => \N__37124\,
            in2 => \_gnd_net_\,
            in3 => \N__36948\,
            lcout => front_order_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59250\,
            ce => \N__35220\,
            sr => \N__35188\
        );

    \pid_front.pid_prereg_esr_RNIMHT91_16_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36831\,
            in1 => \N__36801\,
            in2 => \N__37278\,
            in3 => \N__37245\,
            lcout => \pid_front.m9_e_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIEREV_14_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__36864\,
            in1 => \N__36900\,
            in2 => \_gnd_net_\,
            in3 => \N__37158\,
            lcout => OPEN,
            ltout => \pid_front.m9_e_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIJRCU2_20_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__37179\,
            in1 => \N__37212\,
            in2 => \N__35340\,
            in3 => \N__35337\,
            lcout => \pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_esr_5_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__35296\,
            in1 => \N__35280\,
            in2 => \N__36685\,
            in3 => \N__35241\,
            lcout => front_order_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59265\,
            ce => \N__35219\,
            sr => \N__35193\
        );

    \pid_front.state_RNIVIRQ_0_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__50625\,
            in1 => \N__47709\,
            in2 => \N__50507\,
            in3 => \N__57835\,
            lcout => OPEN,
            ltout => \pid_front.state_RNIVIRQZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.state_RNISV141_0_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35160\,
            in3 => \N__58320\,
            lcout => \pid_front.N_543_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNI9NAB3_10_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54314\,
            in1 => \N__35646\,
            in2 => \N__37082\,
            in3 => \N__35634\,
            lcout => \pid_front.error_d_reg_esr_RNI9NAB3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI653N_0_10_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35153\,
            in2 => \_gnd_net_\,
            in3 => \N__35684\,
            lcout => \pid_front.N_1463_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI653N_10_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__35685\,
            in1 => \_gnd_net_\,
            in2 => \N__35157\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_p_reg_esr_RNI653NZ0Z_10\,
            ltout => \pid_front.error_p_reg_esr_RNI653NZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIESET1_0_10_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35674\,
            in2 => \N__35133\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_10_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54315\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59278\,
            ce => \N__49362\,
            sr => \N__57616\
        );

    \pid_front.error_p_reg_esr_RNIESET1_10_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35675\,
            in2 => \_gnd_net_\,
            in3 => \N__35657\,
            lcout => \pid_front.error_p_reg_esr_RNIESET1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNISPQT1_10_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54308\,
            in1 => \N__35645\,
            in2 => \N__36420\,
            in3 => \N__35633\,
            lcout => \pid_front.error_d_reg_esr_RNISPQT1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNIJOJC1_2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35537\,
            in1 => \N__35464\,
            in2 => \_gnd_net_\,
            in3 => \N__35389\,
            lcout => \uart_drone.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.state_RNIL5IF_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47621\,
            in2 => \_gnd_net_\,
            in3 => \N__57834\,
            lcout => \pid_side.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_3_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__35564\,
            in1 => \N__35497\,
            in2 => \N__35426\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH4data_esr_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56479\,
            lcout => \frame_decoder_CH4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \Commands_frame_decoder.source_CH4data_esr_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56284\,
            lcout => \frame_decoder_CH4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \Commands_frame_decoder.source_CH4data_esr_2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56124\,
            lcout => \frame_decoder_CH4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \Commands_frame_decoder.source_CH4data_esr_3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55353\,
            lcout => \frame_decoder_CH4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \Commands_frame_decoder.source_CH4data_esr_4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53379\,
            lcout => \frame_decoder_CH4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \Commands_frame_decoder.source_CH4data_esr_5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55903\,
            lcout => \frame_decoder_CH4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \Commands_frame_decoder.source_CH4data_esr_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55733\,
            lcout => \frame_decoder_CH4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \Commands_frame_decoder.source_CH4data_ess_7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55567\,
            lcout => \frame_decoder_CH4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59097\,
            ce => \N__35760\,
            sr => \N__57525\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41160\,
            in2 => \N__41206\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35748\,
            in2 => \N__35742\,
            in3 => \N__35730\,
            lcout => \scaler_4.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_0\,
            carryout => \scaler_4.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35727\,
            in2 => \N__35721\,
            in3 => \N__35709\,
            lcout => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_1\,
            carryout => \scaler_4.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35706\,
            in2 => \N__35700\,
            in3 => \N__35688\,
            lcout => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_2\,
            carryout => \scaler_4.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35901\,
            in2 => \N__35895\,
            in3 => \N__35880\,
            lcout => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_3\,
            carryout => \scaler_4.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35877\,
            in2 => \N__35871\,
            in3 => \N__35859\,
            lcout => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_4\,
            carryout => \scaler_4.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35856\,
            in2 => \N__35847\,
            in3 => \N__35838\,
            lcout => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_5\,
            carryout => \scaler_4.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35835\,
            in2 => \_gnd_net_\,
            in3 => \N__35820\,
            lcout => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_6\,
            carryout => \scaler_4.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35766\,
            in2 => \N__42298\,
            in3 => \N__35817\,
            lcout => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35814\,
            lcout => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.N_1849_i_l_ofx_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35811\,
            in2 => \_gnd_net_\,
            in3 => \N__35783\,
            lcout => \scaler_4.N_1849_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_ctle_14_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45203\,
            in2 => \_gnd_net_\,
            in3 => \N__57845\,
            lcout => \ppm_encoder_1.pid_altitude_dv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI4N6K_2_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36148\,
            lcout => \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_6_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__36132\,
            in1 => \N__36126\,
            in2 => \N__40171\,
            in3 => \N__45354\,
            lcout => \ppm_encoder_1.throttleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59121\,
            ce => 'H',
            sr => \N__57542\
        );

    \ppm_encoder_1.throttle_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__36096\,
            in1 => \N__36090\,
            in2 => \N__45398\,
            in3 => \N__44216\,
            lcout => \ppm_encoder_1.throttleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59121\,
            ce => 'H',
            sr => \N__57542\
        );

    \ppm_encoder_1.throttle_9_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__36066\,
            in1 => \N__45344\,
            in2 => \N__40251\,
            in3 => \N__36036\,
            lcout => \ppm_encoder_1.throttleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59133\,
            ce => 'H',
            sr => \N__57552\
        );

    \ppm_encoder_1.aileron_4_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__36030\,
            in1 => \N__43248\,
            in2 => \N__45396\,
            in3 => \N__46951\,
            lcout => \ppm_encoder_1.aileronZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59133\,
            ce => 'H',
            sr => \N__57552\
        );

    \ppm_encoder_1.throttle_4_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__41872\,
            in1 => \N__45343\,
            in2 => \N__36021\,
            in3 => \N__35985\,
            lcout => \ppm_encoder_1.throttleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59133\,
            ce => 'H',
            sr => \N__57552\
        );

    \ppm_encoder_1.throttle_8_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__35979\,
            in1 => \N__35949\,
            in2 => \N__45397\,
            in3 => \N__40469\,
            lcout => \ppm_encoder_1.throttleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59133\,
            ce => 'H',
            sr => \N__57552\
        );

    \ppm_encoder_1.throttle_12_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__35943\,
            in1 => \N__45342\,
            in2 => \N__39952\,
            in3 => \N__35916\,
            lcout => \ppm_encoder_1.throttleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59133\,
            ce => 'H',
            sr => \N__57552\
        );

    \ppm_encoder_1.aileron_2_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__35910\,
            in1 => \N__41123\,
            in2 => \N__43792\,
            in3 => \N__45340\,
            lcout => \ppm_encoder_1.aileronZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59148\,
            ce => 'H',
            sr => \N__57561\
        );

    \ppm_encoder_1.throttle_0_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__45333\,
            in1 => \N__36249\,
            in2 => \_gnd_net_\,
            in3 => \N__43660\,
            lcout => \ppm_encoder_1.throttleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59148\,
            ce => 'H',
            sr => \N__57561\
        );

    \ppm_encoder_1.throttle_7_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__36228\,
            in1 => \N__36214\,
            in2 => \N__45395\,
            in3 => \N__40342\,
            lcout => \ppm_encoder_1.throttleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59148\,
            ce => 'H',
            sr => \N__57561\
        );

    \ppm_encoder_1.elevator_10_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__37917\,
            in1 => \N__37884\,
            in2 => \N__45394\,
            in3 => \N__40520\,
            lcout => \ppm_encoder_1.elevatorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59148\,
            ce => 'H',
            sr => \N__57561\
        );

    \ppm_encoder_1.elevator_2_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__37791\,
            in1 => \N__37773\,
            in2 => \N__47032\,
            in3 => \N__45341\,
            lcout => \ppm_encoder_1.elevatorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59148\,
            ce => 'H',
            sr => \N__57561\
        );

    \ppm_encoder_1.elevator_8_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__37995\,
            in1 => \N__37968\,
            in2 => \N__45388\,
            in3 => \N__40455\,
            lcout => \ppm_encoder_1.elevatorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59160\,
            ce => 'H',
            sr => \N__57572\
        );

    \ppm_encoder_1.aileron_10_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__43043\,
            in1 => \N__36186\,
            in2 => \N__45399\,
            in3 => \N__40496\,
            lcout => \ppm_encoder_1.aileronZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59160\,
            ce => 'H',
            sr => \N__57572\
        );

    \ppm_encoder_1.aileron_13_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__48062\,
            in1 => \N__36180\,
            in2 => \N__38175\,
            in3 => \N__45358\,
            lcout => \ppm_encoder_1.aileronZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59160\,
            ce => 'H',
            sr => \N__57572\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47163\,
            in1 => \N__37821\,
            in2 => \_gnd_net_\,
            in3 => \N__38124\,
            lcout => \ppm_encoder_1.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI14DT_2_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36170\,
            in2 => \_gnd_net_\,
            in3 => \N__57865\,
            lcout => \dron_frame_decoder_1.N_489_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNICVO11_2_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__36291\,
            in1 => \N__38246\,
            in2 => \N__36282\,
            in3 => \N__38230\,
            lcout => \pid_front.error_p_reg_esr_RNICVO11Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__36311\,
            in1 => \N__36263\,
            in2 => \_gnd_net_\,
            in3 => \N__50866\,
            lcout => \pid_front.un1_pid_prereg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101101001"
        )
    port map (
            in0 => \N__50867\,
            in1 => \N__36312\,
            in2 => \N__36267\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.un1_pid_prereg_2\,
            ltout => \pid_front.un1_pid_prereg_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIJCSG_2_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36294\,
            in3 => \N__36290\,
            lcout => \pid_front.error_p_reg_esr_RNIJCSGZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__38103\,
            in1 => \N__38082\,
            in2 => \_gnd_net_\,
            in3 => \N__49301\,
            lcout => \pid_front.un1_pid_prereg_0\,
            ltout => \pid_front.un1_pid_prereg_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIH7Q01_1_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__38568\,
            in1 => \N__36278\,
            in2 => \N__36270\,
            in3 => \N__38551\,
            lcout => \pid_front.error_p_reg_esr_RNIH7Q01Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_3_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59191\,
            ce => \N__49372\,
            sr => \N__57583\
        );

    \pid_front.error_d_reg_prev_esr_2_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59191\,
            ce => \N__49372\,
            sr => \N__57583\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52291\,
            lcout => \drone_H_disp_front_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50779\,
            lcout => \drone_H_disp_front_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50398\,
            lcout => \drone_H_disp_front_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52693\,
            lcout => \drone_H_disp_front_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52598\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52477\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53211\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52391\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59201\,
            ce => \N__36354\,
            sr => \N__57597\
        );

    \pid_front.error_d_reg_prev_esr_0_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49460\,
            in2 => \N__56939\,
            in3 => \N__56935\,
            lcout => \pid_front.error_d_reg_prevZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \pid_front.un1_pid_prereg_cry_0\,
            clk => \N__59216\,
            ce => \N__49369\,
            sr => \N__57603\
        );

    \pid_front.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50519\,
            in2 => \_gnd_net_\,
            in3 => \N__36339\,
            lcout => \pid_front.un1_pid_prereg_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_0\,
            carryout => \pid_front.un1_pid_prereg_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_2_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38208\,
            in2 => \N__38589\,
            in3 => \N__36315\,
            lcout => \pid_front.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_1\,
            carryout => \pid_front.un1_pid_prereg_cry_0_0\,
            clk => \N__59216\,
            ce => \N__49369\,
            sr => \N__57603\
        );

    \pid_front.pid_prereg_esr_3_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38535\,
            in2 => \N__36792\,
            in3 => \N__36756\,
            lcout => \pid_front.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_0_0\,
            carryout => \pid_front.un1_pid_prereg_cry_1_0\,
            clk => \N__59216\,
            ce => \N__49369\,
            sr => \N__57603\
        );

    \pid_front.pid_prereg_esr_4_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36753\,
            in2 => \N__36744\,
            in3 => \N__36690\,
            lcout => \pid_front.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_1_0\,
            carryout => \pid_front.un1_pid_prereg_cry_2\,
            clk => \N__59216\,
            ce => \N__49369\,
            sr => \N__57603\
        );

    \pid_front.pid_prereg_esr_5_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38217\,
            in2 => \N__38070\,
            in3 => \N__36645\,
            lcout => \pid_front.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_2\,
            carryout => \pid_front.un1_pid_prereg_cry_3\,
            clk => \N__59216\,
            ce => \N__49369\,
            sr => \N__57603\
        );

    \pid_front.pid_prereg_esr_6_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38006\,
            in2 => \N__36642\,
            in3 => \N__36609\,
            lcout => \pid_front.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_3\,
            carryout => \pid_front.un1_pid_prereg_cry_4\,
            clk => \N__59216\,
            ce => \N__49369\,
            sr => \N__57603\
        );

    \pid_front.pid_prereg_esr_7_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36605\,
            in2 => \N__36594\,
            in3 => \N__36555\,
            lcout => \pid_front.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_4\,
            carryout => \pid_front.un1_pid_prereg_cry_5\,
            clk => \N__59216\,
            ce => \N__49369\,
            sr => \N__57603\
        );

    \pid_front.pid_prereg_esr_8_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36552\,
            in2 => \N__36540\,
            in3 => \N__36495\,
            lcout => \pid_front.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \pid_front.un1_pid_prereg_cry_6\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_9_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36492\,
            in2 => \N__36474\,
            in3 => \N__36435\,
            lcout => \pid_front.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_6\,
            carryout => \pid_front.un1_pid_prereg_cry_7\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_10_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36432\,
            in2 => \N__36419\,
            in3 => \N__37095\,
            lcout => \pid_front.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_7\,
            carryout => \pid_front.un1_pid_prereg_cry_8\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_11_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37092\,
            in2 => \N__37083\,
            in3 => \N__37038\,
            lcout => \pid_front.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_8\,
            carryout => \pid_front.un1_pid_prereg_cry_9\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_12_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37035\,
            in2 => \N__37023\,
            in3 => \N__36987\,
            lcout => \pid_front.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_9\,
            carryout => \pid_front.un1_pid_prereg_cry_10\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_13_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36984\,
            in2 => \N__36969\,
            in3 => \N__36924\,
            lcout => \pid_front.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_10\,
            carryout => \pid_front.un1_pid_prereg_cry_11\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_14_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36921\,
            in2 => \N__36912\,
            in3 => \N__36894\,
            lcout => \pid_front.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_11\,
            carryout => \pid_front.un1_pid_prereg_cry_12\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_15_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36891\,
            in2 => \N__36879\,
            in3 => \N__36858\,
            lcout => \pid_front.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_12\,
            carryout => \pid_front.un1_pid_prereg_cry_13\,
            clk => \N__59233\,
            ce => \N__49367\,
            sr => \N__57610\
        );

    \pid_front.pid_prereg_esr_16_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36855\,
            in2 => \N__36846\,
            in3 => \N__36825\,
            lcout => \pid_front.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_12_23_0_\,
            carryout => \pid_front.un1_pid_prereg_cry_14\,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \pid_front.pid_prereg_esr_17_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36822\,
            in2 => \N__36813\,
            in3 => \N__36795\,
            lcout => \pid_front.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_14\,
            carryout => \pid_front.un1_pid_prereg_cry_15\,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \pid_front.pid_prereg_esr_18_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37299\,
            in2 => \N__37290\,
            in3 => \N__37269\,
            lcout => \pid_front.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_15\,
            carryout => \pid_front.un1_pid_prereg_cry_16\,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \pid_front.pid_prereg_esr_19_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37266\,
            in2 => \N__37257\,
            in3 => \N__37239\,
            lcout => \pid_front.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_16\,
            carryout => \pid_front.un1_pid_prereg_cry_17\,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \pid_front.pid_prereg_esr_20_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37236\,
            in2 => \N__37227\,
            in3 => \N__37206\,
            lcout => \pid_front.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_17\,
            carryout => \pid_front.un1_pid_prereg_cry_18\,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \pid_front.pid_prereg_esr_21_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37203\,
            in2 => \N__37194\,
            in3 => \N__37173\,
            lcout => \pid_front.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_18\,
            carryout => \pid_front.un1_pid_prereg_cry_19\,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \pid_front.pid_prereg_esr_22_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37170\,
            in2 => \N__42516\,
            in3 => \N__37152\,
            lcout => \pid_front.pid_preregZ0Z_22\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_19\,
            carryout => \pid_front.un1_pid_prereg_cry_20\,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \pid_front.pid_prereg_esr_23_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37320\,
            in2 => \_gnd_net_\,
            in3 => \N__37149\,
            lcout => \pid_front.pid_preregZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59251\,
            ce => \N__49365\,
            sr => \N__57617\
        );

    \Commands_frame_decoder.source_CH3data_esr_0_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56506\,
            lcout => front_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \Commands_frame_decoder.source_CH3data_esr_1_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56311\,
            lcout => front_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \Commands_frame_decoder.source_CH3data_esr_2_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56142\,
            lcout => front_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \Commands_frame_decoder.source_CH3data_esr_3_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__55356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => front_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \Commands_frame_decoder.source_CH3data_esr_4_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53409\,
            lcout => front_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \Commands_frame_decoder.source_CH3data_esr_5_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55932\,
            lcout => front_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \Commands_frame_decoder.source_CH3data_esr_6_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55755\,
            lcout => front_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \Commands_frame_decoder.source_CH3data_ess_7_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55584\,
            lcout => front_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59266\,
            ce => \N__37338\,
            sr => \N__57624\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39417\,
            lcout => \drone_H_disp_front_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNO_0_23_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__42539\,
            in1 => \N__42609\,
            in2 => \N__42552\,
            in3 => \N__42610\,
            lcout => \pid_front.un1_pid_prereg_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_8_l_ofx_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__39411\,
            in1 => \_gnd_net_\,
            in2 => \N__37311\,
            in3 => \N__39398\,
            lcout => \pid_front.error_axb_8_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_7_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37307\,
            in2 => \_gnd_net_\,
            in3 => \N__39410\,
            lcout => \pid_front.error_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39397\,
            lcout => \drone_H_disp_front_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__59501\,
            in1 => \_gnd_net_\,
            in2 => \N__43059\,
            in3 => \N__37362\,
            lcout => \pid_front.un1_pid_prereg_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI8QE61_20_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__37361\,
            in1 => \N__43055\,
            in2 => \_gnd_net_\,
            in3 => \N__59500\,
            lcout => \pid_front.un1_pid_prereg_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIFCSD1_0_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__47684\,
            in1 => \N__39717\,
            in2 => \N__39595\,
            in3 => \N__57828\,
            lcout => \pid_alt.state_RNIFCSD1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_data_valid_esr_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39718\,
            lcout => pid_altitude_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59080\,
            ce => \N__39840\,
            sr => \N__57519\
        );

    \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37595\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \ppm_encoder_1.un1_rudder_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37427\,
            in2 => \_gnd_net_\,
            in3 => \N__37347\,
            lcout => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_6\,
            carryout => \ppm_encoder_1.un1_rudder_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39800\,
            in2 => \_gnd_net_\,
            in3 => \N__37344\,
            lcout => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_7\,
            carryout => \ppm_encoder_1.un1_rudder_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39830\,
            in2 => \_gnd_net_\,
            in3 => \N__37341\,
            lcout => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_8\,
            carryout => \ppm_encoder_1.un1_rudder_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39782\,
            in2 => \_gnd_net_\,
            in3 => \N__37410\,
            lcout => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_9\,
            carryout => \ppm_encoder_1.un1_rudder_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39552\,
            in3 => \N__37407\,
            lcout => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_10\,
            carryout => \ppm_encoder_1.un1_rudder_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39528\,
            in2 => \_gnd_net_\,
            in3 => \N__37404\,
            lcout => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_11\,
            carryout => \ppm_encoder_1.un1_rudder_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39761\,
            in2 => \N__42315\,
            in3 => \N__37401\,
            lcout => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_12\,
            carryout => \ppm_encoder_1.un1_rudder_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_14_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37476\,
            in2 => \_gnd_net_\,
            in3 => \N__37398\,
            lcout => \ppm_encoder_1.rudderZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59088\,
            ce => \N__46776\,
            sr => \N__57529\
        );

    \scaler_4.un2_source_data_0_cry_1_c_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41235\,
            in2 => \N__41139\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_6_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37388\,
            in2 => \N__41245\,
            in3 => \N__37395\,
            lcout => scaler_4_data_6,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_1\,
            carryout => \scaler_4.un2_source_data_0_cry_2\,
            clk => \N__59094\,
            ce => \N__37466\,
            sr => \N__57535\
        );

    \scaler_4.source_data_1_esr_7_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37373\,
            in2 => \N__37392\,
            in3 => \N__37380\,
            lcout => scaler_4_data_7,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_2\,
            carryout => \scaler_4.un2_source_data_0_cry_3\,
            clk => \N__59094\,
            ce => \N__37466\,
            sr => \N__57535\
        );

    \scaler_4.source_data_1_esr_8_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37559\,
            in2 => \N__37377\,
            in3 => \N__37365\,
            lcout => scaler_4_data_8,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_3\,
            carryout => \scaler_4.un2_source_data_0_cry_4\,
            clk => \N__59094\,
            ce => \N__37466\,
            sr => \N__57535\
        );

    \scaler_4.source_data_1_esr_9_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37544\,
            in2 => \N__37563\,
            in3 => \N__37551\,
            lcout => scaler_4_data_9,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_4\,
            carryout => \scaler_4.un2_source_data_0_cry_5\,
            clk => \N__59094\,
            ce => \N__37466\,
            sr => \N__57535\
        );

    \scaler_4.source_data_1_esr_10_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37529\,
            in2 => \N__37548\,
            in3 => \N__37536\,
            lcout => scaler_4_data_10,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_5\,
            carryout => \scaler_4.un2_source_data_0_cry_6\,
            clk => \N__59094\,
            ce => \N__37466\,
            sr => \N__57535\
        );

    \scaler_4.source_data_1_esr_11_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37514\,
            in2 => \N__37533\,
            in3 => \N__37521\,
            lcout => scaler_4_data_11,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_6\,
            carryout => \scaler_4.un2_source_data_0_cry_7\,
            clk => \N__59094\,
            ce => \N__37466\,
            sr => \N__57535\
        );

    \scaler_4.source_data_1_esr_12_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37502\,
            in2 => \N__37518\,
            in3 => \N__37506\,
            lcout => scaler_4_data_12,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_7\,
            carryout => \scaler_4.un2_source_data_0_cry_8\,
            clk => \N__59094\,
            ce => \N__37466\,
            sr => \N__57535\
        );

    \scaler_4.source_data_1_esr_13_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37503\,
            in2 => \N__37491\,
            in3 => \N__37482\,
            lcout => scaler_4_data_13,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_9\,
            clk => \N__59102\,
            ce => \N__37467\,
            sr => \N__57543\
        );

    \scaler_4.source_data_1_esr_14_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37479\,
            lcout => scaler_4_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59102\,
            ce => \N__37467\,
            sr => \N__57543\
        );

    \ppm_encoder_1.rudder_7_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__37437\,
            in1 => \N__37428\,
            in2 => \N__45370\,
            in3 => \N__40576\,
            lcout => \ppm_encoder_1.rudderZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59111\,
            ce => 'H',
            sr => \N__57553\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_0_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43629\,
            in2 => \_gnd_net_\,
            in3 => \N__43538\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_134_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011110100"
        )
    port map (
            in0 => \N__43590\,
            in1 => \N__37634\,
            in2 => \N__37644\,
            in3 => \N__42654\,
            lcout => ppm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59111\,
            ce => 'H',
            sr => \N__57553\
        );

    \ppm_encoder_1.throttle_2_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__37623\,
            in1 => \N__37614\,
            in2 => \N__45371\,
            in3 => \N__46993\,
            lcout => \ppm_encoder_1.throttleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59111\,
            ce => 'H',
            sr => \N__57553\
        );

    \ppm_encoder_1.elevator_4_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__37737\,
            in1 => \N__37761\,
            in2 => \N__45297\,
            in3 => \N__41852\,
            lcout => \ppm_encoder_1.elevatorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \ppm_encoder_1.elevator_5_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__37728\,
            in1 => \N__37698\,
            in2 => \N__43199\,
            in3 => \N__45200\,
            lcout => \ppm_encoder_1.elevatorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \ppm_encoder_1.elevator_9_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__37929\,
            in1 => \N__37959\,
            in2 => \N__45298\,
            in3 => \N__40227\,
            lcout => \ppm_encoder_1.elevatorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \ppm_encoder_1.rudder_6_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__37596\,
            in1 => \N__45190\,
            in2 => \_gnd_net_\,
            in3 => \N__40610\,
            lcout => \ppm_encoder_1.rudderZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \ppm_encoder_1.elevator_11_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__37875\,
            in1 => \N__37842\,
            in2 => \N__45296\,
            in3 => \N__40099\,
            lcout => \ppm_encoder_1.elevatorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \ppm_encoder_1.aileron_5_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__43274\,
            in1 => \N__37578\,
            in2 => \N__45295\,
            in3 => \N__51269\,
            lcout => \ppm_encoder_1.aileronZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \pid_alt.state_1_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39599\,
            lcout => \pid_alt.N_72_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \ppm_encoder_1.elevator_6_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__45186\,
            in1 => \N__37689\,
            in2 => \N__40149\,
            in3 => \N__37656\,
            lcout => \ppm_encoder_1.elevatorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59118\,
            ce => 'H',
            sr => \N__57562\
        );

    \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45428\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41480\,
            in2 => \N__42316\,
            in3 => \N__37794\,
            lcout => \ppm_encoder_1.un1_elevator_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_0\,
            carryout => \ppm_encoder_1.un1_elevator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37790\,
            in2 => \_gnd_net_\,
            in3 => \N__37767\,
            lcout => \ppm_encoder_1.un1_elevator_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_1\,
            carryout => \ppm_encoder_1.un1_elevator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43886\,
            in2 => \N__42317\,
            in3 => \N__37764\,
            lcout => \ppm_encoder_1.un1_elevator_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_2\,
            carryout => \ppm_encoder_1.un1_elevator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37760\,
            in2 => \_gnd_net_\,
            in3 => \N__37731\,
            lcout => \ppm_encoder_1.un1_elevator_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_3\,
            carryout => \ppm_encoder_1.un1_elevator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37727\,
            in2 => \_gnd_net_\,
            in3 => \N__37692\,
            lcout => \ppm_encoder_1.un1_elevator_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_4\,
            carryout => \ppm_encoder_1.un1_elevator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42278\,
            in2 => \N__37688\,
            in3 => \N__37650\,
            lcout => \ppm_encoder_1.un1_elevator_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_5\,
            carryout => \ppm_encoder_1.un1_elevator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40292\,
            in2 => \_gnd_net_\,
            in3 => \N__37647\,
            lcout => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_6\,
            carryout => \ppm_encoder_1.un1_elevator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37994\,
            in2 => \_gnd_net_\,
            in3 => \N__37962\,
            lcout => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37955\,
            in2 => \_gnd_net_\,
            in3 => \N__37920\,
            lcout => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_8\,
            carryout => \ppm_encoder_1.un1_elevator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37916\,
            in2 => \_gnd_net_\,
            in3 => \N__37878\,
            lcout => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_9\,
            carryout => \ppm_encoder_1.un1_elevator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37874\,
            in2 => \_gnd_net_\,
            in3 => \N__37833\,
            lcout => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_10\,
            carryout => \ppm_encoder_1.un1_elevator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39890\,
            in2 => \_gnd_net_\,
            in3 => \N__37830\,
            lcout => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_11\,
            carryout => \ppm_encoder_1.un1_elevator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38153\,
            in2 => \N__42352\,
            in3 => \N__37827\,
            lcout => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_12\,
            carryout => \ppm_encoder_1.un1_elevator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_esr_14_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37824\,
            lcout => \ppm_encoder_1.elevatorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59145\,
            ce => \N__46777\,
            sr => \N__57577\
        );

    \ppm_encoder_1.throttle_RNIM4PT2_13_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__44372\,
            in1 => \N__37820\,
            in2 => \N__41361\,
            in3 => \N__44069\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIMC2D6_13_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44400\,
            in2 => \N__37797\,
            in3 => \N__38187\,
            lcout => \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI68LH2_13_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__38122\,
            in1 => \N__38170\,
            in2 => \N__44202\,
            in3 => \N__45553\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51431\,
            in1 => \N__38181\,
            in2 => \_gnd_net_\,
            in3 => \N__38171\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_13_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__38123\,
            in1 => \N__38157\,
            in2 => \N__45401\,
            in3 => \N__38130\,
            lcout => \ppm_encoder_1.elevatorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59157\,
            ce => 'H',
            sr => \N__57584\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38109\,
            lcout => \drone_H_disp_front_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__38102\,
            in1 => \N__38081\,
            in2 => \_gnd_net_\,
            in3 => \N__49295\,
            lcout => \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNIOBP11_5_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__38232\,
            in1 => \N__38061\,
            in2 => \N__38250\,
            in3 => \N__38055\,
            lcout => \pid_front.error_d_reg_esr_RNIOBP11Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNI1EE8_5_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38046\,
            in1 => \N__38293\,
            in2 => \_gnd_net_\,
            in3 => \N__53080\,
            lcout => \pid_front.un1_pid_prereg_40_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIUAE8_4_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__38279\,
            in1 => \N__38258\,
            in2 => \_gnd_net_\,
            in3 => \N__59425\,
            lcout => \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4\,
            ltout => \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNIVOSG_5_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__38047\,
            in1 => \N__38294\,
            in2 => \N__38016\,
            in3 => \N__53081\,
            lcout => \pid_front.error_d_reg_esr_RNIVOSGZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_5_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__53082\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59188\,
            ce => \N__49373\,
            sr => \N__57604\
        );

    \pid_front.error_d_reg_prev_esr_4_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__59427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_reg_prevZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59188\,
            ce => \N__49373\,
            sr => \N__57604\
        );

    \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__38280\,
            in1 => \N__38259\,
            in2 => \_gnd_net_\,
            in3 => \N__59426\,
            lcout => \pid_front.un1_pid_prereg_17\,
            ltout => \pid_front.un1_pid_prereg_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIPISG_3_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38235\,
            in3 => \N__38231\,
            lcout => \pid_front.error_p_reg_esr_RNIPISGZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI6MF7_0_1_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__46919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38201\,
            lcout => \pid_front.N_1427_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI4KF7_0_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38396\,
            in2 => \_gnd_net_\,
            in3 => \N__38348\,
            lcout => OPEN,
            ltout => \pid_front.error_p_reg_esr_RNI4KF7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNINGRV_1_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011111100"
        )
    port map (
            in0 => \N__38588\,
            in1 => \N__56894\,
            in2 => \N__38211\,
            in3 => \N__38325\,
            lcout => \pid_front.error_d_reg_esr_RNINGRVZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40721\,
            lcout => \drone_H_disp_front_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNI6MF7_1_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__46920\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38202\,
            lcout => \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1\,
            ltout => \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIUQTF_0_1_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38592\,
            in3 => \N__38552\,
            lcout => \pid_front.un1_pid_prereg\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_3_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38574\,
            lcout => \pid_front.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIUQTF_1_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38564\,
            in2 => \_gnd_net_\,
            in3 => \N__38553\,
            lcout => \pid_front.error_p_reg_esr_RNIUQTFZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__38528\,
            in1 => \N__38490\,
            in2 => \_gnd_net_\,
            in3 => \N__38457\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38415\,
            lcout => \drone_H_disp_front_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38406\,
            lcout => \drone_H_disp_front_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_RNIPLTF_1_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__38397\,
            in1 => \N__38347\,
            in2 => \N__56893\,
            in3 => \N__38324\,
            lcout => \pid_front.un1_pid_prereg_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38313\,
            lcout => \drone_H_disp_front_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_2_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38925\,
            lcout => \pid_front.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39360\,
            lcout => \drone_H_disp_front_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_0_c_inv_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38871\,
            in2 => \_gnd_net_\,
            in3 => \N__38902\,
            lcout => \pid_front.error_axb_0\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \pid_front.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_0_c_RNIC7KB_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38865\,
            in2 => \_gnd_net_\,
            in3 => \N__38811\,
            lcout => \pid_front.error_1\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_0\,
            carryout => \pid_front.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_1_c_RNIEALB_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38808\,
            in2 => \_gnd_net_\,
            in3 => \N__38763\,
            lcout => \pid_front.error_2\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_1\,
            carryout => \pid_front.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_2_c_RNIGDMB_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38760\,
            in2 => \_gnd_net_\,
            in3 => \N__38712\,
            lcout => \pid_front.error_3\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_2\,
            carryout => \pid_front.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_3_c_RNIABAG_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38709\,
            in2 => \N__38703\,
            in3 => \N__38652\,
            lcout => \pid_front.error_4\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_3\,
            carryout => \pid_front.error_cry_0_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38649\,
            in2 => \N__38643\,
            in3 => \N__38595\,
            lcout => \pid_front.error_5\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_0_0\,
            carryout => \pid_front.error_cry_1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39342\,
            in2 => \N__39336\,
            in3 => \N__39294\,
            lcout => \pid_front.error_6\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_1_0\,
            carryout => \pid_front.error_cry_2_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_2_0_c_RNIU61K_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39291\,
            in2 => \N__39279\,
            in3 => \N__39231\,
            lcout => \pid_front.error_7\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_2_0\,
            carryout => \pid_front.error_cry_3_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39228\,
            in2 => \N__39219\,
            in3 => \N__39171\,
            lcout => \pid_front.error_8\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \pid_front.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_4_c_RNILNBG_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50799\,
            in2 => \N__39168\,
            in3 => \N__39120\,
            lcout => \pid_front.error_9\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_4\,
            carryout => \pid_front.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_5_c_RNIVNFF_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39117\,
            in2 => \N__39111\,
            in3 => \N__39060\,
            lcout => \pid_front.error_10\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_5\,
            carryout => \pid_front.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_6_c_RNI3VJG_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39057\,
            in2 => \_gnd_net_\,
            in3 => \N__39012\,
            lcout => \pid_front.error_11\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_6\,
            carryout => \pid_front.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_7_c_RNIAPPM_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39009\,
            in2 => \N__39402\,
            in3 => \N__38970\,
            lcout => \pid_front.error_12\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_7\,
            carryout => \pid_front.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_8_c_RNIAC2E_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38967\,
            in2 => \N__40731\,
            in3 => \N__38928\,
            lcout => \pid_front.error_13\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_8\,
            carryout => \pid_front.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_9_c_RNIDG3E_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39507\,
            in2 => \N__39384\,
            in3 => \N__39459\,
            lcout => \pid_front.error_14\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_9\,
            carryout => \pid_front.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_10_c_RNINTDI_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__39369\,
            in1 => \N__39383\,
            in2 => \_gnd_net_\,
            in3 => \N__39456\,
            lcout => \pid_front.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50403\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59263\,
            ce => \N__50697\,
            sr => \N__57636\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52708\,
            lcout => \drone_H_disp_front_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59263\,
            ce => \N__50697\,
            sr => \N__57636\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52597\,
            lcout => \drone_H_disp_front_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59263\,
            ce => \N__50697\,
            sr => \N__57636\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53228\,
            lcout => \drone_H_disp_front_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59263\,
            ce => \N__50697\,
            sr => \N__57636\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52395\,
            lcout => \drone_H_disp_front_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59263\,
            ce => \N__50697\,
            sr => \N__57636\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52300\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59263\,
            ce => \N__50697\,
            sr => \N__57636\
        );

    \pid_alt.state_RNIH1EN_0_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39600\,
            in2 => \_gnd_net_\,
            in3 => \N__57836\,
            lcout => \pid_alt.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_data_valid_esr_RNO_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39588\,
            in2 => \_gnd_net_\,
            in3 => \N__57870\,
            lcout => \pid_alt.state_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_9_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__39831\,
            in1 => \N__39813\,
            in2 => \N__45202\,
            in3 => \N__40204\,
            lcout => \ppm_encoder_1.rudderZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59091\,
            ce => 'H',
            sr => \N__57530\
        );

    \ppm_encoder_1.rudder_8_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__39807\,
            in1 => \N__39801\,
            in2 => \N__46231\,
            in3 => \N__45132\,
            lcout => \ppm_encoder_1.rudderZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59091\,
            ce => 'H',
            sr => \N__57530\
        );

    \ppm_encoder_1.rudder_10_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__39783\,
            in1 => \N__39768\,
            in2 => \N__45201\,
            in3 => \N__46291\,
            lcout => \ppm_encoder_1.rudderZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59091\,
            ce => 'H',
            sr => \N__57530\
        );

    \ppm_encoder_1.rudder_13_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__39762\,
            in1 => \N__39744\,
            in2 => \N__45374\,
            in3 => \N__44365\,
            lcout => \ppm_encoder_1.rudderZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59098\,
            ce => 'H',
            sr => \N__57536\
        );

    \pid_alt.state_0_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__39584\,
            in1 => \N__47705\,
            in2 => \_gnd_net_\,
            in3 => \N__39676\,
            lcout => \pid_alt.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59098\,
            ce => 'H',
            sr => \N__57536\
        );

    \ppm_encoder_1.rudder_11_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__39551\,
            in1 => \N__39534\,
            in2 => \N__45372\,
            in3 => \N__40850\,
            lcout => \ppm_encoder_1.rudderZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59098\,
            ce => 'H',
            sr => \N__57536\
        );

    \ppm_encoder_1.rudder_12_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__39527\,
            in1 => \N__39513\,
            in2 => \N__45373\,
            in3 => \N__46712\,
            lcout => \ppm_encoder_1.rudderZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59098\,
            ce => 'H',
            sr => \N__57536\
        );

    \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__39859\,
            in1 => \N__39907\,
            in2 => \N__45558\,
            in3 => \N__44189\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__39953\,
            in1 => \N__46708\,
            in2 => \N__41353\,
            in3 => \N__44053\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47178\,
            in1 => \N__39954\,
            in2 => \_gnd_net_\,
            in3 => \N__39860\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51409\,
            in2 => \N__39930\,
            in3 => \N__39908\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_12_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__39909\,
            in1 => \N__45294\,
            in2 => \N__39927\,
            in3 => \N__45590\,
            lcout => \ppm_encoder_1.aileronZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59105\,
            ce => 'H',
            sr => \N__57544\
        );

    \ppm_encoder_1.elevator_12_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__39861\,
            in1 => \N__39897\,
            in2 => \N__45375\,
            in3 => \N__39873\,
            lcout => \ppm_encoder_1.elevatorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59105\,
            ce => 'H',
            sr => \N__57544\
        );

    \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__40000\,
            in1 => \N__40851\,
            in2 => \N__44070\,
            in3 => \N__41357\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47490\,
            in2 => \N__39849\,
            in3 => \N__39846\,
            lcout => \ppm_encoder_1.elevator_RNIC22D6Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__40100\,
            in1 => \N__40063\,
            in2 => \N__44201\,
            in3 => \N__45513\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47164\,
            in1 => \N__40001\,
            in2 => \_gnd_net_\,
            in3 => \N__40101\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51426\,
            in2 => \N__40083\,
            in3 => \N__40064\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_11_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__40065\,
            in1 => \N__45389\,
            in2 => \N__43010\,
            in3 => \N__40080\,
            lcout => \ppm_encoder_1.aileronZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59112\,
            ce => 'H',
            sr => \N__57554\
        );

    \ppm_encoder_1.throttle_11_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__40053\,
            in1 => \N__40017\,
            in2 => \N__40005\,
            in3 => \N__45390\,
            lcout => \ppm_encoder_1.throttleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59112\,
            ce => 'H',
            sr => \N__57554\
        );

    \ppm_encoder_1.throttle_RNI04QV2_9_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__40249\,
            in1 => \N__40205\,
            in2 => \N__41352\,
            in3 => \N__44054\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIV9PO6_9_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46161\,
            in2 => \N__39987\,
            in3 => \N__39960\,
            lcout => \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51410\,
            in1 => \N__40212\,
            in2 => \_gnd_net_\,
            in3 => \N__39981\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_9_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44660\,
            in2 => \N__39984\,
            in3 => \N__40188\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59122\,
            ce => \N__44613\,
            sr => \N__57563\
        );

    \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__40225\,
            in1 => \N__39980\,
            in2 => \N__45532\,
            in3 => \N__44166\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47171\,
            in1 => \N__40250\,
            in2 => \_gnd_net_\,
            in3 => \N__40226\,
            lcout => \ppm_encoder_1.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__46389\,
            in1 => \N__46566\,
            in2 => \N__46140\,
            in3 => \N__40206\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__46565\,
            in1 => \N__46388\,
            in2 => \_gnd_net_\,
            in3 => \N__46070\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIQTPV2_6_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__40172\,
            in1 => \N__40606\,
            in2 => \N__44073\,
            in3 => \N__41327\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIGQOO6_6_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45834\,
            in2 => \N__40182\,
            in3 => \N__40179\,
            lcout => \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIAH7O2_6_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__40111\,
            in1 => \N__45483\,
            in2 => \N__40148\,
            in3 => \N__44125\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47165\,
            in1 => \N__40173\,
            in2 => \_gnd_net_\,
            in3 => \N__40144\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_292_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__40112\,
            in1 => \_gnd_net_\,
            in2 => \N__40128\,
            in3 => \N__51456\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_6_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__40125\,
            in1 => \N__40113\,
            in2 => \N__42975\,
            in3 => \N__45363\,
            lcout => \ppm_encoder_1.aileronZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59134\,
            ce => 'H',
            sr => \N__57573\
        );

    \ppm_encoder_1.throttle_RNISVPV2_7_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__40343\,
            in1 => \N__40577\,
            in2 => \N__44071\,
            in3 => \N__41332\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNILVOO6_7_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__45924\,
            in1 => \_gnd_net_\,
            in2 => \N__40353\,
            in3 => \N__40350\,
            lcout => \ppm_encoder_1.throttle_RNILVOO6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNICJ7O2_7_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__40264\,
            in1 => \N__40309\,
            in2 => \N__44200\,
            in3 => \N__45516\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47169\,
            in1 => \N__40344\,
            in2 => \_gnd_net_\,
            in3 => \N__40265\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51436\,
            in2 => \N__40326\,
            in3 => \N__40310\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_7_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__40311\,
            in1 => \N__40323\,
            in2 => \N__42930\,
            in3 => \N__45362\,
            lcout => \ppm_encoder_1.aileronZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59149\,
            ce => 'H',
            sr => \N__57578\
        );

    \ppm_encoder_1.elevator_7_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__40266\,
            in1 => \N__40299\,
            in2 => \N__45400\,
            in3 => \N__40293\,
            lcout => \ppm_encoder_1.elevatorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59149\,
            ce => 'H',
            sr => \N__57578\
        );

    \ppm_encoder_1.throttle_RNIU1QV2_8_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__40475\,
            in1 => \N__46232\,
            in2 => \N__44072\,
            in3 => \N__41348\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__46257\,
            in1 => \_gnd_net_\,
            in2 => \N__40254\,
            in3 => \N__40482\,
            lcout => \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__40453\,
            in1 => \N__40417\,
            in2 => \N__44190\,
            in3 => \N__45546\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47177\,
            in1 => \N__40476\,
            in2 => \_gnd_net_\,
            in3 => \N__40454\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__51415\,
            in1 => \_gnd_net_\,
            in2 => \N__40434\,
            in3 => \N__40418\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_8_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__40419\,
            in1 => \N__42885\,
            in2 => \N__45402\,
            in3 => \N__40431\,
            lcout => \ppm_encoder_1.aileronZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59161\,
            ce => 'H',
            sr => \N__57585\
        );

    \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__44059\,
            in1 => \N__40385\,
            in2 => \N__41356\,
            in3 => \N__44816\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__44325\,
            in1 => \_gnd_net_\,
            in2 => \N__40407\,
            in3 => \N__40404\,
            lcout => \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__40397\,
            in1 => \N__40364\,
            in2 => \N__45561\,
            in3 => \N__44194\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47150\,
            in1 => \N__40398\,
            in2 => \_gnd_net_\,
            in3 => \N__40386\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__51452\,
            in1 => \_gnd_net_\,
            in2 => \N__40368\,
            in3 => \N__40365\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__45759\,
            in1 => \N__46570\,
            in2 => \N__46444\,
            in3 => \N__40611\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIGUOT2_10_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__44058\,
            in1 => \N__40553\,
            in2 => \N__41355\,
            in3 => \N__46302\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48854\,
            lcout => \ppm_encoder_1.N_2150_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI02LH2_10_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__40526\,
            in1 => \N__40502\,
            in2 => \N__45560\,
            in3 => \N__44195\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI7T1D6_10_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__46608\,
            in1 => \_gnd_net_\,
            in2 => \N__40590\,
            in3 => \N__40587\,
            lcout => \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__45900\,
            in1 => \N__46569\,
            in2 => \N__46445\,
            in3 => \N__40581\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40557\,
            in1 => \N__47128\,
            in2 => \_gnd_net_\,
            in3 => \N__40527\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51451\,
            in2 => \N__40506\,
            in3 => \N__40503\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46977\,
            in1 => \N__51450\,
            in2 => \_gnd_net_\,
            in3 => \N__43794\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52467\,
            lcout => \drone_H_disp_front_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59202\,
            ce => \N__50692\,
            sr => \N__57611\
        );

    \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__40689\,
            in1 => \N__42770\,
            in2 => \N__40662\,
            in3 => \N__42810\,
            lcout => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_6_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44704\,
            in1 => \N__40710\,
            in2 => \_gnd_net_\,
            in3 => \N__40698\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59217\,
            ce => \N__44612\,
            sr => \N__57618\
        );

    \ppm_encoder_1.pulses2count_esr_7_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40683\,
            in1 => \N__40674\,
            in2 => \_gnd_net_\,
            in3 => \N__44705\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59217\,
            ce => \N__44612\,
            sr => \N__57618\
        );

    \ppm_encoder_1.pulses2count_esr_13_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44703\,
            in1 => \N__40653\,
            in2 => \_gnd_net_\,
            in3 => \N__44346\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59217\,
            ce => \N__44612\,
            sr => \N__57618\
        );

    \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__42720\,
            in1 => \N__40644\,
            in2 => \N__41925\,
            in3 => \N__41769\,
            lcout => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_8_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44706\,
            in1 => \N__40638\,
            in2 => \_gnd_net_\,
            in3 => \N__46188\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59217\,
            ce => \N__44612\,
            sr => \N__57618\
        );

    \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__40626\,
            in1 => \N__44519\,
            in2 => \N__42696\,
            in3 => \N__40620\,
            lcout => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42076\,
            in1 => \N__42025\,
            in2 => \N__42057\,
            in3 => \N__43586\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_2_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__40800\,
            in1 => \_gnd_net_\,
            in2 => \N__44727\,
            in3 => \N__44301\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59234\,
            ce => \N__44592\,
            sr => \N__57625\
        );

    \ppm_encoder_1.pulses2count_esr_0_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44720\,
            in1 => \N__50214\,
            in2 => \_gnd_net_\,
            in3 => \N__40791\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59234\,
            ce => \N__44592\,
            sr => \N__57625\
        );

    \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__42075\,
            in1 => \N__40779\,
            in2 => \N__40773\,
            in3 => \N__44455\,
            lcout => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_1_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__44721\,
            in1 => \_gnd_net_\,
            in2 => \N__41562\,
            in3 => \N__43824\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59234\,
            ce => \N__44592\,
            sr => \N__57625\
        );

    \ppm_encoder_1.counter_0_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44459\,
            in2 => \N__40764\,
            in3 => \N__40763\,
            lcout => \ppm_encoder_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_0\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_1_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42078\,
            in2 => \_gnd_net_\,
            in3 => \N__40743\,
            lcout => \ppm_encoder_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_0\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_1\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_2_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42026\,
            in2 => \_gnd_net_\,
            in3 => \N__40740\,
            lcout => \ppm_encoder_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_1\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_2\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_3_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42056\,
            in2 => \_gnd_net_\,
            in3 => \N__40737\,
            lcout => \ppm_encoder_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_2\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_3\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_4_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42746\,
            in2 => \_gnd_net_\,
            in3 => \N__40734\,
            lcout => \ppm_encoder_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_3\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_4\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_5_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42789\,
            in2 => \_gnd_net_\,
            in3 => \N__40830\,
            lcout => \ppm_encoder_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_4\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_5\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_6_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42809\,
            in2 => \_gnd_net_\,
            in3 => \N__40827\,
            lcout => \ppm_encoder_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_5\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_6\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_7_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42769\,
            in2 => \_gnd_net_\,
            in3 => \N__40824\,
            lcout => \ppm_encoder_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_6\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_7\,
            clk => \N__59252\,
            ce => 'H',
            sr => \N__41046\
        );

    \ppm_encoder_1.counter_8_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42692\,
            in2 => \_gnd_net_\,
            in3 => \N__40821\,
            lcout => \ppm_encoder_1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_8\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_9_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44518\,
            in2 => \_gnd_net_\,
            in3 => \N__40818\,
            lcout => \ppm_encoder_1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_8\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_9\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_10_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44551\,
            in2 => \_gnd_net_\,
            in3 => \N__40815\,
            lcout => \ppm_encoder_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_9\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_10\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_11_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44491\,
            in2 => \_gnd_net_\,
            in3 => \N__40812\,
            lcout => \ppm_encoder_1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_10\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_11\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_12_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42719\,
            in2 => \_gnd_net_\,
            in3 => \N__40809\,
            lcout => \ppm_encoder_1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_11\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_12\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_13_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41921\,
            in2 => \_gnd_net_\,
            in3 => \N__40806\,
            lcout => \ppm_encoder_1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_12\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_13\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_14_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41945\,
            in2 => \_gnd_net_\,
            in3 => \N__40803\,
            lcout => \ppm_encoder_1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_13\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_14\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_15_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43103\,
            in2 => \_gnd_net_\,
            in3 => \N__41058\,
            lcout => \ppm_encoder_1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_14\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_15\,
            clk => \N__59267\,
            ce => 'H',
            sr => \N__41045\
        );

    \ppm_encoder_1.counter_16_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43143\,
            in2 => \_gnd_net_\,
            in3 => \N__41055\,
            lcout => \ppm_encoder_1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_16\,
            clk => \N__59279\,
            ce => 'H',
            sr => \N__41044\
        );

    \ppm_encoder_1.counter_17_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43124\,
            in2 => \_gnd_net_\,
            in3 => \N__41052\,
            lcout => \ppm_encoder_1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_16\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_17\,
            clk => \N__59279\,
            ce => 'H',
            sr => \N__41044\
        );

    \ppm_encoder_1.counter_18_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43158\,
            in2 => \_gnd_net_\,
            in3 => \N__41049\,
            lcout => \ppm_encoder_1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59279\,
            ce => 'H',
            sr => \N__41044\
        );

    \ppm_encoder_1.aileron_0_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__45405\,
            in1 => \N__43289\,
            in2 => \_gnd_net_\,
            in3 => \N__50233\,
            lcout => \ppm_encoder_1.aileronZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59099\,
            ce => 'H',
            sr => \N__57537\
        );

    \scaler_4.source_data_1_4_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__41021\,
            in1 => \N__41217\,
            in2 => \N__46817\,
            in3 => \N__41173\,
            lcout => scaler_4_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59106\,
            ce => 'H',
            sr => \N__57545\
        );

    \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40982\,
            in2 => \_gnd_net_\,
            in3 => \N__57842\,
            lcout => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__57843\,
            in1 => \N__41072\,
            in2 => \N__46353\,
            in3 => \N__48743\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46332\,
            in1 => \N__48330\,
            in2 => \_gnd_net_\,
            in3 => \N__40849\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46501\,
            in2 => \N__41088\,
            in3 => \N__46664\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__47172\,
            in1 => \N__43482\,
            in2 => \_gnd_net_\,
            in3 => \N__43351\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__47173\,
            in1 => \N__43483\,
            in2 => \_gnd_net_\,
            in3 => \N__43350\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001110"
        )
    port map (
            in0 => \N__48740\,
            in1 => \N__57887\,
            in2 => \N__49082\,
            in3 => \N__43485\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__57886\,
            in1 => \N__43409\,
            in2 => \N__43170\,
            in3 => \N__48742\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43316\,
            in2 => \_gnd_net_\,
            in3 => \N__43699\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__57885\,
            in1 => \N__43388\,
            in2 => \N__41073\,
            in3 => \N__48741\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIH72D6_12_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \N__46641\,
            in1 => \N__41085\,
            in2 => \_gnd_net_\,
            in3 => \N__41079\,
            lcout => \ppm_encoder_1.elevator_RNIH72D6Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__46352\,
            in1 => \N__47162\,
            in2 => \N__51448\,
            in3 => \N__49061\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__48739\,
            in1 => \N__57888\,
            in2 => \N__41262\,
            in3 => \N__41103\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__41259\,
            in1 => \N__41213\,
            in2 => \_gnd_net_\,
            in3 => \N__41175\,
            lcout => \scaler_4.un2_source_data_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.source_pid_1_esr_1_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__47745\,
            in1 => \N__44854\,
            in2 => \N__49695\,
            in3 => \N__45625\,
            lcout => side_order_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59135\,
            ce => \N__48036\,
            sr => \N__47994\
        );

    \pid_side.source_pid_1_esr_2_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__45626\,
            in1 => \N__49681\,
            in2 => \N__44859\,
            in3 => \N__49755\,
            lcout => side_order_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59135\,
            ce => \N__48036\,
            sr => \N__47994\
        );

    \pid_side.source_pid_1_esr_3_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__49728\,
            in1 => \N__44858\,
            in2 => \N__49696\,
            in3 => \N__45627\,
            lcout => side_order_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59135\,
            ce => \N__48036\,
            sr => \N__47994\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__43481\,
            in1 => \N__43692\,
            in2 => \N__43445\,
            in3 => \N__43517\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__43480\,
            in1 => \N__43436\,
            in2 => \N__48735\,
            in3 => \N__43691\,
            lcout => \ppm_encoder_1.init_pulses_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43410\,
            in3 => \N__41102\,
            lcout => \ppm_encoder_1.N_221\,
            ltout => \ppm_encoder_1.N_221_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48635\,
            in1 => \N__43479\,
            in2 => \N__41091\,
            in3 => \N__43435\,
            lcout => \ppm_encoder_1.init_pulses_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__41848\,
            in1 => \N__46952\,
            in2 => \N__45514\,
            in3 => \N__44123\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__41873\,
            in1 => \N__46800\,
            in2 => \N__41354\,
            in3 => \N__44048\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIFISN6_4_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__44424\,
            in1 => \_gnd_net_\,
            in2 => \N__41385\,
            in3 => \N__41382\,
            lcout => \ppm_encoder_1.elevator_RNIFISN6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__43189\,
            in1 => \N__51265\,
            in2 => \N__45515\,
            in3 => \N__44124\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__43357\,
            in1 => \N__43389\,
            in2 => \N__43317\,
            in3 => \N__48642\,
            lcout => \ppm_encoder_1.init_pulses_3_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__44049\,
            in1 => \N__43223\,
            in2 => \N__41376\,
            in3 => \N__45971\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIKNSN6_5_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46004\,
            in2 => \N__41373\,
            in3 => \N__41370\,
            lcout => \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI077O2_1_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__41461\,
            in1 => \N__41509\,
            in2 => \N__45545\,
            in3 => \N__44170\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIUINC6_1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \N__43845\,
            in1 => \N__41268\,
            in2 => \N__41364\,
            in3 => \N__41328\,
            lcout => \ppm_encoder_1.throttle_RNIUINC6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIEES71_1_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41410\,
            in1 => \N__43703\,
            in2 => \N__43809\,
            in3 => \N__48696\,
            lcout => \ppm_encoder_1.throttle_m_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47170\,
            in1 => \N__41462\,
            in2 => \_gnd_net_\,
            in3 => \N__41411\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51411\,
            in2 => \N__41565\,
            in3 => \N__41510\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_1_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__45376\,
            in1 => \N__41546\,
            in2 => \N__41526\,
            in3 => \N__41511\,
            lcout => \ppm_encoder_1.aileronZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59162\,
            ce => 'H',
            sr => \N__57586\
        );

    \ppm_encoder_1.elevator_1_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__41463\,
            in1 => \N__41496\,
            in2 => \N__41487\,
            in3 => \N__45380\,
            lcout => \ppm_encoder_1.elevatorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59162\,
            ce => 'H',
            sr => \N__57586\
        );

    \ppm_encoder_1.throttle_1_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__41451\,
            in1 => \N__41439\,
            in2 => \N__45403\,
            in3 => \N__41412\,
            lcout => \ppm_encoder_1.throttleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59162\,
            ce => 'H',
            sr => \N__57586\
        );

    \ppm_encoder_1.elevator_RNINSH16_0_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43638\,
            in2 => \N__46044\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43841\,
            in2 => \N__41400\,
            in3 => \N__41391\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44276\,
            in2 => \N__43758\,
            in3 => \N__41388\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44237\,
            in2 => \N__43968\,
            in3 => \N__41685\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44417\,
            in2 => \N__41682\,
            in3 => \N__41670\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46005\,
            in2 => \N__41667\,
            in3 => \N__41655\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45833\,
            in2 => \N__41652\,
            in3 => \N__41640\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45923\,
            in2 => \N__41637\,
            in3 => \N__41628\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46253\,
            in2 => \N__41625\,
            in3 => \N__41616\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_8\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46160\,
            in2 => \N__41613\,
            in3 => \N__41598\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46604\,
            in2 => \N__41595\,
            in3 => \N__41586\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47483\,
            in2 => \N__41583\,
            in3 => \N__41568\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46637\,
            in2 => \N__41757\,
            in3 => \N__41742\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44393\,
            in2 => \N__41739\,
            in3 => \N__41727\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44321\,
            in2 => \N__41724\,
            in3 => \N__41715\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45795\,
            in2 => \N__45816\,
            in3 => \N__41712\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43071\,
            in2 => \_gnd_net_\,
            in3 => \N__41709\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_16\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44259\,
            in2 => \_gnd_net_\,
            in3 => \N__41706\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41700\,
            in2 => \_gnd_net_\,
            in3 => \N__41703\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_2_18_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__48851\,
            in1 => \N__47883\,
            in2 => \N__49105\,
            in3 => \N__49074\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41694\,
            in2 => \_gnd_net_\,
            in3 => \N__43618\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47127\,
            in1 => \N__41877\,
            in2 => \_gnd_net_\,
            in3 => \N__41853\,
            lcout => \ppm_encoder_1.N_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__47109\,
            in1 => \N__57896\,
            in2 => \N__51449\,
            in3 => \N__48852\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_4_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__46092\,
            in1 => \N__44684\,
            in2 => \_gnd_net_\,
            in3 => \N__46932\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59218\,
            ce => \N__44602\,
            sr => \N__57619\
        );

    \ppm_encoder_1.pulses2count_esr_5_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44685\,
            in1 => \N__51246\,
            in2 => \_gnd_net_\,
            in3 => \N__45951\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59218\,
            ce => \N__44602\,
            sr => \N__57619\
        );

    \ppm_encoder_1.pulses2count_esr_10_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41829\,
            in1 => \N__47511\,
            in2 => \_gnd_net_\,
            in3 => \N__44681\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59218\,
            ce => \N__44602\,
            sr => \N__57619\
        );

    \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__44492\,
            in1 => \N__41823\,
            in2 => \N__41793\,
            in3 => \N__44552\,
            lcout => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_11_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41817\,
            in1 => \N__44682\,
            in2 => \_gnd_net_\,
            in3 => \N__41805\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59218\,
            ce => \N__44602\,
            sr => \N__57619\
        );

    \ppm_encoder_1.pulses2count_esr_12_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44683\,
            in1 => \N__41784\,
            in2 => \_gnd_net_\,
            in3 => \N__46653\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59218\,
            ce => \N__44602\,
            sr => \N__57619\
        );

    \ppm_encoder_1.counter24_0_I_1_c_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41763\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42003\,
            in2 => \N__42449\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_0\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41979\,
            in2 => \N__42439\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_1\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41901\,
            in2 => \N__42446\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_2\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41895\,
            in2 => \N__42440\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_3\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41889\,
            in2 => \N__42447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_4\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41883\,
            in2 => \N__42441\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_5\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42084\,
            in2 => \N__42448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_6\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42504\,
            in2 => \N__42450\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42468\,
            in2 => \N__42442\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_8\,
            carryout => \ppm_encoder_1.counter24_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42087\,
            lcout => \ppm_encoder_1.counter24_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__44733\,
            in1 => \N__43104\,
            in2 => \N__46869\,
            in3 => \N__41946\,
            lcout => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__43536\,
            in1 => \N__42052\,
            in2 => \N__42027\,
            in3 => \N__42077\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__42051\,
            in1 => \N__42033\,
            in2 => \N__44622\,
            in3 => \N__42021\,
            lcout => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__42787\,
            in1 => \N__41997\,
            in2 => \N__42747\,
            in3 => \N__41988\,
            lcout => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41973\,
            in1 => \N__44438\,
            in2 => \N__43083\,
            in3 => \N__42672\,
            lcout => \ppm_encoder_1.N_232\,
            ltout => \ppm_encoder_1.N_232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__44988\,
            in1 => \N__43608\,
            in2 => \N__41967\,
            in3 => \N__43537\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41944\,
            in2 => \_gnd_net_\,
            in3 => \N__41920\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIUS1G_4_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42808\,
            in1 => \N__42788\,
            in2 => \N__42771\,
            in3 => \N__42745\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIAEV01_8_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__42726\,
            in1 => \N__42718\,
            in2 => \N__42699\,
            in3 => \N__42691\,
            lcout => \ppm_encoder_1.N_139_17\,
            ltout => \ppm_encoder_1.N_139_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_1_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44439\,
            in1 => \N__42666\,
            in2 => \N__42657\,
            in3 => \N__43082\,
            lcout => \ppm_encoder_1.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_esr_RNIGKTC2_20_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42627\,
            in2 => \_gnd_net_\,
            in3 => \N__42561\,
            lcout => \pid_front.error_p_reg_esr_RNIGKTC2Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__42491\,
            in1 => \N__43120\,
            in2 => \N__45011\,
            in3 => \N__43141\,
            lcout => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_16_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__46907\,
            in1 => \N__44772\,
            in2 => \N__42495\,
            in3 => \N__48870\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59280\,
            ce => 'H',
            sr => \N__57640\
        );

    \ppm_encoder_1.pulses2count_18_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__48869\,
            in1 => \N__46908\,
            in2 => \N__42480\,
            in3 => \N__49113\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59280\,
            ce => 'H',
            sr => \N__57640\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42476\,
            in2 => \_gnd_net_\,
            in3 => \N__43156\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNI637H_18_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43157\,
            in1 => \N__43142\,
            in2 => \N__43128\,
            in3 => \N__43102\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49083\,
            in1 => \N__44771\,
            in2 => \_gnd_net_\,
            in3 => \N__48868\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_20_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59502\,
            lcout => \pid_front.error_d_reg_prevZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59289\,
            ce => \N__49368\,
            sr => \N__57644\
        );

    \pid_side.source_pid_1_10_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__47578\,
            in1 => \N__45695\,
            in2 => \N__43033\,
            in3 => \N__49967\,
            lcout => side_order_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59107\,
            ce => 'H',
            sr => \N__47986\
        );

    \pid_side.source_pid_1_11_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__45696\,
            in1 => \N__47579\,
            in2 => \N__43006\,
            in3 => \N__49928\,
            lcout => side_order_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59107\,
            ce => 'H',
            sr => \N__47986\
        );

    \pid_side.source_pid_1_6_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111010"
        )
    port map (
            in0 => \N__47580\,
            in1 => \N__49568\,
            in2 => \N__42961\,
            in3 => \N__45697\,
            lcout => side_order_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59107\,
            ce => 'H',
            sr => \N__47986\
        );

    \pid_side.source_pid_1_7_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__45698\,
            in1 => \N__49542\,
            in2 => \N__42916\,
            in3 => \N__47581\,
            lcout => side_order_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59107\,
            ce => 'H',
            sr => \N__47986\
        );

    \pid_side.source_pid_1_8_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__47582\,
            in1 => \N__45699\,
            in2 => \N__42871\,
            in3 => \N__49509\,
            lcout => side_order_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59107\,
            ce => 'H',
            sr => \N__47986\
        );

    \pid_side.source_pid_1_9_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__45700\,
            in1 => \N__47583\,
            in2 => \N__42835\,
            in3 => \N__49488\,
            lcout => side_order_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59107\,
            ce => 'H',
            sr => \N__47986\
        );

    \pid_side.state_RNID6CB8_1_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47577\,
            in2 => \_gnd_net_\,
            in3 => \N__47982\,
            lcout => \pid_side.state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.source_pid_1_esr_0_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__47769\,
            in1 => \N__44843\,
            in2 => \N__49697\,
            in3 => \N__45613\,
            lcout => side_order_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59114\,
            ce => \N__48020\,
            sr => \N__47983\
        );

    \pid_side.source_pid_1_esr_5_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__45643\,
            in1 => \N__45701\,
            in2 => \N__49619\,
            in3 => \N__45663\,
            lcout => side_order_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59114\,
            ce => \N__48020\,
            sr => \N__47983\
        );

    \pid_side.source_pid_1_esr_4_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__49698\,
            in1 => \N__45702\,
            in2 => \N__49620\,
            in3 => \N__45614\,
            lcout => side_order_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59124\,
            ce => \N__48021\,
            sr => \N__47987\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43437\,
            in1 => \N__45870\,
            in2 => \_gnd_net_\,
            in3 => \N__43668\,
            lcout => \ppm_encoder_1.N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47151\,
            in1 => \N__43227\,
            in2 => \_gnd_net_\,
            in3 => \N__43200\,
            lcout => \ppm_encoder_1.N_291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48274\,
            in2 => \_gnd_net_\,
            in3 => \N__48736\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010101010"
        )
    port map (
            in0 => \N__43355\,
            in1 => \N__47152\,
            in2 => \N__51432\,
            in3 => \N__46360\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__57889\,
            in1 => \N__43356\,
            in2 => \N__43161\,
            in3 => \N__48738\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59136\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43438\,
            in1 => \N__43387\,
            in2 => \N__43359\,
            in3 => \N__43484\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_153_d\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48275\,
            in2 => \N__43449\,
            in3 => \N__48737\,
            lcout => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__57890\,
            in1 => \N__51382\,
            in2 => \N__43446\,
            in3 => \N__48645\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43722\,
            in2 => \_gnd_net_\,
            in3 => \N__43743\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43382\,
            in2 => \_gnd_net_\,
            in3 => \N__43408\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001110"
        )
    port map (
            in0 => \N__43383\,
            in1 => \N__43358\,
            in2 => \N__43320\,
            in3 => \N__43312\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43296\,
            in3 => \N__48643\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010010"
        )
    port map (
            in0 => \N__48644\,
            in1 => \N__48994\,
            in2 => \N__43728\,
            in3 => \N__57894\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__43745\,
            in1 => \N__51381\,
            in2 => \N__57902\,
            in3 => \N__48646\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43744\,
            in2 => \_gnd_net_\,
            in3 => \N__43723\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__47000\,
            in1 => \N__43793\,
            in2 => \N__44159\,
            in3 => \N__44020\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001111"
        )
    port map (
            in0 => \N__45504\,
            in1 => \N__47039\,
            in2 => \N__43761\,
            in3 => \N__44280\,
            lcout => \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__43746\,
            in1 => \N__43724\,
            in2 => \N__43704\,
            in3 => \N__48636\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIGCMK2_0_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__43667\,
            in1 => \N__50240\,
            in2 => \N__43644\,
            in3 => \N__44126\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_0\,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__45879\,
            in1 => \N__46040\,
            in2 => \N__43641\,
            in3 => \N__45503\,
            lcout => \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43510\,
            in2 => \_gnd_net_\,
            in3 => \N__43573\,
            lcout => \ppm_encoder_1.PPM_STATE_53_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_1_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__43511\,
            in1 => \_gnd_net_\,
            in2 => \N__43560\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59163\,
            ce => 'H',
            sr => \N__57587\
        );

    \ppm_encoder_1.PPM_STATE_0_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__43628\,
            in1 => \N__43574\,
            in2 => \N__43539\,
            in3 => \N__43556\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59163\,
            ce => 'H',
            sr => \N__57587\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43865\,
            in1 => \N__47161\,
            in2 => \_gnd_net_\,
            in3 => \N__44226\,
            lcout => \ppm_encoder_1.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIMIMK2_3_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__44225\,
            in1 => \N__43915\,
            in2 => \N__44199\,
            in3 => \N__44021\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIT3R05_3_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__43864\,
            in1 => \N__44241\,
            in2 => \N__43971\,
            in3 => \N__45559\,
            lcout => \ppm_encoder_1.elevator_RNIT3R05Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51404\,
            in1 => \N__43959\,
            in2 => \_gnd_net_\,
            in3 => \N__43916\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_3_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__45381\,
            in1 => \N__43917\,
            in2 => \N__43953\,
            in3 => \N__43929\,
            lcout => \ppm_encoder_1.aileronZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59176\,
            ce => 'H',
            sr => \N__57598\
        );

    \ppm_encoder_1.elevator_3_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__43866\,
            in1 => \N__43902\,
            in2 => \N__45404\,
            in3 => \N__43890\,
            lcout => \ppm_encoder_1.elevatorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59176\,
            ce => 'H',
            sr => \N__57598\
        );

    \ppm_encoder_1.init_pulses_1_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__47277\,
            in1 => \N__47467\,
            in2 => \N__43854\,
            in3 => \N__48189\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59192\,
            ce => 'H',
            sr => \N__57605\
        );

    \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__47815\,
            in1 => \N__49025\,
            in2 => \_gnd_net_\,
            in3 => \N__48789\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001010101"
        )
    port map (
            in0 => \N__46684\,
            in1 => \N__46447\,
            in2 => \N__47822\,
            in3 => \N__46553\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__46448\,
            in1 => \N__45779\,
            in2 => \N__46572\,
            in3 => \N__46685\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_2_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47466\,
            in1 => \N__48153\,
            in2 => \N__47318\,
            in3 => \N__44286\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59192\,
            ce => 'H',
            sr => \N__57605\
        );

    \ppm_encoder_1.init_pulses_RNI87N01_2_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__45778\,
            in1 => \N__49026\,
            in2 => \_gnd_net_\,
            in3 => \N__48790\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000001111"
        )
    port map (
            in0 => \N__48236\,
            in1 => \N__46449\,
            in2 => \N__46689\,
            in3 => \N__46554\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_17_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47422\,
            in1 => \N__49128\,
            in2 => \N__47319\,
            in3 => \N__44265\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59204\,
            ce => 'H',
            sr => \N__57612\
        );

    \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__48794\,
            in1 => \N__45025\,
            in2 => \_gnd_net_\,
            in3 => \N__49078\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__49077\,
            in1 => \_gnd_net_\,
            in2 => \N__45032\,
            in3 => \N__48793\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_3_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__47327\,
            in1 => \N__48132\,
            in2 => \N__44253\,
            in3 => \N__47424\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59204\,
            ce => 'H',
            sr => \N__57612\
        );

    \ppm_encoder_1.init_pulses_RNI98N01_3_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49075\,
            in1 => \N__48232\,
            in2 => \_gnd_net_\,
            in3 => \N__48791\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_4_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47423\,
            in1 => \N__48111\,
            in2 => \N__47320\,
            in3 => \N__44430\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59204\,
            ce => 'H',
            sr => \N__57612\
        );

    \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__48792\,
            in1 => \N__46108\,
            in2 => \_gnd_net_\,
            in3 => \N__49076\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48291\,
            in2 => \_gnd_net_\,
            in3 => \N__48832\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_13_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47417\,
            in1 => \N__49233\,
            in2 => \N__47348\,
            in3 => \N__44406\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59219\,
            ce => 'H',
            sr => \N__57620\
        );

    \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49073\,
            in1 => \N__47836\,
            in2 => \_gnd_net_\,
            in3 => \N__48833\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_18_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47418\,
            in1 => \N__48519\,
            in2 => \N__47349\,
            in3 => \N__44382\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59219\,
            ce => 'H',
            sr => \N__57620\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__47837\,
            in1 => \N__46573\,
            in2 => \N__46453\,
            in3 => \N__44376\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_14_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47419\,
            in1 => \N__49206\,
            in2 => \N__47350\,
            in3 => \N__44334\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59235\,
            ce => 'H',
            sr => \N__57626\
        );

    \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__44830\,
            in1 => \_gnd_net_\,
            in2 => \N__48867\,
            in3 => \N__49069\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__49067\,
            in1 => \N__48834\,
            in2 => \_gnd_net_\,
            in3 => \N__44831\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__44832\,
            in1 => \N__46574\,
            in2 => \N__46454\,
            in3 => \N__44820\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_15_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47420\,
            in1 => \N__49182\,
            in2 => \N__47351\,
            in3 => \N__44787\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59235\,
            ce => 'H',
            sr => \N__57626\
        );

    \ppm_encoder_1.init_pulses_16_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47421\,
            in1 => \N__49155\,
            in2 => \N__47352\,
            in3 => \N__44778\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59235\,
            ce => 'H',
            sr => \N__57626\
        );

    \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__44765\,
            in1 => \_gnd_net_\,
            in2 => \N__48866\,
            in3 => \N__49068\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_14_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44751\,
            in1 => \N__44725\,
            in2 => \_gnd_net_\,
            in3 => \N__44739\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59253\,
            ce => \N__44580\,
            sr => \N__57632\
        );

    \ppm_encoder_1.pulses2count_esr_3_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44726\,
            in1 => \N__44640\,
            in2 => \_gnd_net_\,
            in3 => \N__44631\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59253\,
            ce => \N__44580\,
            sr => \N__57632\
        );

    \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57844\,
            in2 => \_gnd_net_\,
            in3 => \N__48853\,
            lcout => \ppm_encoder_1.N_2150_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIK1KG_0_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__44553\,
            in1 => \N__44523\,
            in2 => \N__44496\,
            in3 => \N__44463\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_14_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59458\,
            lcout => \pid_front.error_d_reg_prevZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59281\,
            ce => \N__49374\,
            sr => \N__57641\
        );

    \ppm_encoder_1.pulses2count_17_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__45033\,
            in1 => \N__46900\,
            in2 => \N__45012\,
            in3 => \N__48871\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59290\,
            ce => 'H',
            sr => \N__57645\
        );

    \pid_side.pid_prereg_esr_RNIOPAK1_2_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__49748\,
            in1 => \N__47731\,
            in2 => \N__49724\,
            in3 => \N__47761\,
            lcout => \pid_side.m32_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIKRVH2_5_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__44994\,
            in1 => \N__47552\,
            in2 => \N__49618\,
            in3 => \N__44980\,
            lcout => \pid_side.un1_reset_0_i_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNI2NBO1_6_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__49564\,
            in1 => \N__49486\,
            in2 => \N__49541\,
            in3 => \N__49507\,
            lcout => \pid_side.m26_e_5\,
            ltout => \pid_side.m26_e_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNI7JSP1_10_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__49927\,
            in1 => \_gnd_net_\,
            in2 => \N__44865\,
            in3 => \N__49966\,
            lcout => \pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNI2NBO1_0_6_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__49487\,
            in1 => \N__49537\,
            in2 => \N__49569\,
            in3 => \N__49508\,
            lcout => \pid_side.m18_s_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIQEI8_13_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__50014\,
            in1 => \N__49854\,
            in2 => \_gnd_net_\,
            in3 => \N__48084\,
            lcout => \pid_side.N_11_0\,
            ltout => \pid_side.N_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNILRSP2_5_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49611\,
            in1 => \N__45645\,
            in2 => \N__44862\,
            in3 => \N__45694\,
            lcout => \pid_side.pid_prereg_esr_RNILRSP2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIGJDR1_10_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__49929\,
            in1 => \N__49968\,
            in2 => \N__45735\,
            in3 => \N__47517\,
            lcout => OPEN,
            ltout => \pid_side.pid_prereg_esr_RNIGJDR1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIQBAH2_23_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__48085\,
            in1 => \N__49664\,
            in2 => \N__45726\,
            in3 => \N__50015\,
            lcout => OPEN,
            ltout => \pid_side.pid_prereg_esr_RNIQBAH2Z0Z_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIKNK25_10_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__47592\,
            in1 => \N__45723\,
            in2 => \N__45717\,
            in3 => \N__45661\,
            lcout => OPEN,
            ltout => \pid_side.i19_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIKC058_23_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45714\,
            in2 => \N__45705\,
            in3 => \N__47523\,
            lcout => \pid_side.un1_reset_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIEUA9_12_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__50016\,
            in1 => \N__49855\,
            in2 => \N__49893\,
            in3 => \N__48086\,
            lcout => \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12\,
            ltout => \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIF0QB2_10_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__45662\,
            in1 => \_gnd_net_\,
            in2 => \N__45648\,
            in3 => \N__45644\,
            lcout => \pid_side.N_82_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.source_pid_1_esr_12_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__49857\,
            in1 => \N__48087\,
            in2 => \N__50028\,
            in3 => \N__49892\,
            lcout => side_order_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59137\,
            ce => \N__48025\,
            sr => \N__47984\
        );

    \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001100110"
        )
    port map (
            in0 => \N__45570\,
            in1 => \N__46036\,
            in2 => \N__45878\,
            in3 => \N__45557\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_0_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__45429\,
            in1 => \N__45385\,
            in2 => \_gnd_net_\,
            in3 => \N__45874\,
            lcout => \ppm_encoder_1.elevatorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59151\,
            ce => 'H',
            sr => \N__57579\
        );

    \ppm_encoder_1.init_pulses_6_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47468\,
            in1 => \N__48465\,
            in2 => \N__47315\,
            in3 => \N__45849\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59151\,
            ce => 'H',
            sr => \N__57579\
        );

    \ppm_encoder_1.init_pulses_RNICBN01_6_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__45751\,
            in1 => \N__48990\,
            in2 => \_gnd_net_\,
            in3 => \N__48797\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__48798\,
            in1 => \_gnd_net_\,
            in2 => \N__49043\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48931\,
            in2 => \_gnd_net_\,
            in3 => \N__48637\,
            lcout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\,
            ltout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNILVE13_0_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__48640\,
            in1 => \N__46063\,
            in2 => \N__45798\,
            in3 => \N__48286\,
            lcout => \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47871\,
            in1 => \N__48935\,
            in2 => \N__48864\,
            in3 => \N__47912\,
            lcout => \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__48641\,
            in1 => \N__45783\,
            in2 => \N__48296\,
            in3 => \N__47869\,
            lcout => \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47870\,
            in1 => \N__48290\,
            in2 => \N__48865\,
            in3 => \N__45752\,
            lcout => \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__48639\,
            in1 => \N__48285\,
            in2 => \N__46071\,
            in3 => \N__47872\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_0_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__47241\,
            in1 => \N__46080\,
            in2 => \N__46074\,
            in3 => \N__47469\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59164\,
            ce => 'H',
            sr => \N__57588\
        );

    \ppm_encoder_1.init_pulses_RNI65N01_0_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__48638\,
            in1 => \_gnd_net_\,
            in2 => \N__48995\,
            in3 => \N__46062\,
            lcout => \ppm_encoder_1.un1_init_pulses_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_5_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47456\,
            in1 => \N__48495\,
            in2 => \N__47316\,
            in3 => \N__46017\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59177\,
            ce => 'H',
            sr => \N__57599\
        );

    \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__48986\,
            in1 => \N__45983\,
            in2 => \_gnd_net_\,
            in3 => \N__48702\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__45982\,
            in1 => \_gnd_net_\,
            in2 => \N__48795\,
            in3 => \N__48987\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__46575\,
            in1 => \N__45984\,
            in2 => \N__46446\,
            in3 => \N__45972\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_7_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47457\,
            in1 => \N__48441\,
            in2 => \N__47317\,
            in3 => \N__45936\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59177\,
            ce => 'H',
            sr => \N__57599\
        );

    \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__48989\,
            in1 => \N__48709\,
            in2 => \_gnd_net_\,
            in3 => \N__45892\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__45893\,
            in1 => \_gnd_net_\,
            in2 => \N__48796\,
            in3 => \N__48988\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_8_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47461\,
            in1 => \N__48423\,
            in2 => \N__47346\,
            in3 => \N__46269\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59193\,
            ce => 'H',
            sr => \N__57606\
        );

    \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__46198\,
            in1 => \N__49021\,
            in2 => \_gnd_net_\,
            in3 => \N__48700\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__48698\,
            in1 => \_gnd_net_\,
            in2 => \N__49065\,
            in3 => \N__46199\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__46236\,
            in1 => \N__46436\,
            in2 => \N__46203\,
            in3 => \N__46564\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_9_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__47462\,
            in1 => \N__48408\,
            in2 => \N__47347\,
            in3 => \N__46173\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59193\,
            ce => 'H',
            sr => \N__57606\
        );

    \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__46127\,
            in1 => \N__49022\,
            in2 => \_gnd_net_\,
            in3 => \N__48701\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__48699\,
            in1 => \_gnd_net_\,
            in2 => \N__49066\,
            in3 => \N__46126\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__46113\,
            in1 => \N__49014\,
            in2 => \_gnd_net_\,
            in3 => \N__48697\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__46567\,
            in1 => \N__46112\,
            in2 => \N__46437\,
            in3 => \N__46796\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_4_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46824\,
            lcout => \ppm_encoder_1.rudderZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59205\,
            ce => \N__46781\,
            sr => \N__57613\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46407\,
            in1 => \N__47190\,
            in2 => \_gnd_net_\,
            in3 => \N__46716\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46568\,
            in2 => \N__46692\,
            in3 => \N__46676\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__49023\,
            in1 => \N__48815\,
            in2 => \_gnd_net_\,
            in3 => \N__47189\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101001101010"
        )
    port map (
            in0 => \N__47188\,
            in1 => \N__49024\,
            in2 => \N__48863\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_10_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__47343\,
            in1 => \N__47464\,
            in2 => \N__48390\,
            in3 => \N__46617\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59220\,
            ce => 'H',
            sr => \N__57621\
        );

    \ppm_encoder_1.init_pulses_RNINSJT_10_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__46585\,
            in1 => \_gnd_net_\,
            in2 => \N__48861\,
            in3 => \N__49080\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__49079\,
            in1 => \N__48808\,
            in2 => \_gnd_net_\,
            in3 => \N__46586\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__46587\,
            in1 => \N__46571\,
            in2 => \N__46455\,
            in3 => \N__46301\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_11_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__47344\,
            in1 => \N__47465\,
            in2 => \N__48366\,
            in3 => \N__47499\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59220\,
            ce => 'H',
            sr => \N__57621\
        );

    \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__48313\,
            in1 => \_gnd_net_\,
            in2 => \N__48862\,
            in3 => \N__49081\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_12_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__47463\,
            in1 => \N__47345\,
            in2 => \N__48345\,
            in3 => \N__47199\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59220\,
            ce => 'H',
            sr => \N__57621\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47126\,
            in1 => \N__47040\,
            in2 => \_gnd_net_\,
            in3 => \N__47004\,
            lcout => \ppm_encoder_1.N_288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51427\,
            in1 => \N__46968\,
            in2 => \_gnd_net_\,
            in3 => \N__46959\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_prev_esr_1_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56895\,
            lcout => \pid_front.error_d_reg_prevZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59268\,
            ce => \N__49376\,
            sr => \N__57637\
        );

    \ppm_encoder_1.pulses2count_15_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__47905\,
            in1 => \N__46865\,
            in2 => \N__46906\,
            in3 => \N__48873\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59282\,
            ce => 'H',
            sr => \N__57642\
        );

    \pid_front.error_d_reg_prev_esr_11_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56822\,
            lcout => \pid_front.error_d_reg_prevZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59291\,
            ce => \N__49375\,
            sr => \N__57646\
        );

    \pid_alt.state_RNICP2N1_0_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47796\,
            in2 => \_gnd_net_\,
            in3 => \N__58319\,
            lcout => \pid_alt.N_664_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_0_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__47618\,
            in1 => \N__50940\,
            in2 => \N__53511\,
            in3 => \N__47762\,
            lcout => \pid_side.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59115\,
            ce => 'H',
            sr => \N__57555\
        );

    \pid_side.pid_prereg_1_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__49266\,
            in1 => \N__50832\,
            in2 => \N__47741\,
            in3 => \N__47619\,
            lcout => \pid_side.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59115\,
            ce => 'H',
            sr => \N__57555\
        );

    \pid_side.state_0_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__47711\,
            in1 => \N__47617\,
            in2 => \_gnd_net_\,
            in3 => \N__47554\,
            lcout => \pid_side.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59115\,
            ce => 'H',
            sr => \N__57555\
        );

    \pid_side.state_RNINK4U_0_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__47553\,
            in1 => \N__47710\,
            in2 => \N__47622\,
            in3 => \N__57830\,
            lcout => \pid_side.state_RNINK4UZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.state_1_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59115\,
            ce => 'H',
            sr => \N__57555\
        );

    \pid_side.pid_prereg_esr_RNIU5CG_10_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__49926\,
            in1 => \N__49965\,
            in2 => \N__49694\,
            in3 => \N__49882\,
            lcout => \pid_side.m18_s_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNICPBG_23_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__57829\,
            in1 => \N__47551\,
            in2 => \_gnd_net_\,
            in3 => \N__50024\,
            lcout => \pid_side.un1_reset_0_i_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNI90H1_12_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49881\,
            in2 => \_gnd_net_\,
            in3 => \N__49842\,
            lcout => \pid_side.m26_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNI2MA2_14_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__49821\,
            in1 => \N__50046\,
            in2 => \_gnd_net_\,
            in3 => \N__49806\,
            lcout => \pid_side.m9_e_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50085\,
            in1 => \N__49794\,
            in2 => \N__49770\,
            in3 => \N__49782\,
            lcout => OPEN,
            ltout => \pid_side.m9_e_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIFB07_20_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__48096\,
            in1 => \N__50070\,
            in2 => \N__48090\,
            in3 => \N__50058\,
            lcout => \pid_side.pid_prereg_esr_RNIFB07Z0Z_20\,
            ltout => \pid_side.pid_prereg_esr_RNIFB07Z0Z_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.source_pid_1_esr_13_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__50020\,
            in1 => \_gnd_net_\,
            in2 => \N__48069\,
            in3 => \N__49856\,
            lcout => side_order_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59138\,
            ce => \N__48035\,
            sr => \N__47985\
        );

    \Commands_frame_decoder.state_RNIC08S_3_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47945\,
            in2 => \_gnd_net_\,
            in3 => \N__57858\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__47913\,
            in1 => \N__48999\,
            in2 => \_gnd_net_\,
            in3 => \N__48823\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__48825\,
            in1 => \N__47873\,
            in2 => \N__48297\,
            in3 => \N__47847\,
            lcout => \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__47823\,
            in1 => \N__48996\,
            in2 => \_gnd_net_\,
            in3 => \N__48819\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011011110"
        )
    port map (
            in0 => \N__48824\,
            in1 => \N__57895\,
            in2 => \N__51400\,
            in3 => \N__49013\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__48326\,
            in1 => \N__48998\,
            in2 => \_gnd_net_\,
            in3 => \N__48821\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48822\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48292\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__48240\,
            in1 => \N__48997\,
            in2 => \_gnd_net_\,
            in3 => \N__48820\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48216\,
            in2 => \N__48204\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48195\,
            in2 => \_gnd_net_\,
            in3 => \N__48177\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48174\,
            in2 => \N__48168\,
            in3 => \N__48141\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48138\,
            in2 => \_gnd_net_\,
            in3 => \N__48120\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48117\,
            in2 => \_gnd_net_\,
            in3 => \N__48099\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48501\,
            in2 => \_gnd_net_\,
            in3 => \N__48489\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48486\,
            in2 => \N__48480\,
            in3 => \N__48453\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48450\,
            in3 => \N__48435\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48432\,
            in2 => \_gnd_net_\,
            in3 => \N__48417\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_8\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48414\,
            in2 => \_gnd_net_\,
            in3 => \N__48402\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48399\,
            in2 => \_gnd_net_\,
            in3 => \N__48378\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48375\,
            in2 => \_gnd_net_\,
            in3 => \N__48354\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48351\,
            in2 => \_gnd_net_\,
            in3 => \N__48333\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49254\,
            in2 => \N__49245\,
            in3 => \N__49221\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49218\,
            in2 => \_gnd_net_\,
            in3 => \N__49194\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49191\,
            in2 => \_gnd_net_\,
            in3 => \N__49170\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49167\,
            in2 => \_gnd_net_\,
            in3 => \N__49143\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_16\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49140\,
            in2 => \_gnd_net_\,
            in3 => \N__49116\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__49112\,
            in1 => \N__49060\,
            in2 => \N__48872\,
            in3 => \N__48522\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48507\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \drone_H_disp_side_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52484\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59236\,
            ce => \N__50297\,
            sr => \N__57627\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53224\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59236\,
            ce => \N__50297\,
            sr => \N__57627\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52374\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59236\,
            ce => \N__50297\,
            sr => \N__57627\
        );

    \pid_front.pid_prereg_0_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__50508\,
            in1 => \N__49461\,
            in2 => \N__56940\,
            in3 => \N__49423\,
            lcout => \pid_front.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59269\,
            ce => 'H',
            sr => \N__57638\
        );

    \pid_front.error_d_reg_prev_esr_18_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59573\,
            lcout => \pid_front.error_d_reg_prevZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59292\,
            ce => \N__49377\,
            sr => \N__57647\
        );

    \pid_front.error_d_reg_esr_2_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49311\,
            lcout => \pid_front.error_d_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59302\,
            ce => \N__58455\,
            sr => \N__58179\
        );

    \GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57827\,
            lcout => \GB_BUFFER_reset_system_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_1_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53436\,
            lcout => \pid_side.error_d_reg_prevZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59125\,
            ce => \N__57948\,
            sr => \N__57564\
        );

    \pid_side.error_d_reg_prev_esr_0_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50936\,
            in2 => \N__53510\,
            in3 => \N__53509\,
            lcout => \pid_side.error_d_reg_prevZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_20_9_0_\,
            carryout => \pid_side.un1_pid_prereg_cry_0\,
            clk => \N__59140\,
            ce => \N__57950\,
            sr => \N__57574\
        );

    \pid_side.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50828\,
            in2 => \_gnd_net_\,
            in3 => \N__49257\,
            lcout => \pid_side.un1_pid_prereg_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_0\,
            carryout => \pid_side.un1_pid_prereg_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_2_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50814\,
            in2 => \N__50967\,
            in3 => \N__49731\,
            lcout => \pid_side.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_1\,
            carryout => \pid_side.un1_pid_prereg_cry_0_0\,
            clk => \N__59140\,
            ce => \N__57950\,
            sr => \N__57574\
        );

    \pid_side.pid_prereg_esr_3_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50925\,
            in2 => \N__53043\,
            in3 => \N__49701\,
            lcout => \pid_side.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_0_0\,
            carryout => \pid_side.un1_pid_prereg_cry_1_0\,
            clk => \N__59140\,
            ce => \N__57950\,
            sr => \N__57574\
        );

    \pid_side.pid_prereg_esr_4_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53655\,
            in2 => \N__52803\,
            in3 => \N__49623\,
            lcout => \pid_side.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_1_0\,
            carryout => \pid_side.un1_pid_prereg_cry_2\,
            clk => \N__59140\,
            ce => \N__57950\,
            sr => \N__57574\
        );

    \pid_side.pid_prereg_esr_5_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52833\,
            in2 => \N__52857\,
            in3 => \N__49572\,
            lcout => \pid_side.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_2\,
            carryout => \pid_side.un1_pid_prereg_cry_3\,
            clk => \N__59140\,
            ce => \N__57950\,
            sr => \N__57574\
        );

    \pid_side.pid_prereg_esr_6_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52877\,
            in2 => \N__50847\,
            in3 => \N__49545\,
            lcout => \pid_side.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_3\,
            carryout => \pid_side.un1_pid_prereg_cry_4\,
            clk => \N__59140\,
            ce => \N__57950\,
            sr => \N__57574\
        );

    \pid_side.pid_prereg_esr_7_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54633\,
            in2 => \N__54612\,
            in3 => \N__49512\,
            lcout => \pid_side.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_4\,
            carryout => \pid_side.un1_pid_prereg_cry_5\,
            clk => \N__59140\,
            ce => \N__57950\,
            sr => \N__57574\
        );

    \pid_side.pid_prereg_esr_8_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54942\,
            in2 => \N__54591\,
            in3 => \N__49491\,
            lcout => \pid_side.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_20_10_0_\,
            carryout => \pid_side.un1_pid_prereg_cry_6\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_9_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53703\,
            in2 => \N__53727\,
            in3 => \N__49464\,
            lcout => \pid_side.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_6\,
            carryout => \pid_side.un1_pid_prereg_cry_7\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_10_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51078\,
            in2 => \N__53757\,
            in3 => \N__49932\,
            lcout => \pid_side.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_7\,
            carryout => \pid_side.un1_pid_prereg_cry_8\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_11_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51063\,
            in2 => \N__51183\,
            in3 => \N__49896\,
            lcout => \pid_side.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_8\,
            carryout => \pid_side.un1_pid_prereg_cry_9\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_12_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51195\,
            in2 => \N__51135\,
            in3 => \N__49860\,
            lcout => \pid_side.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_9\,
            carryout => \pid_side.un1_pid_prereg_cry_10\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_13_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51102\,
            in2 => \N__51122\,
            in3 => \N__49824\,
            lcout => \pid_side.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_10\,
            carryout => \pid_side.un1_pid_prereg_cry_11\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_14_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51093\,
            in2 => \N__51003\,
            in3 => \N__49809\,
            lcout => \pid_side.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_11\,
            carryout => \pid_side.un1_pid_prereg_cry_12\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_15_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51057\,
            in2 => \N__50916\,
            in3 => \N__49797\,
            lcout => \pid_side.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_12\,
            carryout => \pid_side.un1_pid_prereg_cry_13\,
            clk => \N__59153\,
            ce => \N__57951\,
            sr => \N__57581\
        );

    \pid_side.pid_prereg_esr_16_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51084\,
            in2 => \N__50181\,
            in3 => \N__49785\,
            lcout => \pid_side.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_20_11_0_\,
            carryout => \pid_side.un1_pid_prereg_cry_14\,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.pid_prereg_esr_17_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49974\,
            in2 => \N__50106\,
            in3 => \N__49773\,
            lcout => \pid_side.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_14\,
            carryout => \pid_side.un1_pid_prereg_cry_15\,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.pid_prereg_esr_18_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50157\,
            in2 => \N__52923\,
            in3 => \N__49758\,
            lcout => \pid_side.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_15\,
            carryout => \pid_side.un1_pid_prereg_cry_16\,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.pid_prereg_esr_19_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50172\,
            in2 => \N__53553\,
            in3 => \N__50073\,
            lcout => \pid_side.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_16\,
            carryout => \pid_side.un1_pid_prereg_cry_17\,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.pid_prereg_esr_20_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49980\,
            in2 => \N__50166\,
            in3 => \N__50061\,
            lcout => \pid_side.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_17\,
            carryout => \pid_side.un1_pid_prereg_cry_18\,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.pid_prereg_esr_21_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50094\,
            in2 => \N__50196\,
            in3 => \N__50049\,
            lcout => \pid_side.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_18\,
            carryout => \pid_side.un1_pid_prereg_cry_19\,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.pid_prereg_esr_22_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50274\,
            in2 => \N__51204\,
            in3 => \N__50034\,
            lcout => \pid_side.pid_preregZ0Z_22\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_19\,
            carryout => \pid_side.un1_pid_prereg_cry_20\,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.pid_prereg_esr_23_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50265\,
            in2 => \_gnd_net_\,
            in3 => \N__50031\,
            lcout => \pid_side.pid_preregZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59166\,
            ce => \N__57952\,
            sr => \N__57590\
        );

    \pid_side.error_d_reg_prev_esr_RNILHF23_18_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__51833\,
            in1 => \N__51227\,
            in2 => \N__53991\,
            in3 => \N__52956\,
            lcout => \pid_side.error_d_reg_prev_esr_RNILHF23Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIJV5H1_15_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50117\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIJV5H1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54378\,
            in1 => \N__52989\,
            in2 => \_gnd_net_\,
            in3 => \N__54813\,
            lcout => \pid_side.un1_pid_prereg_30\,
            ltout => \pid_side.un1_pid_prereg_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI0PB23_14_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__50135\,
            in1 => \N__50994\,
            in2 => \N__50184\,
            in3 => \N__52974\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI0PB23Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI4UC23_17_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__52896\,
            in1 => \N__52954\,
            in2 => \N__51228\,
            in3 => \N__54102\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI4UC23Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI5I6H1_18_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51226\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI5I6H1Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIP56H1_16_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__54121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52934\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIP56H1Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_16_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59195\,
            ce => \N__57956\,
            sr => \N__57607\
        );

    \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54179\,
            in1 => \N__50144\,
            in2 => \_gnd_net_\,
            in3 => \N__56626\,
            lcout => \pid_side.un1_pid_prereg_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__56627\,
            in1 => \_gnd_net_\,
            in2 => \N__50148\,
            in3 => \N__54180\,
            lcout => \pid_side.un1_pid_prereg_36\,
            ltout => \pid_side.un1_pid_prereg_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIC5C23_15_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__54122\,
            in1 => \N__50136\,
            in2 => \N__50121\,
            in3 => \N__50118\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIC5C23Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI89K23_19_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__54029\,
            in1 => \N__53983\,
            in2 => \N__51834\,
            in3 => \N__53980\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI89K23Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIGJM23_20_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__54028\,
            in1 => \N__53979\,
            in2 => \N__54035\,
            in3 => \N__53978\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIGJM23Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNO_0_23_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__54030\,
            in1 => \N__53981\,
            in2 => \N__54036\,
            in3 => \N__53982\,
            lcout => \pid_side.un1_pid_prereg_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51365\,
            in1 => \N__50256\,
            in2 => \_gnd_net_\,
            in3 => \N__50244\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIGV8H1_19_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53974\,
            in2 => \_gnd_net_\,
            in3 => \N__51826\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIGV8H1Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH2data_esr_1_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56285\,
            lcout => side_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59238\,
            ce => \N__51810\,
            sr => \N__57628\
        );

    \Commands_frame_decoder.source_CH2data_esr_2_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56132\,
            lcout => side_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59238\,
            ce => \N__51810\,
            sr => \N__57628\
        );

    \Commands_frame_decoder.source_CH2data_esr_0_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56507\,
            lcout => side_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59238\,
            ce => \N__51810\,
            sr => \N__57628\
        );

    \Commands_frame_decoder.source_CH2data_esr_4_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53397\,
            lcout => side_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59238\,
            ce => \N__51810\,
            sr => \N__57628\
        );

    \Commands_frame_decoder.source_CH2data_esr_5_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55926\,
            lcout => side_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59238\,
            ce => \N__51810\,
            sr => \N__57628\
        );

    \Commands_frame_decoder.source_CH2data_esr_6_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__55749\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => side_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59238\,
            ce => \N__51810\,
            sr => \N__57628\
        );

    \Commands_frame_decoder.source_CH2data_ess_7_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55574\,
            lcout => side_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59238\,
            ce => \N__51810\,
            sr => \N__57628\
        );

    \pid_side.error_axb_1_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50409\,
            lcout => \pid_side.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50780\,
            lcout => \drone_H_disp_side_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59254\,
            ce => \N__50298\,
            sr => \N__57633\
        );

    \pid_side.error_axb_2_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50310\,
            lcout => \pid_side.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50402\,
            lcout => \drone_H_disp_side_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59254\,
            ce => \N__50298\,
            sr => \N__57633\
        );

    \pid_side.error_axb_3_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50304\,
            lcout => \pid_side.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52709\,
            lcout => \drone_H_disp_side_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59254\,
            ce => \N__50298\,
            sr => \N__57633\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52307\,
            lcout => \drone_H_disp_side_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59254\,
            ce => \N__50298\,
            sr => \N__57633\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52605\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59254\,
            ce => \N__50298\,
            sr => \N__57633\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50703\,
            lcout => \drone_H_disp_front_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50781\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59271\,
            ce => \N__50696\,
            sr => \N__57639\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52406\,
            lcout => \drone_H_disp_side_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50649\,
            lcout => \drone_H_disp_side_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50643\,
            lcout => \drone_H_disp_side_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50634\,
            lcout => \drone_H_disp_side_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52236\,
            lcout => \drone_H_disp_side_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.state_1_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50505\,
            lcout => \pid_front.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59284\,
            ce => 'H',
            sr => \N__57643\
        );

    \pid_front.pid_prereg_1_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__50544\,
            in1 => \N__50529\,
            in2 => \N__50434\,
            in3 => \N__50506\,
            lcout => \pid_front.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59284\,
            ce => 'H',
            sr => \N__57643\
        );

    \pid_side.error_axb_8_l_ofx_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__52614\,
            in1 => \_gnd_net_\,
            in2 => \N__50892\,
            in3 => \N__52502\,
            lcout => \pid_side.error_axb_8_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_axb_7_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50888\,
            in2 => \_gnd_net_\,
            in3 => \N__52613\,
            lcout => \pid_side.error_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52501\,
            lcout => \drone_H_disp_side_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_3_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50877\,
            lcout => \pid_front.error_d_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59315\,
            ce => \N__58494\,
            sr => \N__58180\
        );

    \pid_side.error_p_reg_esr_RNI5QI23_5_LC_21_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100100111001"
        )
    port map (
            in0 => \N__53784\,
            in1 => \N__54894\,
            in2 => \N__53823\,
            in3 => \N__52878\,
            lcout => \pid_side.error_p_reg_esr_RNI5QI23Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_5_LC_21_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54753\,
            lcout => \pid_side.error_d_reg_prevZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59126\,
            ce => \N__57949\,
            sr => \N__57565\
        );

    \pid_side.error_d_reg_esr_RNI5QKD1_1_LC_21_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__53022\,
            in1 => \N__50952\,
            in2 => \N__53435\,
            in3 => \N__50807\,
            lcout => \pid_side.un1_pid_prereg_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNISH6J_0_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__50950\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53020\,
            lcout => OPEN,
            ltout => \pid_side.error_p_reg_esr_RNISH6JZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNIFP9R2_1_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011111010"
        )
    port map (
            in0 => \N__53431\,
            in1 => \N__50966\,
            in2 => \N__50817\,
            in3 => \N__50808\,
            lcout => \pid_side.error_d_reg_esr_RNIFP9R2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIUJ6J_0_1_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54257\,
            in2 => \_gnd_net_\,
            in3 => \N__50978\,
            lcout => \pid_side.N_1546_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIUJ6J_1_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__50979\,
            in1 => \_gnd_net_\,
            in2 => \N__54261\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1\,
            ltout => \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIAVKD1_0_1_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53645\,
            in2 => \N__50970\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.un1_pid_prereg\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNISH6J_0_0_LC_21_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__53021\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50951\,
            lcout => \pid_side.un1_pid_prereg_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIAVKD1_1_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53646\,
            in2 => \_gnd_net_\,
            in3 => \N__53054\,
            lcout => \pid_side.error_p_reg_esr_RNIAVKD1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54512\,
            in1 => \N__50900\,
            in2 => \_gnd_net_\,
            in3 => \N__55102\,
            lcout => \pid_side.un1_pid_prereg_18\,
            ltout => \pid_side.un1_pid_prereg_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50919\,
            in3 => \N__51048\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54513\,
            in1 => \N__50901\,
            in2 => \_gnd_net_\,
            in3 => \N__55103\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13\,
            ltout => \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI4NA21_0_12_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50904\,
            in3 => \N__51523\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_13_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55104\,
            lcout => \pid_side.error_d_reg_prevZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59167\,
            ce => \N__57953\,
            sr => \N__57591\
        );

    \pid_side.error_d_reg_prev_esr_RNI4NA21_12_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51026\,
            in2 => \_gnd_net_\,
            in3 => \N__51524\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI4NA21Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54431\,
            in1 => \N__53574\,
            in2 => \_gnd_net_\,
            in3 => \N__55169\,
            lcout => \pid_side.un1_pid_prereg_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIDP5H1_14_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50993\,
            in2 => \_gnd_net_\,
            in3 => \N__52970\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIDP5H1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNIKMFP2_10_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__55078\,
            in1 => \N__51072\,
            in2 => \N__53756\,
            in3 => \N__52997\,
            lcout => \pid_side.error_d_reg_esr_RNIKMFP2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIUQN9_0_10_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54401\,
            in2 => \_gnd_net_\,
            in3 => \N__53538\,
            lcout => \pid_side.N_1582_i\,
            ltout => \pid_side.N_1582_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNI104E2_10_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__55079\,
            in1 => \N__51179\,
            in2 => \N__51066\,
            in3 => \N__52998\,
            lcout => \pid_side.error_d_reg_esr_RNI104E2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIKCB23_13_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__51047\,
            in1 => \N__50992\,
            in2 => \N__51015\,
            in3 => \N__52969\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIKCB23Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIBAGJ2_12_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__51525\,
            in1 => \N__51046\,
            in2 => \N__51033\,
            in3 => \N__51011\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIBAGJ2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54377\,
            in1 => \N__52985\,
            in2 => \_gnd_net_\,
            in3 => \N__54808\,
            lcout => \pid_side.un1_pid_prereg_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIO9BH1_20_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53990\,
            in2 => \_gnd_net_\,
            in3 => \N__54034\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIO9BH1Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNILJFJ2_12_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51548\,
            in1 => \N__51144\,
            in2 => \N__51165\,
            in3 => \N__51555\,
            lcout => \pid_side.error_d_reg_prev_esr_RNILJFJ2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIUQN9_10_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__53537\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54405\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10\,
            ltout => \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIQCA21_0_10_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51186\,
            in3 => \N__51158\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__51506\,
            in1 => \N__51483\,
            in2 => \_gnd_net_\,
            in3 => \N__54870\,
            lcout => \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11\,
            ltout => \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIQCA21_10_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51147\,
            in3 => \N__51143\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIQCA21Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_12_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54711\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59207\,
            ce => \N__57958\,
            sr => \N__57614\
        );

    \pid_side.error_d_reg_prev_esr_RNI2VN9_0_12_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__51537\,
            in1 => \_gnd_net_\,
            in2 => \N__54657\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \pid_side.N_1590_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNIVTFJ2_12_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__54710\,
            in1 => \N__51123\,
            in2 => \N__51105\,
            in3 => \N__51549\,
            lcout => \pid_side.error_d_reg_esr_RNIVTFJ2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIVKIO_12_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__51536\,
            in1 => \_gnd_net_\,
            in2 => \N__54656\,
            in3 => \N__54709\,
            lcout => \pid_side.un1_pid_prereg_107_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__51482\,
            in1 => \N__51507\,
            in2 => \_gnd_net_\,
            in3 => \N__54868\,
            lcout => \pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNI2VN9_12_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54649\,
            in2 => \_gnd_net_\,
            in3 => \N__51535\,
            lcout => \pid_side.error_d_reg_prev_esr_RNI2VN9Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_11_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59207\,
            ce => \N__57958\,
            sr => \N__57614\
        );

    \pid_side.error_p_reg_esr_11_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51495\,
            lcout => \pid_side.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59222\,
            ce => \N__56607\,
            sr => \N__58188\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__51468\,
            in1 => \N__51405\,
            in2 => \_gnd_net_\,
            in3 => \N__51273\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54681\,
            in1 => \N__51843\,
            in2 => \_gnd_net_\,
            in3 => \N__55043\,
            lcout => \pid_side.un1_pid_prereg_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_19_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__55044\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59239\,
            ce => \N__57962\,
            sr => \N__57629\
        );

    \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54680\,
            in1 => \N__51842\,
            in2 => \_gnd_net_\,
            in3 => \N__55042\,
            lcout => \pid_side.un1_pid_prereg_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH2data_esr_3_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55372\,
            lcout => side_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59255\,
            ce => \N__51809\,
            sr => \N__57634\
        );

    \pid_side.error_cry_0_c_inv_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51756\,
            in2 => \_gnd_net_\,
            in3 => \N__51772\,
            lcout => \pid_side.error_axb_0\,
            ltout => OPEN,
            carryin => \bfn_21_17_0_\,
            carryout => \pid_side.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_0_c_RNI43F5_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51750\,
            in2 => \_gnd_net_\,
            in3 => \N__51717\,
            lcout => \pid_side.error_1\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_0\,
            carryout => \pid_side.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_1_c_RNI66G5_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51714\,
            in2 => \_gnd_net_\,
            in3 => \N__51681\,
            lcout => \pid_side.error_2\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_1\,
            carryout => \pid_side.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_2_c_RNI89H5_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51678\,
            in2 => \_gnd_net_\,
            in3 => \N__51648\,
            lcout => \pid_side.error_3\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_2\,
            carryout => \pid_side.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_3_c_RNI1SDJ_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51645\,
            in2 => \N__51639\,
            in3 => \N__51603\,
            lcout => \pid_side.error_4\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_3\,
            carryout => \pid_side.error_cry_0_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_0_0_c_RNIF3ET_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51600\,
            in2 => \N__51591\,
            in3 => \N__51558\,
            lcout => \pid_side.error_5\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_0_0\,
            carryout => \pid_side.error_cry_1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_1_0_c_RNII9K11_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52191\,
            in2 => \N__52185\,
            in3 => \N__52149\,
            lcout => \pid_side.error_6\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_1_0\,
            carryout => \pid_side.error_cry_2_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_2_0_c_RNILFQL_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52146\,
            in2 => \N__52140\,
            in3 => \N__52110\,
            lcout => \pid_side.error_7\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_2_0\,
            carryout => \pid_side.error_cry_3_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_3_0_c_RNIOL0Q_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52107\,
            in2 => \N__52101\,
            in3 => \N__52065\,
            lcout => \pid_side.error_8\,
            ltout => OPEN,
            carryin => \bfn_21_18_0_\,
            carryout => \pid_side.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_4_c_RNIC8FJ_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52062\,
            in2 => \N__52044\,
            in3 => \N__52011\,
            lcout => \pid_side.error_9\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_4\,
            carryout => \pid_side.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_5_c_RNIM4IS_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52008\,
            in2 => \N__51996\,
            in3 => \N__51954\,
            lcout => \pid_side.error_10\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_5\,
            carryout => \pid_side.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_6_c_RNIQBMT_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51951\,
            in2 => \_gnd_net_\,
            in3 => \N__51918\,
            lcout => \pid_side.error_11\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_6\,
            carryout => \pid_side.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_7_c_RNIPRDP1_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51915\,
            in2 => \N__52506\,
            in3 => \N__51882\,
            lcout => \pid_side.error_12\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_7\,
            carryout => \pid_side.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_8_c_RNIUUKS_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51879\,
            in2 => \N__52410\,
            in3 => \N__51846\,
            lcout => \pid_side.error_13\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_8\,
            carryout => \pid_side.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_9_c_RNI13MS_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53141\,
            in2 => \N__52779\,
            in3 => \N__52746\,
            lcout => \pid_side.error_14\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_9\,
            carryout => \pid_side.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_10_c_RNIBCT11_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__53142\,
            in1 => \N__52317\,
            in2 => \_gnd_net_\,
            in3 => \N__52743\,
            lcout => \pid_side.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52713\,
            lcout => \drone_H_disp_side_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59294\,
            ce => \N__53129\,
            sr => \N__57648\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__52586\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \drone_H_disp_side_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59294\,
            ce => \N__53129\,
            sr => \N__57648\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52488\,
            lcout => \drone_H_disp_side_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59294\,
            ce => \N__53129\,
            sr => \N__57648\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52384\,
            lcout => \drone_H_disp_side_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59294\,
            ce => \N__53129\,
            sr => \N__57648\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52311\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59294\,
            ce => \N__53129\,
            sr => \N__57648\
        );

    \pid_front.error_d_reg_esr_6_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52230\,
            lcout => \pid_front.error_d_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59319\,
            ce => \N__58502\,
            sr => \N__58181\
        );

    \pid_side.error_d_reg_esr_RNI76TK1_5_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000101000"
        )
    port map (
            in0 => \N__54752\,
            in1 => \N__53815\,
            in2 => \N__53795\,
            in3 => \N__52845\,
            lcout => \pid_side.error_d_reg_esr_RNI76TK1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNILKEQ_5_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__53814\,
            in1 => \N__53788\,
            in2 => \_gnd_net_\,
            in3 => \N__54751\,
            lcout => OPEN,
            ltout => \pid_side.un1_pid_prereg_40_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNI86Q93_5_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__52812\,
            in1 => \N__53601\,
            in2 => \N__52860\,
            in3 => \N__52844\,
            lcout => \pid_side.error_d_reg_esr_RNI86Q93Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54278\,
            in1 => \N__52820\,
            in2 => \_gnd_net_\,
            in3 => \N__53458\,
            lcout => \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__53459\,
            in1 => \_gnd_net_\,
            in2 => \N__52824\,
            in3 => \N__54279\,
            lcout => \pid_side.un1_pid_prereg_17\,
            ltout => \pid_side.un1_pid_prereg_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNI10TK1_3_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52836\,
            in3 => \N__53600\,
            lcout => \pid_side.error_p_reg_esr_RNI10TK1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_4_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__53460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59168\,
            ce => \N__57954\,
            sr => \N__57592\
        );

    \pid_side.error_p_reg_esr_RNISPP93_2_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__53672\,
            in1 => \N__53599\,
            in2 => \N__53628\,
            in3 => \N__52811\,
            lcout => \pid_side.error_p_reg_esr_RNISPP93Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_5_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__52791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59180\,
            ce => \N__56592\,
            sr => \N__58196\
        );

    \pid_side.error_p_reg_esr_0_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53031\,
            lcout => \pid_side.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59180\,
            ce => \N__56592\,
            sr => \N__58196\
        );

    \pid_side.state_RNIK1B71_0_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53010\,
            in2 => \_gnd_net_\,
            in3 => \N__58321\,
            lcout => \pid_side.N_599_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIE47J_9_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54348\,
            in2 => \_gnd_net_\,
            in3 => \N__54139\,
            lcout => \pid_side.error_p_reg_esr_RNIE47JZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_15_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54812\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59208\,
            ce => \N__57959\,
            sr => \N__57615\
        );

    \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__53573\,
            in1 => \N__54432\,
            in2 => \_gnd_net_\,
            in3 => \N__55168\,
            lcout => \pid_side.un1_pid_prereg_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54218\,
            in1 => \N__52904\,
            in2 => \_gnd_net_\,
            in3 => \N__54982\,
            lcout => \pid_side.un1_pid_prereg_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_18_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54984\,
            lcout => \pid_side.error_d_reg_prevZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59223\,
            ce => \N__57960\,
            sr => \N__57622\
        );

    \pid_side.error_d_reg_prev_esr_RNIOHC23_16_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__52938\,
            in1 => \N__52889\,
            in2 => \N__54123\,
            in3 => \N__54094\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIOHC23Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_22_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__54983\,
            in1 => \_gnd_net_\,
            in2 => \N__52908\,
            in3 => \N__54219\,
            lcout => \pid_side.un1_pid_prereg_47\,
            ltout => \pid_side.un1_pid_prereg_47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIVB6H1_17_LC_22_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__54095\,
            in1 => \_gnd_net_\,
            in2 => \N__53556\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prev_esr_RNIVB6H1Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_10_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55080\,
            lcout => \pid_side.error_d_reg_prevZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59240\,
            ce => \N__57963\,
            sr => \N__57630\
        );

    \pid_side.error_d_reg_esr_0_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53520\,
            lcout => \pid_side.error_d_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59256\,
            ce => \N__56593\,
            sr => \N__58189\
        );

    \pid_side.error_d_reg_esr_4_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53472\,
            lcout => \pid_side.error_d_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59256\,
            ce => \N__56593\,
            sr => \N__58189\
        );

    \pid_side.error_d_reg_esr_1_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53445\,
            lcout => \pid_side.error_d_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59256\,
            ce => \N__56593\,
            sr => \N__58189\
        );

    \Commands_frame_decoder.source_xy_kd_4_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53396\,
            in2 => \_gnd_net_\,
            in3 => \N__58322\,
            lcout => xy_kd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59285\,
            ce => \N__55205\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53229\,
            lcout => \drone_H_disp_side_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59295\,
            ce => \N__53133\,
            sr => \N__57649\
        );

    \pid_front.error_d_reg_esr_5_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__53094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59322\,
            ce => \N__58495\,
            sr => \N__58182\
        );

    \pid_side.error_p_reg_esr_RNI5PH23_1_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__53058\,
            in1 => \N__53623\,
            in2 => \N__53673\,
            in3 => \N__53644\,
            lcout => \pid_side.error_p_reg_esr_RNI5PH23Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54240\,
            in1 => \N__53610\,
            in2 => \_gnd_net_\,
            in3 => \N__55133\,
            lcout => \pid_side.un1_pid_prereg_2\,
            ltout => \pid_side.un1_pid_prereg_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIRPSK1_2_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__53658\,
            in3 => \N__53624\,
            lcout => \pid_side.error_p_reg_esr_RNIRPSK1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54197\,
            in1 => \N__53582\,
            in2 => \_gnd_net_\,
            in3 => \N__54535\,
            lcout => \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNICBEQ_2_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__54536\,
            in1 => \_gnd_net_\,
            in2 => \N__53586\,
            in3 => \N__54198\,
            lcout => \pid_side.un1_pid_prereg_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_3_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__55134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59181\,
            ce => \N__57955\,
            sr => \N__57600\
        );

    \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_23_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54239\,
            in1 => \N__53609\,
            in2 => \_gnd_net_\,
            in3 => \N__55132\,
            lcout => \pid_side.un1_pid_prereg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_2_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54537\,
            lcout => \pid_side.error_d_reg_prevZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59196\,
            ce => \N__57957\,
            sr => \N__57608\
        );

    \pid_side.error_d_reg_prev_esr_14_LC_23_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55170\,
            lcout => \pid_side.error_d_reg_prevZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59196\,
            ce => \N__57957\,
            sr => \N__57608\
        );

    \pid_side.error_p_reg_esr_RNI8U6J_6_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54930\,
            in2 => \_gnd_net_\,
            in3 => \N__54912\,
            lcout => OPEN,
            ltout => \pid_side.N_1566_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNIUJLD1_6_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__53819\,
            in1 => \N__53796\,
            in2 => \N__53763\,
            in3 => \N__55014\,
            lcout => \pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIE47J_0_9_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54347\,
            in2 => \_gnd_net_\,
            in3 => \N__54141\,
            lcout => OPEN,
            ltout => \pid_side.N_1578_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNID3MD1_9_LC_23_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__54057\,
            in1 => \N__54489\,
            in2 => \N__53760\,
            in3 => \N__53691\,
            lcout => \pid_side.error_d_reg_esr_RNID3MD1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNI11FQ_9_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54052\,
            in1 => \N__54346\,
            in2 => \_gnd_net_\,
            in3 => \N__54140\,
            lcout => \pid_side.un1_pid_prereg_80_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_8_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54777\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59224\,
            ce => \N__57961\,
            sr => \N__57623\
        );

    \pid_side.error_p_reg_esr_RNIC27J_8_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__53689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54493\,
            lcout => OPEN,
            ltout => \pid_side.N_1574_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNI8ULD1_8_LC_23_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__54776\,
            in1 => \N__54570\,
            in2 => \N__53730\,
            in3 => \N__54960\,
            lcout => \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8\,
            ltout => \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIL1CR2_8_LC_23_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110011001"
        )
    port map (
            in0 => \N__53690\,
            in1 => \N__53712\,
            in2 => \N__53706\,
            in3 => \N__54494\,
            lcout => \pid_side.error_p_reg_esr_RNIL1CR2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNIUTEQ_8_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__54775\,
            in1 => \_gnd_net_\,
            in2 => \N__54495\,
            in3 => \N__53688\,
            lcout => \pid_side.un1_pid_prereg_70_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_9_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59224\,
            ce => \N__57961\,
            sr => \N__57623\
        );

    \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__54836\,
            in1 => \_gnd_net_\,
            in2 => \N__54081\,
            in3 => \N__54153\,
            lcout => \pid_side.un1_pid_prereg_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__54152\,
            in1 => \N__54077\,
            in2 => \_gnd_net_\,
            in3 => \N__54835\,
            lcout => \pid_side.un1_pid_prereg_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_17_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54837\,
            lcout => \pid_side.error_d_reg_prevZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59257\,
            ce => \N__57965\,
            sr => \N__57635\
        );

    \pid_side.error_d_reg_esr_9_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54069\,
            lcout => \pid_side.error_d_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59272\,
            ce => \N__56598\,
            sr => \N__58190\
        );

    \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__57980\,
            in1 => \N__54458\,
            in2 => \_gnd_net_\,
            in3 => \N__57997\,
            lcout => \pid_side.un1_pid_prereg_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__54462\,
            in1 => \N__57981\,
            in2 => \_gnd_net_\,
            in3 => \N__58004\,
            lcout => \pid_side.un1_pid_prereg_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_d_reg_esr_8_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53928\,
            lcout => \pid_front.error_d_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59327\,
            ce => \N__58523\,
            sr => \N__58183\
        );

    \pid_front.error_d_reg_esr_12_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53865\,
            lcout => \pid_front.error_d_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59327\,
            ce => \N__58523\,
            sr => \N__58183\
        );

    \pid_front.error_d_reg_esr_10_LC_23_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54327\,
            lcout => \pid_front.error_d_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59327\,
            ce => \N__58523\,
            sr => \N__58183\
        );

    \pid_side.error_p_reg_esr_4_LC_24_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54288\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59197\,
            ce => \N__56603\,
            sr => \N__58204\
        );

    \pid_side.error_p_reg_esr_1_LC_24_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54267\,
            lcout => \pid_side.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59197\,
            ce => \N__56603\,
            sr => \N__58204\
        );

    \pid_side.error_p_reg_esr_3_LC_24_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54246\,
            lcout => \pid_side.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59197\,
            ce => \N__56603\,
            sr => \N__58204\
        );

    \pid_side.error_p_reg_esr_18_LC_24_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54231\,
            lcout => \pid_side.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59197\,
            ce => \N__56603\,
            sr => \N__58204\
        );

    \pid_side.error_p_reg_esr_2_LC_24_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54204\,
            lcout => \pid_side.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59197\,
            ce => \N__56603\,
            sr => \N__58204\
        );

    \pid_side.error_p_reg_esr_16_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54189\,
            lcout => \pid_side.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59209\,
            ce => \N__56608\,
            sr => \N__58202\
        );

    \pid_side.error_p_reg_esr_17_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54162\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59209\,
            ce => \N__56608\,
            sr => \N__58202\
        );

    \pid_side.error_d_reg_esr_2_LC_24_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54549\,
            lcout => \pid_side.error_d_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59209\,
            ce => \N__56608\,
            sr => \N__58202\
        );

    \pid_side.error_p_reg_esr_13_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54522\,
            lcout => \pid_side.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59209\,
            ce => \N__56608\,
            sr => \N__58202\
        );

    \pid_side.error_p_reg_esr_8_LC_24_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54501\,
            lcout => \pid_side.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59209\,
            ce => \N__56608\,
            sr => \N__58202\
        );

    \pid_side.error_p_reg_esr_20_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54471\,
            lcout => \pid_side.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59209\,
            ce => \N__56608\,
            sr => \N__58202\
        );

    \pid_side.error_p_reg_esr_14_LC_24_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54441\,
            lcout => \pid_side.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59209\,
            ce => \N__56608\,
            sr => \N__58202\
        );

    \pid_side.error_p_reg_esr_10_LC_24_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54411\,
            lcout => \pid_side.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59225\,
            ce => \N__56564\,
            sr => \N__58199\
        );

    \pid_side.error_p_reg_esr_15_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54384\,
            lcout => \pid_side.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59225\,
            ce => \N__56564\,
            sr => \N__58199\
        );

    \pid_side.error_p_reg_esr_6_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54360\,
            lcout => \pid_side.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59225\,
            ce => \N__56564\,
            sr => \N__58199\
        );

    \pid_side.error_p_reg_esr_9_LC_24_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54354\,
            lcout => \pid_side.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59225\,
            ce => \N__56564\,
            sr => \N__58199\
        );

    \pid_side.error_p_reg_esr_7_LC_24_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54693\,
            lcout => \pid_side.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59225\,
            ce => \N__56564\,
            sr => \N__58199\
        );

    \pid_side.error_p_reg_esr_19_LC_24_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54687\,
            lcout => \pid_side.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59225\,
            ce => \N__56564\,
            sr => \N__58199\
        );

    \pid_side.error_p_reg_esr_12_LC_24_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54663\,
            lcout => \pid_side.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59225\,
            ce => \N__56564\,
            sr => \N__58199\
        );

    \pid_side.error_d_reg_prev_esr_7_LC_24_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56649\,
            lcout => \pid_side.error_d_reg_prevZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59241\,
            ce => \N__57964\,
            sr => \N__57631\
        );

    \pid_side.error_d_reg_esr_RNIRQEQ_7_LC_24_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56647\,
            in1 => \N__54567\,
            in2 => \_gnd_net_\,
            in3 => \N__54957\,
            lcout => OPEN,
            ltout => \pid_side.un1_pid_prereg_60_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNI1DBR2_6_LC_24_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110100101"
        )
    port map (
            in0 => \N__54910\,
            in1 => \N__54629\,
            in2 => \N__54615\,
            in3 => \N__54928\,
            lcout => \pid_side.error_p_reg_esr_RNI1DBR2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIA07J_7_LC_24_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54568\,
            in2 => \_gnd_net_\,
            in3 => \N__54958\,
            lcout => OPEN,
            ltout => \pid_side.N_1570_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_RNI3PLD1_7_LC_24_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101001101"
        )
    port map (
            in0 => \N__54911\,
            in1 => \N__56648\,
            in2 => \N__54594\,
            in3 => \N__54929\,
            lcout => \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7\,
            ltout => \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_esr_RNIBNBR2_7_LC_24_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001010101"
        )
    port map (
            in0 => \N__54576\,
            in1 => \N__54569\,
            in2 => \N__54552\,
            in3 => \N__54959\,
            lcout => \pid_side.error_p_reg_esr_RNIBNBR2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_6_LC_24_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__55010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_reg_prevZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59241\,
            ce => \N__57964\,
            sr => \N__57631\
        );

    \pid_side.error_d_reg_esr_RNIONEQ_6_LC_24_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54927\,
            in1 => \N__54909\,
            in2 => \_gnd_net_\,
            in3 => \N__55009\,
            lcout => \pid_side.un1_pid_prereg_50_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_esr_11_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54882\,
            lcout => \pid_side.error_d_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59258\,
            ce => \N__56597\,
            sr => \N__58195\
        );

    \pid_side.error_d_reg_esr_17_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_d_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_15_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54822\,
            lcout => \pid_side.error_d_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_8_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54786\,
            lcout => \pid_side.error_d_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_5_LC_24_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54762\,
            lcout => \pid_side.error_d_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_12_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54720\,
            lcout => \pid_side.error_d_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_14_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55179\,
            lcout => \pid_side.error_d_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_3_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55140\,
            lcout => \pid_side.error_d_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_13_LC_24_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55116\,
            lcout => \pid_side.error_d_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59273\,
            ce => \N__56610\,
            sr => \N__58194\
        );

    \pid_side.error_d_reg_esr_10_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55086\,
            lcout => \pid_side.error_d_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59286\,
            ce => \N__56599\,
            sr => \N__58192\
        );

    \pid_side.error_d_reg_esr_19_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55053\,
            lcout => \pid_side.error_d_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59286\,
            ce => \N__56599\,
            sr => \N__58192\
        );

    \pid_side.error_d_reg_esr_20_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55029\,
            lcout => \pid_side.error_d_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59286\,
            ce => \N__56599\,
            sr => \N__58192\
        );

    \pid_side.error_d_reg_esr_6_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55020\,
            lcout => \pid_side.error_d_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59286\,
            ce => \N__56599\,
            sr => \N__58192\
        );

    \pid_side.error_d_reg_esr_18_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54993\,
            lcout => \pid_side.error_d_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59286\,
            ce => \N__56599\,
            sr => \N__58192\
        );

    \pid_side.error_d_reg_esr_7_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54966\,
            lcout => \pid_side.error_d_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59286\,
            ce => \N__56599\,
            sr => \N__58192\
        );

    \pid_side.error_d_reg_esr_16_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56634\,
            lcout => \pid_side.error_d_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59296\,
            ce => \N__56609\,
            sr => \N__58191\
        );

    \Commands_frame_decoder.source_xy_kd_0_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56508\,
            in2 => \_gnd_net_\,
            in3 => \N__58323\,
            lcout => xy_kd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59304\,
            ce => \N__55212\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kd_1_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56313\,
            lcout => xy_kd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59304\,
            ce => \N__55212\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kd_2_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56140\,
            in2 => \_gnd_net_\,
            in3 => \N__58325\,
            lcout => xy_kd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59304\,
            ce => \N__55212\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kd_5_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55931\,
            in2 => \_gnd_net_\,
            in3 => \N__58327\,
            lcout => xy_kd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59304\,
            ce => \N__55212\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kd_6_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58328\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55754\,
            lcout => xy_kd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59304\,
            ce => \N__55212\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kd_7_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55582\,
            in2 => \_gnd_net_\,
            in3 => \N__58329\,
            lcout => xy_kd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59304\,
            ce => \N__55212\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kd_3_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55362\,
            lcout => xy_kd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59304\,
            ce => \N__55212\,
            sr => \_gnd_net_\
        );

    \pid_side.error_d_reg_prev_esr_20_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58005\,
            lcout => \pid_side.error_d_reg_prevZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59316\,
            ce => \N__57966\,
            sr => \N__57650\
        );

    \pid_front.error_d_reg_esr_0_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56949\,
            lcout => \pid_front.error_d_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59323\,
            ce => \N__58536\,
            sr => \N__58187\
        );

    \pid_front.error_d_reg_esr_1_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56901\,
            lcout => \pid_front.error_d_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59328\,
            ce => \N__58534\,
            sr => \N__58186\
        );

    \pid_front.error_d_reg_esr_13_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56859\,
            lcout => \pid_front.error_d_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59328\,
            ce => \N__58534\,
            sr => \N__58186\
        );

    \pid_front.error_d_reg_esr_11_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56832\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59328\,
            ce => \N__58534\,
            sr => \N__58186\
        );

    \pid_front.error_d_reg_esr_9_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56784\,
            lcout => \pid_front.error_d_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59328\,
            ce => \N__58534\,
            sr => \N__58186\
        );

    \pid_front.error_d_reg_esr_16_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56736\,
            lcout => \pid_front.error_d_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59332\,
            ce => \N__58524\,
            sr => \N__58185\
        );

    \pid_front.error_d_reg_esr_17_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56682\,
            lcout => \pid_front.error_d_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59332\,
            ce => \N__58524\,
            sr => \N__58185\
        );

    \pid_front.error_d_reg_esr_18_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__59583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59332\,
            ce => \N__58524\,
            sr => \N__58185\
        );

    \pid_front.error_d_reg_esr_19_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59538\,
            lcout => \pid_front.error_d_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59332\,
            ce => \N__58524\,
            sr => \N__58185\
        );

    \pid_front.error_d_reg_esr_20_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__59511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_d_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59332\,
            ce => \N__58524\,
            sr => \N__58185\
        );

    \pid_front.error_d_reg_esr_14_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59475\,
            lcout => \pid_front.error_d_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59332\,
            ce => \N__58524\,
            sr => \N__58185\
        );

    \pid_front.error_d_reg_esr_4_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59433\,
            lcout => \pid_front.error_d_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59332\,
            ce => \N__58524\,
            sr => \N__58185\
        );

    \pid_front.error_d_reg_esr_7_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59403\,
            lcout => \pid_front.error_d_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59335\,
            ce => \N__58535\,
            sr => \N__58184\
        );

    \pid_front.error_d_reg_esr_15_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59367\,
            lcout => \pid_front.error_d_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__59335\,
            ce => \N__58535\,
            sr => \N__58184\
        );
end \INTERFACE\;
