// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 10 2019 19:42:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2Drone" view "INTERFACE"

module Pc2Drone (
    data,
    uart_input,
    data_rdy,
    uart_input_debug,
    clk_system);

    output [7:0] data;
    input uart_input;
    output data_rdy;
    output uart_input_debug;
    input clk_system;

    wire N__3233;
    wire N__3232;
    wire N__3231;
    wire N__3222;
    wire N__3221;
    wire N__3220;
    wire N__3213;
    wire N__3212;
    wire N__3211;
    wire N__3204;
    wire N__3203;
    wire N__3202;
    wire N__3195;
    wire N__3194;
    wire N__3193;
    wire N__3186;
    wire N__3185;
    wire N__3184;
    wire N__3177;
    wire N__3176;
    wire N__3175;
    wire N__3168;
    wire N__3167;
    wire N__3166;
    wire N__3159;
    wire N__3158;
    wire N__3157;
    wire N__3150;
    wire N__3149;
    wire N__3148;
    wire N__3141;
    wire N__3140;
    wire N__3139;
    wire N__3132;
    wire N__3131;
    wire N__3130;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2922;
    wire N__2917;
    wire N__2914;
    wire N__2909;
    wire N__2908;
    wire N__2907;
    wire N__2906;
    wire N__2903;
    wire N__2902;
    wire N__2901;
    wire N__2898;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2875;
    wire N__2870;
    wire N__2867;
    wire N__2866;
    wire N__2859;
    wire N__2858;
    wire N__2857;
    wire N__2856;
    wire N__2851;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2812;
    wire N__2807;
    wire N__2806;
    wire N__2803;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2761;
    wire N__2760;
    wire N__2759;
    wire N__2758;
    wire N__2757;
    wire N__2756;
    wire N__2755;
    wire N__2754;
    wire N__2753;
    wire N__2752;
    wire N__2751;
    wire N__2750;
    wire N__2749;
    wire N__2748;
    wire N__2747;
    wire N__2746;
    wire N__2745;
    wire N__2744;
    wire N__2743;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2676;
    wire N__2675;
    wire N__2670;
    wire N__2667;
    wire N__2664;
    wire N__2663;
    wire N__2662;
    wire N__2661;
    wire N__2660;
    wire N__2659;
    wire N__2654;
    wire N__2651;
    wire N__2650;
    wire N__2649;
    wire N__2648;
    wire N__2647;
    wire N__2646;
    wire N__2645;
    wire N__2640;
    wire N__2635;
    wire N__2632;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2616;
    wire N__2611;
    wire N__2606;
    wire N__2591;
    wire N__2588;
    wire N__2587;
    wire N__2586;
    wire N__2585;
    wire N__2582;
    wire N__2581;
    wire N__2580;
    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2574;
    wire N__2573;
    wire N__2572;
    wire N__2571;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2556;
    wire N__2553;
    wire N__2546;
    wire N__2541;
    wire N__2536;
    wire N__2519;
    wire N__2518;
    wire N__2517;
    wire N__2514;
    wire N__2511;
    wire N__2510;
    wire N__2509;
    wire N__2508;
    wire N__2503;
    wire N__2500;
    wire N__2497;
    wire N__2494;
    wire N__2491;
    wire N__2490;
    wire N__2489;
    wire N__2488;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2472;
    wire N__2469;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2455;
    wire N__2452;
    wire N__2449;
    wire N__2438;
    wire N__2437;
    wire N__2436;
    wire N__2435;
    wire N__2434;
    wire N__2433;
    wire N__2430;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2418;
    wire N__2415;
    wire N__2410;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2248;
    wire N__2245;
    wire N__2242;
    wire N__2237;
    wire N__2236;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2213;
    wire N__2210;
    wire N__2209;
    wire N__2206;
    wire N__2205;
    wire N__2204;
    wire N__2203;
    wire N__2202;
    wire N__2201;
    wire N__2200;
    wire N__2199;
    wire N__2196;
    wire N__2193;
    wire N__2186;
    wire N__2179;
    wire N__2178;
    wire N__2177;
    wire N__2176;
    wire N__2175;
    wire N__2174;
    wire N__2171;
    wire N__2168;
    wire N__2161;
    wire N__2158;
    wire N__2155;
    wire N__2148;
    wire N__2135;
    wire N__2134;
    wire N__2133;
    wire N__2132;
    wire N__2131;
    wire N__2130;
    wire N__2127;
    wire N__2124;
    wire N__2117;
    wire N__2116;
    wire N__2115;
    wire N__2114;
    wire N__2111;
    wire N__2104;
    wire N__2099;
    wire N__2098;
    wire N__2097;
    wire N__2096;
    wire N__2093;
    wire N__2086;
    wire N__2081;
    wire N__2078;
    wire N__2069;
    wire N__2068;
    wire N__2065;
    wire N__2064;
    wire N__2057;
    wire N__2054;
    wire N__2051;
    wire N__2050;
    wire N__2049;
    wire N__2048;
    wire N__2039;
    wire N__2036;
    wire N__2033;
    wire N__2032;
    wire N__2031;
    wire N__2028;
    wire N__2027;
    wire N__2024;
    wire N__2023;
    wire N__2022;
    wire N__2019;
    wire N__2018;
    wire N__2017;
    wire N__2014;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__1996;
    wire N__1985;
    wire N__1982;
    wire N__1981;
    wire N__1980;
    wire N__1979;
    wire N__1978;
    wire N__1977;
    wire N__1976;
    wire N__1975;
    wire N__1974;
    wire N__1971;
    wire N__1966;
    wire N__1963;
    wire N__1960;
    wire N__1951;
    wire N__1940;
    wire N__1939;
    wire N__1938;
    wire N__1937;
    wire N__1936;
    wire N__1935;
    wire N__1934;
    wire N__1933;
    wire N__1932;
    wire N__1931;
    wire N__1928;
    wire N__1927;
    wire N__1924;
    wire N__1923;
    wire N__1920;
    wire N__1917;
    wire N__1914;
    wire N__1911;
    wire N__1904;
    wire N__1901;
    wire N__1900;
    wire N__1897;
    wire N__1894;
    wire N__1891;
    wire N__1884;
    wire N__1881;
    wire N__1876;
    wire N__1871;
    wire N__1856;
    wire N__1853;
    wire N__1852;
    wire N__1847;
    wire N__1846;
    wire N__1845;
    wire N__1844;
    wire N__1843;
    wire N__1842;
    wire N__1839;
    wire N__1838;
    wire N__1837;
    wire N__1836;
    wire N__1833;
    wire N__1832;
    wire N__1831;
    wire N__1830;
    wire N__1829;
    wire N__1828;
    wire N__1819;
    wire N__1816;
    wire N__1809;
    wire N__1806;
    wire N__1799;
    wire N__1794;
    wire N__1781;
    wire N__1780;
    wire N__1779;
    wire N__1776;
    wire N__1773;
    wire N__1770;
    wire N__1767;
    wire N__1762;
    wire N__1759;
    wire N__1756;
    wire N__1751;
    wire N__1750;
    wire N__1749;
    wire N__1748;
    wire N__1747;
    wire N__1744;
    wire N__1739;
    wire N__1734;
    wire N__1727;
    wire N__1726;
    wire N__1725;
    wire N__1724;
    wire N__1723;
    wire N__1718;
    wire N__1713;
    wire N__1710;
    wire N__1703;
    wire N__1702;
    wire N__1699;
    wire N__1696;
    wire N__1693;
    wire N__1692;
    wire N__1689;
    wire N__1686;
    wire N__1683;
    wire N__1680;
    wire N__1675;
    wire N__1670;
    wire N__1667;
    wire N__1666;
    wire N__1665;
    wire N__1664;
    wire N__1661;
    wire N__1660;
    wire N__1659;
    wire N__1658;
    wire N__1657;
    wire N__1654;
    wire N__1651;
    wire N__1648;
    wire N__1645;
    wire N__1638;
    wire N__1635;
    wire N__1632;
    wire N__1629;
    wire N__1616;
    wire N__1615;
    wire N__1612;
    wire N__1611;
    wire N__1610;
    wire N__1609;
    wire N__1608;
    wire N__1607;
    wire N__1606;
    wire N__1605;
    wire N__1604;
    wire N__1599;
    wire N__1592;
    wire N__1591;
    wire N__1590;
    wire N__1589;
    wire N__1588;
    wire N__1585;
    wire N__1582;
    wire N__1575;
    wire N__1570;
    wire N__1565;
    wire N__1560;
    wire N__1547;
    wire N__1544;
    wire N__1541;
    wire N__1538;
    wire N__1535;
    wire N__1532;
    wire N__1529;
    wire N__1526;
    wire N__1523;
    wire N__1520;
    wire N__1517;
    wire N__1516;
    wire N__1515;
    wire N__1512;
    wire N__1509;
    wire N__1508;
    wire N__1507;
    wire N__1506;
    wire N__1503;
    wire N__1500;
    wire N__1497;
    wire N__1494;
    wire N__1489;
    wire N__1478;
    wire N__1477;
    wire N__1476;
    wire N__1473;
    wire N__1470;
    wire N__1467;
    wire N__1464;
    wire N__1457;
    wire N__1454;
    wire N__1451;
    wire N__1448;
    wire N__1445;
    wire N__1442;
    wire N__1441;
    wire N__1438;
    wire N__1435;
    wire N__1430;
    wire N__1427;
    wire N__1424;
    wire N__1421;
    wire N__1418;
    wire N__1415;
    wire N__1412;
    wire N__1409;
    wire N__1406;
    wire N__1403;
    wire N__1402;
    wire N__1399;
    wire N__1396;
    wire N__1393;
    wire N__1388;
    wire N__1385;
    wire N__1382;
    wire N__1379;
    wire N__1376;
    wire N__1373;
    wire N__1372;
    wire N__1371;
    wire N__1370;
    wire N__1367;
    wire N__1366;
    wire N__1365;
    wire N__1364;
    wire N__1361;
    wire N__1356;
    wire N__1355;
    wire N__1350;
    wire N__1345;
    wire N__1340;
    wire N__1337;
    wire N__1328;
    wire N__1325;
    wire N__1322;
    wire N__1319;
    wire N__1316;
    wire N__1313;
    wire N__1310;
    wire N__1307;
    wire N__1306;
    wire N__1303;
    wire N__1300;
    wire N__1295;
    wire N__1292;
    wire N__1291;
    wire N__1286;
    wire N__1283;
    wire N__1280;
    wire N__1277;
    wire N__1274;
    wire N__1271;
    wire N__1268;
    wire N__1265;
    wire N__1262;
    wire N__1261;
    wire N__1260;
    wire N__1257;
    wire N__1254;
    wire N__1253;
    wire N__1244;
    wire N__1241;
    wire N__1240;
    wire N__1237;
    wire N__1236;
    wire N__1229;
    wire N__1226;
    wire N__1223;
    wire N__1220;
    wire N__1217;
    wire N__1214;
    wire N__1211;
    wire N__1208;
    wire N__1205;
    wire GNDG0;
    wire VCCG0;
    wire \uart.CO0_0_cascade_ ;
    wire \uart.bit_Count_RNO_1Z0Z_2_cascade_ ;
    wire \uart.CO1_1_cascade_ ;
    wire \uart.bit_Count_RNO_2Z0Z_2 ;
    wire \uart.bit_Count_RNO_1Z0Z_1 ;
    wire \uart.state_RNO_1Z0Z_2_cascade_ ;
    wire \uart.state_RNO_2Z0Z_2 ;
    wire \uart.N_170_cascade_ ;
    wire \uart.stateZ0Z_2 ;
    wire \uart.stateZ0Z_1 ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_7_cascade_ ;
    wire \uart.N_44_0 ;
    wire \uart.N_147_0_cascade_ ;
    wire \uart.timer_Count_RNITC202Z0Z_6 ;
    wire \uart.timer_Count_RNIGLM11Z0Z_6_cascade_ ;
    wire \uart.un1_state_7_0_0 ;
    wire \uart.un1_state_7_0_0_cascade_ ;
    wire \uart.N_177 ;
    wire \uart.un1_state_5 ;
    wire \uart.state_RNO_0Z0Z_3 ;
    wire \uart.state_RNO_1Z0Z_3 ;
    wire \uart.N_147_0 ;
    wire \uart.N_159 ;
    wire \uart.timer_Count_6_rep1_RNIRC5SZ0Z1_cascade_ ;
    wire \uart.un1_state_2_0_a3_0_cascade_ ;
    wire \uart.timer_CountZ0Z_6 ;
    wire \uart.timer_Count_fastZ0Z_6 ;
    wire \uart.un1_state_4_0_a2_iso_cascade_ ;
    wire \uart.N_38_0 ;
    wire \uart.N_165_1 ;
    wire \uart.timer_Count_RNIICSG1Z0Z_6 ;
    wire \uart.N_175_cascade_ ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_1 ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_ ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_ ;
    wire \uart.timer_Count_6_repZ0Z1 ;
    wire \uart.un4_timer_Count_1_c2 ;
    wire \uart.timer_Count_RNIMLMA1Z0Z_1_cascade_ ;
    wire \uart.un4_timer_Count_1_c5 ;
    wire \uart.un4_timer_Count_1_c5_cascade_ ;
    wire \uart.timer_CountZ0Z_3 ;
    wire \uart.timer_CountZ0Z_2 ;
    wire \uart.stateZ0Z_3 ;
    wire \uart.timer_Count_RNIHJ661Z0Z_3_cascade_ ;
    wire \uart.timer_CountZ0Z_5 ;
    wire \uart.state_0_sqmuxa_1_d ;
    wire \uart.timer_CountZ0Z_0 ;
    wire \uart.timer_CountZ0Z_1 ;
    wire \uart.un1_timer_Count_0_sqmuxa_0 ;
    wire \uart.timer_CountZ0Z_4 ;
    wire \uart.timer_CountZ0Z_7 ;
    wire \uart.N_28_mux_i_i_0 ;
    wire \uart.N_22_mux ;
    wire data_rdy_c;
    wire \uart.data_Aux_esr_RNO_0Z0Z_0 ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_4 ;
    wire \uart.N_39_0 ;
    wire \uart.N_40_0 ;
    wire \uart.timer_Count_6_rep1_RNI1B4SZ0 ;
    wire \uart.timer_Count_6_rep1_RNI02QZ0Z61 ;
    wire \uart.N_145_0 ;
    wire \uart.timer_Count28 ;
    wire \uart.timer_Count28_cascade_ ;
    wire \uart.stateZ0Z_4 ;
    wire \uart.bit_CountZ0Z_1 ;
    wire \uart.bit_CountZ0Z_0 ;
    wire \uart.bit_CountZ0Z_2 ;
    wire \uart.N_175 ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_5_cascade_ ;
    wire \uart.data_Aux_esr_RNO_0Z0Z_6 ;
    wire \uart.state_1_sqmuxa ;
    wire \uart.N_42_0 ;
    wire \uart.N_41_0 ;
    wire \uart.N_37_0 ;
    wire \uart.data_AuxZ0Z_0 ;
    wire data_c_0;
    wire \uart.data_AuxZ0Z_1 ;
    wire data_c_1;
    wire \uart.data_AuxZ0Z_2 ;
    wire data_c_2;
    wire \uart.data_AuxZ0Z_3 ;
    wire data_c_3;
    wire \uart.data_AuxZ0Z_5 ;
    wire data_c_5;
    wire data_c_6;
    wire \uart.data_AuxZ0Z_7 ;
    wire data_c_7;
    wire \uart.data_AuxZ0Z_4 ;
    wire data_c_4;
    wire \uart.state_1_sqmuxa_0 ;
    wire \uart.state_RNIVF8I3Z0Z_4 ;
    wire uart_input_c;
    wire \uart.data_AuxZ0Z_6 ;
    wire _gnd_net_;
    wire clk_system_c_g;
    wire \uart.N_43_0 ;
    wire \uart.un1_state_4_0_a2_iso ;

    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3231),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__3233),
            .DIN(N__3232),
            .DOUT(N__3231),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__3233),
            .PADOUT(N__3232),
            .PADIN(N__3231),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD data_obuf_2_iopad (
            .OE(N__3222),
            .DIN(N__3221),
            .DOUT(N__3220),
            .PACKAGEPIN(data[2]));
    defparam data_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_2_preio (
            .PADOEN(N__3222),
            .PADOUT(N__3221),
            .PADIN(N__3220),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3107),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD data_obuf_6_iopad (
            .OE(N__3213),
            .DIN(N__3212),
            .DOUT(N__3211),
            .PACKAGEPIN(data[6]));
    defparam data_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_6_preio (
            .PADOEN(N__3213),
            .PADOUT(N__3212),
            .PADIN(N__3211),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3032),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_ibuf_iopad (
            .OE(N__3204),
            .DIN(N__3203),
            .DOUT(N__3202),
            .PACKAGEPIN(uart_input));
    defparam uart_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_ibuf_preio (
            .PADOEN(N__3204),
            .PADOUT(N__3203),
            .PADIN(N__3202),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD data_obuf_1_iopad (
            .OE(N__3195),
            .DIN(N__3194),
            .DOUT(N__3193),
            .PACKAGEPIN(data[1]));
    defparam data_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_1_preio (
            .PADOEN(N__3195),
            .PADOUT(N__3194),
            .PADIN(N__3193),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2330),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD data_obuf_5_iopad (
            .OE(N__3186),
            .DIN(N__3185),
            .DOUT(N__3184),
            .PACKAGEPIN(data[5]));
    defparam data_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_5_preio (
            .PADOEN(N__3186),
            .PADOUT(N__3185),
            .PADIN(N__3184),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3047),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam data_obuf_0_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD data_obuf_0_iopad (
            .OE(N__3177),
            .DIN(N__3176),
            .DOUT(N__3175),
            .PACKAGEPIN(data[0]));
    defparam data_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_0_preio (
            .PADOEN(N__3177),
            .PADOUT(N__3176),
            .PADIN(N__3175),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2357),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD data_obuf_4_iopad (
            .OE(N__3168),
            .DIN(N__3167),
            .DOUT(N__3166),
            .PACKAGEPIN(data[4]));
    defparam data_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_4_preio (
            .PADOEN(N__3168),
            .PADOUT(N__3167),
            .PADIN(N__3166),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2972),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam data_rdy_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD data_rdy_obuf_iopad (
            .OE(N__3159),
            .DIN(N__3158),
            .DOUT(N__3157),
            .PACKAGEPIN(data_rdy));
    defparam data_rdy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam data_rdy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO data_rdy_obuf_preio (
            .PADOEN(N__3159),
            .PADOUT(N__3158),
            .PADIN(N__3157),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2309),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD data_obuf_3_iopad (
            .OE(N__3150),
            .DIN(N__3149),
            .DOUT(N__3148),
            .PACKAGEPIN(data[3]));
    defparam data_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_3_preio (
            .PADOEN(N__3150),
            .PADOUT(N__3149),
            .PADIN(N__3148),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3080),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_debug_obuf_iopad (
            .OE(N__3141),
            .DIN(N__3140),
            .DOUT(N__3139),
            .PACKAGEPIN(uart_input_debug));
    defparam uart_input_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_input_debug_obuf_preio (
            .PADOEN(N__3141),
            .PADOUT(N__3140),
            .PADIN(N__3139),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2806),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD data_obuf_7_iopad (
            .OE(N__3132),
            .DIN(N__3131),
            .DOUT(N__3130),
            .PACKAGEPIN(data[7]));
    defparam data_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam data_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO data_obuf_7_preio (
            .PADOEN(N__3132),
            .PADOUT(N__3131),
            .PADIN(N__3130),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2999),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__739 (
            .O(N__3113),
            .I(N__3110));
    LocalMux I__738 (
            .O(N__3110),
            .I(\uart.data_AuxZ0Z_2 ));
    IoInMux I__737 (
            .O(N__3107),
            .I(N__3104));
    LocalMux I__736 (
            .O(N__3104),
            .I(N__3101));
    Span4Mux_s3_v I__735 (
            .O(N__3101),
            .I(N__3098));
    Sp12to4 I__734 (
            .O(N__3098),
            .I(N__3095));
    Span12Mux_s8_h I__733 (
            .O(N__3095),
            .I(N__3092));
    Span12Mux_v I__732 (
            .O(N__3092),
            .I(N__3089));
    Odrv12 I__731 (
            .O(N__3089),
            .I(data_c_2));
    InMux I__730 (
            .O(N__3086),
            .I(N__3083));
    LocalMux I__729 (
            .O(N__3083),
            .I(\uart.data_AuxZ0Z_3 ));
    IoInMux I__728 (
            .O(N__3080),
            .I(N__3077));
    LocalMux I__727 (
            .O(N__3077),
            .I(N__3074));
    Span4Mux_s3_v I__726 (
            .O(N__3074),
            .I(N__3071));
    Span4Mux_h I__725 (
            .O(N__3071),
            .I(N__3068));
    Span4Mux_h I__724 (
            .O(N__3068),
            .I(N__3065));
    Sp12to4 I__723 (
            .O(N__3065),
            .I(N__3062));
    Span12Mux_v I__722 (
            .O(N__3062),
            .I(N__3059));
    Odrv12 I__721 (
            .O(N__3059),
            .I(data_c_3));
    InMux I__720 (
            .O(N__3056),
            .I(N__3053));
    LocalMux I__719 (
            .O(N__3053),
            .I(N__3050));
    Odrv4 I__718 (
            .O(N__3050),
            .I(\uart.data_AuxZ0Z_5 ));
    IoInMux I__717 (
            .O(N__3047),
            .I(N__3044));
    LocalMux I__716 (
            .O(N__3044),
            .I(N__3041));
    Sp12to4 I__715 (
            .O(N__3041),
            .I(N__3038));
    Span12Mux_v I__714 (
            .O(N__3038),
            .I(N__3035));
    Odrv12 I__713 (
            .O(N__3035),
            .I(data_c_5));
    IoInMux I__712 (
            .O(N__3032),
            .I(N__3029));
    LocalMux I__711 (
            .O(N__3029),
            .I(N__3026));
    IoSpan4Mux I__710 (
            .O(N__3026),
            .I(N__3023));
    Span4Mux_s0_v I__709 (
            .O(N__3023),
            .I(N__3020));
    Sp12to4 I__708 (
            .O(N__3020),
            .I(N__3017));
    Span12Mux_v I__707 (
            .O(N__3017),
            .I(N__3014));
    Odrv12 I__706 (
            .O(N__3014),
            .I(data_c_6));
    InMux I__705 (
            .O(N__3011),
            .I(N__3008));
    LocalMux I__704 (
            .O(N__3008),
            .I(N__3005));
    Span4Mux_h I__703 (
            .O(N__3005),
            .I(N__3002));
    Odrv4 I__702 (
            .O(N__3002),
            .I(\uart.data_AuxZ0Z_7 ));
    IoInMux I__701 (
            .O(N__2999),
            .I(N__2996));
    LocalMux I__700 (
            .O(N__2996),
            .I(N__2993));
    IoSpan4Mux I__699 (
            .O(N__2993),
            .I(N__2990));
    Sp12to4 I__698 (
            .O(N__2990),
            .I(N__2987));
    Span12Mux_v I__697 (
            .O(N__2987),
            .I(N__2984));
    Odrv12 I__696 (
            .O(N__2984),
            .I(data_c_7));
    InMux I__695 (
            .O(N__2981),
            .I(N__2978));
    LocalMux I__694 (
            .O(N__2978),
            .I(N__2975));
    Odrv4 I__693 (
            .O(N__2975),
            .I(\uart.data_AuxZ0Z_4 ));
    IoInMux I__692 (
            .O(N__2972),
            .I(N__2969));
    LocalMux I__691 (
            .O(N__2969),
            .I(N__2966));
    Span4Mux_s3_v I__690 (
            .O(N__2966),
            .I(N__2963));
    Span4Mux_v I__689 (
            .O(N__2963),
            .I(N__2960));
    Span4Mux_v I__688 (
            .O(N__2960),
            .I(N__2957));
    Odrv4 I__687 (
            .O(N__2957),
            .I(data_c_4));
    CEMux I__686 (
            .O(N__2954),
            .I(N__2950));
    CEMux I__685 (
            .O(N__2953),
            .I(N__2947));
    LocalMux I__684 (
            .O(N__2950),
            .I(N__2944));
    LocalMux I__683 (
            .O(N__2947),
            .I(N__2941));
    Odrv4 I__682 (
            .O(N__2944),
            .I(\uart.state_1_sqmuxa_0 ));
    Odrv4 I__681 (
            .O(N__2941),
            .I(\uart.state_1_sqmuxa_0 ));
    SRMux I__680 (
            .O(N__2936),
            .I(N__2933));
    LocalMux I__679 (
            .O(N__2933),
            .I(N__2930));
    Span4Mux_v I__678 (
            .O(N__2930),
            .I(N__2926));
    SRMux I__677 (
            .O(N__2929),
            .I(N__2923));
    Sp12to4 I__676 (
            .O(N__2926),
            .I(N__2917));
    LocalMux I__675 (
            .O(N__2923),
            .I(N__2917));
    InMux I__674 (
            .O(N__2922),
            .I(N__2914));
    Odrv12 I__673 (
            .O(N__2917),
            .I(\uart.state_RNIVF8I3Z0Z_4 ));
    LocalMux I__672 (
            .O(N__2914),
            .I(\uart.state_RNIVF8I3Z0Z_4 ));
    InMux I__671 (
            .O(N__2909),
            .I(N__2903));
    InMux I__670 (
            .O(N__2908),
            .I(N__2898));
    InMux I__669 (
            .O(N__2907),
            .I(N__2894));
    InMux I__668 (
            .O(N__2906),
            .I(N__2891));
    LocalMux I__667 (
            .O(N__2903),
            .I(N__2887));
    InMux I__666 (
            .O(N__2902),
            .I(N__2884));
    InMux I__665 (
            .O(N__2901),
            .I(N__2881));
    LocalMux I__664 (
            .O(N__2898),
            .I(N__2878));
    InMux I__663 (
            .O(N__2897),
            .I(N__2875));
    LocalMux I__662 (
            .O(N__2894),
            .I(N__2870));
    LocalMux I__661 (
            .O(N__2891),
            .I(N__2870));
    InMux I__660 (
            .O(N__2890),
            .I(N__2867));
    Span4Mux_h I__659 (
            .O(N__2887),
            .I(N__2859));
    LocalMux I__658 (
            .O(N__2884),
            .I(N__2859));
    LocalMux I__657 (
            .O(N__2881),
            .I(N__2859));
    Span4Mux_v I__656 (
            .O(N__2878),
            .I(N__2851));
    LocalMux I__655 (
            .O(N__2875),
            .I(N__2851));
    Span4Mux_v I__654 (
            .O(N__2870),
            .I(N__2846));
    LocalMux I__653 (
            .O(N__2867),
            .I(N__2846));
    InMux I__652 (
            .O(N__2866),
            .I(N__2843));
    Span4Mux_v I__651 (
            .O(N__2859),
            .I(N__2840));
    InMux I__650 (
            .O(N__2858),
            .I(N__2837));
    InMux I__649 (
            .O(N__2857),
            .I(N__2834));
    InMux I__648 (
            .O(N__2856),
            .I(N__2831));
    Span4Mux_v I__647 (
            .O(N__2851),
            .I(N__2828));
    Span4Mux_v I__646 (
            .O(N__2846),
            .I(N__2825));
    LocalMux I__645 (
            .O(N__2843),
            .I(N__2822));
    Span4Mux_h I__644 (
            .O(N__2840),
            .I(N__2819));
    LocalMux I__643 (
            .O(N__2837),
            .I(N__2812));
    LocalMux I__642 (
            .O(N__2834),
            .I(N__2812));
    LocalMux I__641 (
            .O(N__2831),
            .I(N__2812));
    Sp12to4 I__640 (
            .O(N__2828),
            .I(N__2807));
    Sp12to4 I__639 (
            .O(N__2825),
            .I(N__2807));
    Span12Mux_h I__638 (
            .O(N__2822),
            .I(N__2803));
    Sp12to4 I__637 (
            .O(N__2819),
            .I(N__2798));
    Span12Mux_h I__636 (
            .O(N__2812),
            .I(N__2798));
    Span12Mux_h I__635 (
            .O(N__2807),
            .I(N__2795));
    IoInMux I__634 (
            .O(N__2806),
            .I(N__2792));
    Span12Mux_v I__633 (
            .O(N__2803),
            .I(N__2789));
    Span12Mux_v I__632 (
            .O(N__2798),
            .I(N__2786));
    Span12Mux_v I__631 (
            .O(N__2795),
            .I(N__2783));
    LocalMux I__630 (
            .O(N__2792),
            .I(N__2780));
    Odrv12 I__629 (
            .O(N__2789),
            .I(uart_input_c));
    Odrv12 I__628 (
            .O(N__2786),
            .I(uart_input_c));
    Odrv12 I__627 (
            .O(N__2783),
            .I(uart_input_c));
    Odrv4 I__626 (
            .O(N__2780),
            .I(uart_input_c));
    InMux I__625 (
            .O(N__2771),
            .I(N__2768));
    LocalMux I__624 (
            .O(N__2768),
            .I(N__2765));
    Odrv4 I__623 (
            .O(N__2765),
            .I(\uart.data_AuxZ0Z_6 ));
    ClkMux I__622 (
            .O(N__2762),
            .I(N__2702));
    ClkMux I__621 (
            .O(N__2761),
            .I(N__2702));
    ClkMux I__620 (
            .O(N__2760),
            .I(N__2702));
    ClkMux I__619 (
            .O(N__2759),
            .I(N__2702));
    ClkMux I__618 (
            .O(N__2758),
            .I(N__2702));
    ClkMux I__617 (
            .O(N__2757),
            .I(N__2702));
    ClkMux I__616 (
            .O(N__2756),
            .I(N__2702));
    ClkMux I__615 (
            .O(N__2755),
            .I(N__2702));
    ClkMux I__614 (
            .O(N__2754),
            .I(N__2702));
    ClkMux I__613 (
            .O(N__2753),
            .I(N__2702));
    ClkMux I__612 (
            .O(N__2752),
            .I(N__2702));
    ClkMux I__611 (
            .O(N__2751),
            .I(N__2702));
    ClkMux I__610 (
            .O(N__2750),
            .I(N__2702));
    ClkMux I__609 (
            .O(N__2749),
            .I(N__2702));
    ClkMux I__608 (
            .O(N__2748),
            .I(N__2702));
    ClkMux I__607 (
            .O(N__2747),
            .I(N__2702));
    ClkMux I__606 (
            .O(N__2746),
            .I(N__2702));
    ClkMux I__605 (
            .O(N__2745),
            .I(N__2702));
    ClkMux I__604 (
            .O(N__2744),
            .I(N__2702));
    ClkMux I__603 (
            .O(N__2743),
            .I(N__2702));
    GlobalMux I__602 (
            .O(N__2702),
            .I(N__2699));
    gio2CtrlBuf I__601 (
            .O(N__2699),
            .I(clk_system_c_g));
    CEMux I__600 (
            .O(N__2696),
            .I(N__2693));
    LocalMux I__599 (
            .O(N__2693),
            .I(N__2690));
    Span4Mux_h I__598 (
            .O(N__2690),
            .I(N__2687));
    Odrv4 I__597 (
            .O(N__2687),
            .I(\uart.N_43_0 ));
    SRMux I__596 (
            .O(N__2684),
            .I(N__2680));
    SRMux I__595 (
            .O(N__2683),
            .I(N__2677));
    LocalMux I__594 (
            .O(N__2680),
            .I(N__2670));
    LocalMux I__593 (
            .O(N__2677),
            .I(N__2670));
    SRMux I__592 (
            .O(N__2676),
            .I(N__2667));
    SRMux I__591 (
            .O(N__2675),
            .I(N__2664));
    Span4Mux_v I__590 (
            .O(N__2670),
            .I(N__2654));
    LocalMux I__589 (
            .O(N__2667),
            .I(N__2654));
    LocalMux I__588 (
            .O(N__2664),
            .I(N__2651));
    InMux I__587 (
            .O(N__2663),
            .I(N__2640));
    InMux I__586 (
            .O(N__2662),
            .I(N__2640));
    InMux I__585 (
            .O(N__2661),
            .I(N__2635));
    InMux I__584 (
            .O(N__2660),
            .I(N__2635));
    SRMux I__583 (
            .O(N__2659),
            .I(N__2632));
    Span4Mux_v I__582 (
            .O(N__2654),
            .I(N__2627));
    Span4Mux_h I__581 (
            .O(N__2651),
            .I(N__2627));
    SRMux I__580 (
            .O(N__2650),
            .I(N__2624));
    SRMux I__579 (
            .O(N__2649),
            .I(N__2621));
    InMux I__578 (
            .O(N__2648),
            .I(N__2616));
    InMux I__577 (
            .O(N__2647),
            .I(N__2616));
    SRMux I__576 (
            .O(N__2646),
            .I(N__2611));
    InMux I__575 (
            .O(N__2645),
            .I(N__2611));
    LocalMux I__574 (
            .O(N__2640),
            .I(N__2606));
    LocalMux I__573 (
            .O(N__2635),
            .I(N__2606));
    LocalMux I__572 (
            .O(N__2632),
            .I(\uart.un1_state_4_0_a2_iso ));
    Odrv4 I__571 (
            .O(N__2627),
            .I(\uart.un1_state_4_0_a2_iso ));
    LocalMux I__570 (
            .O(N__2624),
            .I(\uart.un1_state_4_0_a2_iso ));
    LocalMux I__569 (
            .O(N__2621),
            .I(\uart.un1_state_4_0_a2_iso ));
    LocalMux I__568 (
            .O(N__2616),
            .I(\uart.un1_state_4_0_a2_iso ));
    LocalMux I__567 (
            .O(N__2611),
            .I(\uart.un1_state_4_0_a2_iso ));
    Odrv4 I__566 (
            .O(N__2606),
            .I(\uart.un1_state_4_0_a2_iso ));
    InMux I__565 (
            .O(N__2591),
            .I(N__2588));
    LocalMux I__564 (
            .O(N__2588),
            .I(N__2582));
    InMux I__563 (
            .O(N__2587),
            .I(N__2577));
    InMux I__562 (
            .O(N__2586),
            .I(N__2567));
    InMux I__561 (
            .O(N__2585),
            .I(N__2564));
    Span4Mux_v I__560 (
            .O(N__2582),
            .I(N__2561));
    InMux I__559 (
            .O(N__2581),
            .I(N__2556));
    InMux I__558 (
            .O(N__2580),
            .I(N__2556));
    LocalMux I__557 (
            .O(N__2577),
            .I(N__2553));
    InMux I__556 (
            .O(N__2576),
            .I(N__2546));
    InMux I__555 (
            .O(N__2575),
            .I(N__2546));
    InMux I__554 (
            .O(N__2574),
            .I(N__2546));
    InMux I__553 (
            .O(N__2573),
            .I(N__2541));
    InMux I__552 (
            .O(N__2572),
            .I(N__2541));
    InMux I__551 (
            .O(N__2571),
            .I(N__2536));
    InMux I__550 (
            .O(N__2570),
            .I(N__2536));
    LocalMux I__549 (
            .O(N__2567),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__548 (
            .O(N__2564),
            .I(\uart.bit_CountZ0Z_0 ));
    Odrv4 I__547 (
            .O(N__2561),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__546 (
            .O(N__2556),
            .I(\uart.bit_CountZ0Z_0 ));
    Odrv4 I__545 (
            .O(N__2553),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__544 (
            .O(N__2546),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__543 (
            .O(N__2541),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__542 (
            .O(N__2536),
            .I(\uart.bit_CountZ0Z_0 ));
    CascadeMux I__541 (
            .O(N__2519),
            .I(N__2514));
    CascadeMux I__540 (
            .O(N__2518),
            .I(N__2511));
    InMux I__539 (
            .O(N__2517),
            .I(N__2503));
    InMux I__538 (
            .O(N__2514),
            .I(N__2503));
    InMux I__537 (
            .O(N__2511),
            .I(N__2500));
    CascadeMux I__536 (
            .O(N__2510),
            .I(N__2497));
    CascadeMux I__535 (
            .O(N__2509),
            .I(N__2494));
    CascadeMux I__534 (
            .O(N__2508),
            .I(N__2491));
    LocalMux I__533 (
            .O(N__2503),
            .I(N__2485));
    LocalMux I__532 (
            .O(N__2500),
            .I(N__2482));
    InMux I__531 (
            .O(N__2497),
            .I(N__2479));
    InMux I__530 (
            .O(N__2494),
            .I(N__2472));
    InMux I__529 (
            .O(N__2491),
            .I(N__2472));
    InMux I__528 (
            .O(N__2490),
            .I(N__2472));
    CascadeMux I__527 (
            .O(N__2489),
            .I(N__2469));
    InMux I__526 (
            .O(N__2488),
            .I(N__2465));
    Span4Mux_h I__525 (
            .O(N__2485),
            .I(N__2462));
    Span4Mux_v I__524 (
            .O(N__2482),
            .I(N__2455));
    LocalMux I__523 (
            .O(N__2479),
            .I(N__2455));
    LocalMux I__522 (
            .O(N__2472),
            .I(N__2455));
    InMux I__521 (
            .O(N__2469),
            .I(N__2452));
    InMux I__520 (
            .O(N__2468),
            .I(N__2449));
    LocalMux I__519 (
            .O(N__2465),
            .I(\uart.bit_CountZ0Z_2 ));
    Odrv4 I__518 (
            .O(N__2462),
            .I(\uart.bit_CountZ0Z_2 ));
    Odrv4 I__517 (
            .O(N__2455),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__516 (
            .O(N__2452),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__515 (
            .O(N__2449),
            .I(\uart.bit_CountZ0Z_2 ));
    CascadeMux I__514 (
            .O(N__2438),
            .I(N__2430));
    InMux I__513 (
            .O(N__2437),
            .I(N__2426));
    InMux I__512 (
            .O(N__2436),
            .I(N__2423));
    InMux I__511 (
            .O(N__2435),
            .I(N__2418));
    InMux I__510 (
            .O(N__2434),
            .I(N__2418));
    InMux I__509 (
            .O(N__2433),
            .I(N__2415));
    InMux I__508 (
            .O(N__2430),
            .I(N__2410));
    InMux I__507 (
            .O(N__2429),
            .I(N__2410));
    LocalMux I__506 (
            .O(N__2426),
            .I(\uart.N_175 ));
    LocalMux I__505 (
            .O(N__2423),
            .I(\uart.N_175 ));
    LocalMux I__504 (
            .O(N__2418),
            .I(\uart.N_175 ));
    LocalMux I__503 (
            .O(N__2415),
            .I(\uart.N_175 ));
    LocalMux I__502 (
            .O(N__2410),
            .I(\uart.N_175 ));
    CascadeMux I__501 (
            .O(N__2399),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_5_cascade_ ));
    InMux I__500 (
            .O(N__2396),
            .I(N__2393));
    LocalMux I__499 (
            .O(N__2393),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_6 ));
    InMux I__498 (
            .O(N__2390),
            .I(N__2387));
    LocalMux I__497 (
            .O(N__2387),
            .I(\uart.state_1_sqmuxa ));
    CEMux I__496 (
            .O(N__2384),
            .I(N__2381));
    LocalMux I__495 (
            .O(N__2381),
            .I(\uart.N_42_0 ));
    CEMux I__494 (
            .O(N__2378),
            .I(N__2375));
    LocalMux I__493 (
            .O(N__2375),
            .I(N__2372));
    Odrv4 I__492 (
            .O(N__2372),
            .I(\uart.N_41_0 ));
    CEMux I__491 (
            .O(N__2369),
            .I(N__2366));
    LocalMux I__490 (
            .O(N__2366),
            .I(\uart.N_37_0 ));
    InMux I__489 (
            .O(N__2363),
            .I(N__2360));
    LocalMux I__488 (
            .O(N__2360),
            .I(\uart.data_AuxZ0Z_0 ));
    IoInMux I__487 (
            .O(N__2357),
            .I(N__2354));
    LocalMux I__486 (
            .O(N__2354),
            .I(N__2351));
    Span12Mux_s5_v I__485 (
            .O(N__2351),
            .I(N__2348));
    Span12Mux_v I__484 (
            .O(N__2348),
            .I(N__2345));
    Odrv12 I__483 (
            .O(N__2345),
            .I(data_c_0));
    InMux I__482 (
            .O(N__2342),
            .I(N__2339));
    LocalMux I__481 (
            .O(N__2339),
            .I(N__2336));
    Span4Mux_v I__480 (
            .O(N__2336),
            .I(N__2333));
    Odrv4 I__479 (
            .O(N__2333),
            .I(\uart.data_AuxZ0Z_1 ));
    IoInMux I__478 (
            .O(N__2330),
            .I(N__2327));
    LocalMux I__477 (
            .O(N__2327),
            .I(N__2324));
    IoSpan4Mux I__476 (
            .O(N__2324),
            .I(N__2321));
    Span4Mux_s3_v I__475 (
            .O(N__2321),
            .I(N__2318));
    Sp12to4 I__474 (
            .O(N__2318),
            .I(N__2315));
    Span12Mux_v I__473 (
            .O(N__2315),
            .I(N__2312));
    Odrv12 I__472 (
            .O(N__2312),
            .I(data_c_1));
    IoInMux I__471 (
            .O(N__2309),
            .I(N__2306));
    LocalMux I__470 (
            .O(N__2306),
            .I(N__2303));
    IoSpan4Mux I__469 (
            .O(N__2303),
            .I(N__2300));
    Span4Mux_s3_v I__468 (
            .O(N__2300),
            .I(N__2297));
    Sp12to4 I__467 (
            .O(N__2297),
            .I(N__2294));
    Odrv12 I__466 (
            .O(N__2294),
            .I(data_rdy_c));
    InMux I__465 (
            .O(N__2291),
            .I(N__2288));
    LocalMux I__464 (
            .O(N__2288),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_0 ));
    InMux I__463 (
            .O(N__2285),
            .I(N__2282));
    LocalMux I__462 (
            .O(N__2282),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_4 ));
    CEMux I__461 (
            .O(N__2279),
            .I(N__2276));
    LocalMux I__460 (
            .O(N__2276),
            .I(N__2273));
    Odrv4 I__459 (
            .O(N__2273),
            .I(\uart.N_39_0 ));
    CEMux I__458 (
            .O(N__2270),
            .I(N__2267));
    LocalMux I__457 (
            .O(N__2267),
            .I(N__2264));
    Odrv4 I__456 (
            .O(N__2264),
            .I(\uart.N_40_0 ));
    InMux I__455 (
            .O(N__2261),
            .I(N__2258));
    LocalMux I__454 (
            .O(N__2258),
            .I(\uart.timer_Count_6_rep1_RNI1B4SZ0 ));
    InMux I__453 (
            .O(N__2255),
            .I(N__2252));
    LocalMux I__452 (
            .O(N__2252),
            .I(\uart.timer_Count_6_rep1_RNI02QZ0Z61 ));
    InMux I__451 (
            .O(N__2249),
            .I(N__2245));
    InMux I__450 (
            .O(N__2248),
            .I(N__2242));
    LocalMux I__449 (
            .O(N__2245),
            .I(\uart.N_145_0 ));
    LocalMux I__448 (
            .O(N__2242),
            .I(\uart.N_145_0 ));
    InMux I__447 (
            .O(N__2237),
            .I(N__2232));
    InMux I__446 (
            .O(N__2236),
            .I(N__2229));
    InMux I__445 (
            .O(N__2235),
            .I(N__2226));
    LocalMux I__444 (
            .O(N__2232),
            .I(N__2223));
    LocalMux I__443 (
            .O(N__2229),
            .I(N__2220));
    LocalMux I__442 (
            .O(N__2226),
            .I(\uart.timer_Count28 ));
    Odrv4 I__441 (
            .O(N__2223),
            .I(\uart.timer_Count28 ));
    Odrv12 I__440 (
            .O(N__2220),
            .I(\uart.timer_Count28 ));
    CascadeMux I__439 (
            .O(N__2213),
            .I(\uart.timer_Count28_cascade_ ));
    InMux I__438 (
            .O(N__2210),
            .I(N__2206));
    InMux I__437 (
            .O(N__2209),
            .I(N__2196));
    LocalMux I__436 (
            .O(N__2206),
            .I(N__2193));
    InMux I__435 (
            .O(N__2205),
            .I(N__2186));
    InMux I__434 (
            .O(N__2204),
            .I(N__2186));
    InMux I__433 (
            .O(N__2203),
            .I(N__2186));
    InMux I__432 (
            .O(N__2202),
            .I(N__2179));
    InMux I__431 (
            .O(N__2201),
            .I(N__2179));
    InMux I__430 (
            .O(N__2200),
            .I(N__2179));
    InMux I__429 (
            .O(N__2199),
            .I(N__2171));
    LocalMux I__428 (
            .O(N__2196),
            .I(N__2168));
    Span4Mux_v I__427 (
            .O(N__2193),
            .I(N__2161));
    LocalMux I__426 (
            .O(N__2186),
            .I(N__2161));
    LocalMux I__425 (
            .O(N__2179),
            .I(N__2161));
    InMux I__424 (
            .O(N__2178),
            .I(N__2158));
    InMux I__423 (
            .O(N__2177),
            .I(N__2155));
    InMux I__422 (
            .O(N__2176),
            .I(N__2148));
    InMux I__421 (
            .O(N__2175),
            .I(N__2148));
    InMux I__420 (
            .O(N__2174),
            .I(N__2148));
    LocalMux I__419 (
            .O(N__2171),
            .I(\uart.stateZ0Z_4 ));
    Odrv12 I__418 (
            .O(N__2168),
            .I(\uart.stateZ0Z_4 ));
    Odrv4 I__417 (
            .O(N__2161),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__416 (
            .O(N__2158),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__415 (
            .O(N__2155),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__414 (
            .O(N__2148),
            .I(\uart.stateZ0Z_4 ));
    InMux I__413 (
            .O(N__2135),
            .I(N__2127));
    InMux I__412 (
            .O(N__2134),
            .I(N__2124));
    InMux I__411 (
            .O(N__2133),
            .I(N__2117));
    InMux I__410 (
            .O(N__2132),
            .I(N__2117));
    InMux I__409 (
            .O(N__2131),
            .I(N__2117));
    InMux I__408 (
            .O(N__2130),
            .I(N__2111));
    LocalMux I__407 (
            .O(N__2127),
            .I(N__2104));
    LocalMux I__406 (
            .O(N__2124),
            .I(N__2104));
    LocalMux I__405 (
            .O(N__2117),
            .I(N__2104));
    InMux I__404 (
            .O(N__2116),
            .I(N__2099));
    InMux I__403 (
            .O(N__2115),
            .I(N__2099));
    InMux I__402 (
            .O(N__2114),
            .I(N__2093));
    LocalMux I__401 (
            .O(N__2111),
            .I(N__2086));
    Span4Mux_v I__400 (
            .O(N__2104),
            .I(N__2086));
    LocalMux I__399 (
            .O(N__2099),
            .I(N__2086));
    InMux I__398 (
            .O(N__2098),
            .I(N__2081));
    InMux I__397 (
            .O(N__2097),
            .I(N__2081));
    InMux I__396 (
            .O(N__2096),
            .I(N__2078));
    LocalMux I__395 (
            .O(N__2093),
            .I(\uart.bit_CountZ0Z_1 ));
    Odrv4 I__394 (
            .O(N__2086),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__393 (
            .O(N__2081),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__392 (
            .O(N__2078),
            .I(\uart.bit_CountZ0Z_1 ));
    CascadeMux I__391 (
            .O(N__2069),
            .I(N__2065));
    InMux I__390 (
            .O(N__2068),
            .I(N__2057));
    InMux I__389 (
            .O(N__2065),
            .I(N__2057));
    InMux I__388 (
            .O(N__2064),
            .I(N__2057));
    LocalMux I__387 (
            .O(N__2057),
            .I(\uart.un4_timer_Count_1_c2 ));
    CascadeMux I__386 (
            .O(N__2054),
            .I(\uart.timer_Count_RNIMLMA1Z0Z_1_cascade_ ));
    InMux I__385 (
            .O(N__2051),
            .I(N__2039));
    InMux I__384 (
            .O(N__2050),
            .I(N__2039));
    InMux I__383 (
            .O(N__2049),
            .I(N__2039));
    InMux I__382 (
            .O(N__2048),
            .I(N__2039));
    LocalMux I__381 (
            .O(N__2039),
            .I(\uart.un4_timer_Count_1_c5 ));
    CascadeMux I__380 (
            .O(N__2036),
            .I(\uart.un4_timer_Count_1_c5_cascade_ ));
    InMux I__379 (
            .O(N__2033),
            .I(N__2028));
    CascadeMux I__378 (
            .O(N__2032),
            .I(N__2024));
    CascadeMux I__377 (
            .O(N__2031),
            .I(N__2019));
    LocalMux I__376 (
            .O(N__2028),
            .I(N__2014));
    InMux I__375 (
            .O(N__2027),
            .I(N__2009));
    InMux I__374 (
            .O(N__2024),
            .I(N__2009));
    InMux I__373 (
            .O(N__2023),
            .I(N__2006));
    InMux I__372 (
            .O(N__2022),
            .I(N__2003));
    InMux I__371 (
            .O(N__2019),
            .I(N__1996));
    InMux I__370 (
            .O(N__2018),
            .I(N__1996));
    InMux I__369 (
            .O(N__2017),
            .I(N__1996));
    Odrv4 I__368 (
            .O(N__2014),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__367 (
            .O(N__2009),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__366 (
            .O(N__2006),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__365 (
            .O(N__2003),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__364 (
            .O(N__1996),
            .I(\uart.timer_CountZ0Z_3 ));
    InMux I__363 (
            .O(N__1985),
            .I(N__1982));
    LocalMux I__362 (
            .O(N__1982),
            .I(N__1971));
    InMux I__361 (
            .O(N__1981),
            .I(N__1966));
    InMux I__360 (
            .O(N__1980),
            .I(N__1966));
    InMux I__359 (
            .O(N__1979),
            .I(N__1963));
    InMux I__358 (
            .O(N__1978),
            .I(N__1960));
    InMux I__357 (
            .O(N__1977),
            .I(N__1951));
    InMux I__356 (
            .O(N__1976),
            .I(N__1951));
    InMux I__355 (
            .O(N__1975),
            .I(N__1951));
    InMux I__354 (
            .O(N__1974),
            .I(N__1951));
    Odrv4 I__353 (
            .O(N__1971),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__352 (
            .O(N__1966),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__351 (
            .O(N__1963),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__350 (
            .O(N__1960),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__349 (
            .O(N__1951),
            .I(\uart.timer_CountZ0Z_2 ));
    CascadeMux I__348 (
            .O(N__1940),
            .I(N__1928));
    InMux I__347 (
            .O(N__1939),
            .I(N__1924));
    CascadeMux I__346 (
            .O(N__1938),
            .I(N__1920));
    CascadeMux I__345 (
            .O(N__1937),
            .I(N__1917));
    CascadeMux I__344 (
            .O(N__1936),
            .I(N__1914));
    InMux I__343 (
            .O(N__1935),
            .I(N__1911));
    InMux I__342 (
            .O(N__1934),
            .I(N__1904));
    InMux I__341 (
            .O(N__1933),
            .I(N__1904));
    InMux I__340 (
            .O(N__1932),
            .I(N__1904));
    CascadeMux I__339 (
            .O(N__1931),
            .I(N__1901));
    InMux I__338 (
            .O(N__1928),
            .I(N__1897));
    InMux I__337 (
            .O(N__1927),
            .I(N__1894));
    LocalMux I__336 (
            .O(N__1924),
            .I(N__1891));
    InMux I__335 (
            .O(N__1923),
            .I(N__1884));
    InMux I__334 (
            .O(N__1920),
            .I(N__1884));
    InMux I__333 (
            .O(N__1917),
            .I(N__1884));
    InMux I__332 (
            .O(N__1914),
            .I(N__1881));
    LocalMux I__331 (
            .O(N__1911),
            .I(N__1876));
    LocalMux I__330 (
            .O(N__1904),
            .I(N__1876));
    InMux I__329 (
            .O(N__1901),
            .I(N__1871));
    InMux I__328 (
            .O(N__1900),
            .I(N__1871));
    LocalMux I__327 (
            .O(N__1897),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__326 (
            .O(N__1894),
            .I(\uart.stateZ0Z_3 ));
    Odrv4 I__325 (
            .O(N__1891),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__324 (
            .O(N__1884),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__323 (
            .O(N__1881),
            .I(\uart.stateZ0Z_3 ));
    Odrv4 I__322 (
            .O(N__1876),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__321 (
            .O(N__1871),
            .I(\uart.stateZ0Z_3 ));
    CascadeMux I__320 (
            .O(N__1856),
            .I(\uart.timer_Count_RNIHJ661Z0Z_3_cascade_ ));
    InMux I__319 (
            .O(N__1853),
            .I(N__1847));
    InMux I__318 (
            .O(N__1852),
            .I(N__1847));
    LocalMux I__317 (
            .O(N__1847),
            .I(N__1839));
    InMux I__316 (
            .O(N__1846),
            .I(N__1833));
    InMux I__315 (
            .O(N__1845),
            .I(N__1819));
    InMux I__314 (
            .O(N__1844),
            .I(N__1819));
    InMux I__313 (
            .O(N__1843),
            .I(N__1819));
    InMux I__312 (
            .O(N__1842),
            .I(N__1819));
    Span4Mux_h I__311 (
            .O(N__1839),
            .I(N__1816));
    InMux I__310 (
            .O(N__1838),
            .I(N__1809));
    InMux I__309 (
            .O(N__1837),
            .I(N__1809));
    InMux I__308 (
            .O(N__1836),
            .I(N__1809));
    LocalMux I__307 (
            .O(N__1833),
            .I(N__1806));
    InMux I__306 (
            .O(N__1832),
            .I(N__1799));
    InMux I__305 (
            .O(N__1831),
            .I(N__1799));
    InMux I__304 (
            .O(N__1830),
            .I(N__1799));
    InMux I__303 (
            .O(N__1829),
            .I(N__1794));
    InMux I__302 (
            .O(N__1828),
            .I(N__1794));
    LocalMux I__301 (
            .O(N__1819),
            .I(\uart.timer_CountZ0Z_5 ));
    Odrv4 I__300 (
            .O(N__1816),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__299 (
            .O(N__1809),
            .I(\uart.timer_CountZ0Z_5 ));
    Odrv4 I__298 (
            .O(N__1806),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__297 (
            .O(N__1799),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__296 (
            .O(N__1794),
            .I(\uart.timer_CountZ0Z_5 ));
    InMux I__295 (
            .O(N__1781),
            .I(N__1776));
    InMux I__294 (
            .O(N__1780),
            .I(N__1773));
    InMux I__293 (
            .O(N__1779),
            .I(N__1770));
    LocalMux I__292 (
            .O(N__1776),
            .I(N__1767));
    LocalMux I__291 (
            .O(N__1773),
            .I(N__1762));
    LocalMux I__290 (
            .O(N__1770),
            .I(N__1762));
    Span4Mux_h I__289 (
            .O(N__1767),
            .I(N__1759));
    Span4Mux_v I__288 (
            .O(N__1762),
            .I(N__1756));
    Odrv4 I__287 (
            .O(N__1759),
            .I(\uart.state_0_sqmuxa_1_d ));
    Odrv4 I__286 (
            .O(N__1756),
            .I(\uart.state_0_sqmuxa_1_d ));
    InMux I__285 (
            .O(N__1751),
            .I(N__1744));
    InMux I__284 (
            .O(N__1750),
            .I(N__1739));
    InMux I__283 (
            .O(N__1749),
            .I(N__1739));
    InMux I__282 (
            .O(N__1748),
            .I(N__1734));
    InMux I__281 (
            .O(N__1747),
            .I(N__1734));
    LocalMux I__280 (
            .O(N__1744),
            .I(\uart.timer_CountZ0Z_0 ));
    LocalMux I__279 (
            .O(N__1739),
            .I(\uart.timer_CountZ0Z_0 ));
    LocalMux I__278 (
            .O(N__1734),
            .I(\uart.timer_CountZ0Z_0 ));
    InMux I__277 (
            .O(N__1727),
            .I(N__1718));
    InMux I__276 (
            .O(N__1726),
            .I(N__1718));
    InMux I__275 (
            .O(N__1725),
            .I(N__1713));
    InMux I__274 (
            .O(N__1724),
            .I(N__1713));
    InMux I__273 (
            .O(N__1723),
            .I(N__1710));
    LocalMux I__272 (
            .O(N__1718),
            .I(\uart.timer_CountZ0Z_1 ));
    LocalMux I__271 (
            .O(N__1713),
            .I(\uart.timer_CountZ0Z_1 ));
    LocalMux I__270 (
            .O(N__1710),
            .I(\uart.timer_CountZ0Z_1 ));
    SRMux I__269 (
            .O(N__1703),
            .I(N__1699));
    SRMux I__268 (
            .O(N__1702),
            .I(N__1696));
    LocalMux I__267 (
            .O(N__1699),
            .I(N__1693));
    LocalMux I__266 (
            .O(N__1696),
            .I(N__1689));
    Span4Mux_h I__265 (
            .O(N__1693),
            .I(N__1686));
    SRMux I__264 (
            .O(N__1692),
            .I(N__1683));
    Span4Mux_v I__263 (
            .O(N__1689),
            .I(N__1680));
    Sp12to4 I__262 (
            .O(N__1686),
            .I(N__1675));
    LocalMux I__261 (
            .O(N__1683),
            .I(N__1675));
    Odrv4 I__260 (
            .O(N__1680),
            .I(\uart.un1_timer_Count_0_sqmuxa_0 ));
    Odrv12 I__259 (
            .O(N__1675),
            .I(\uart.un1_timer_Count_0_sqmuxa_0 ));
    CascadeMux I__258 (
            .O(N__1670),
            .I(N__1667));
    InMux I__257 (
            .O(N__1667),
            .I(N__1661));
    CascadeMux I__256 (
            .O(N__1666),
            .I(N__1654));
    CascadeMux I__255 (
            .O(N__1665),
            .I(N__1651));
    InMux I__254 (
            .O(N__1664),
            .I(N__1648));
    LocalMux I__253 (
            .O(N__1661),
            .I(N__1645));
    InMux I__252 (
            .O(N__1660),
            .I(N__1638));
    InMux I__251 (
            .O(N__1659),
            .I(N__1638));
    InMux I__250 (
            .O(N__1658),
            .I(N__1638));
    InMux I__249 (
            .O(N__1657),
            .I(N__1635));
    InMux I__248 (
            .O(N__1654),
            .I(N__1632));
    InMux I__247 (
            .O(N__1651),
            .I(N__1629));
    LocalMux I__246 (
            .O(N__1648),
            .I(\uart.timer_CountZ0Z_4 ));
    Odrv12 I__245 (
            .O(N__1645),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__244 (
            .O(N__1638),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__243 (
            .O(N__1635),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__242 (
            .O(N__1632),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__241 (
            .O(N__1629),
            .I(\uart.timer_CountZ0Z_4 ));
    CascadeMux I__240 (
            .O(N__1616),
            .I(N__1612));
    InMux I__239 (
            .O(N__1615),
            .I(N__1599));
    InMux I__238 (
            .O(N__1612),
            .I(N__1599));
    InMux I__237 (
            .O(N__1611),
            .I(N__1592));
    InMux I__236 (
            .O(N__1610),
            .I(N__1592));
    InMux I__235 (
            .O(N__1609),
            .I(N__1592));
    InMux I__234 (
            .O(N__1608),
            .I(N__1585));
    InMux I__233 (
            .O(N__1607),
            .I(N__1582));
    InMux I__232 (
            .O(N__1606),
            .I(N__1575));
    InMux I__231 (
            .O(N__1605),
            .I(N__1575));
    InMux I__230 (
            .O(N__1604),
            .I(N__1575));
    LocalMux I__229 (
            .O(N__1599),
            .I(N__1570));
    LocalMux I__228 (
            .O(N__1592),
            .I(N__1570));
    InMux I__227 (
            .O(N__1591),
            .I(N__1565));
    InMux I__226 (
            .O(N__1590),
            .I(N__1565));
    InMux I__225 (
            .O(N__1589),
            .I(N__1560));
    InMux I__224 (
            .O(N__1588),
            .I(N__1560));
    LocalMux I__223 (
            .O(N__1585),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__222 (
            .O(N__1582),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__221 (
            .O(N__1575),
            .I(\uart.timer_CountZ0Z_7 ));
    Odrv4 I__220 (
            .O(N__1570),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__219 (
            .O(N__1565),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__218 (
            .O(N__1560),
            .I(\uart.timer_CountZ0Z_7 ));
    CascadeMux I__217 (
            .O(N__1547),
            .I(N__1544));
    InMux I__216 (
            .O(N__1544),
            .I(N__1541));
    LocalMux I__215 (
            .O(N__1541),
            .I(\uart.N_28_mux_i_i_0 ));
    InMux I__214 (
            .O(N__1538),
            .I(N__1535));
    LocalMux I__213 (
            .O(N__1535),
            .I(\uart.N_22_mux ));
    CascadeMux I__212 (
            .O(N__1532),
            .I(\uart.N_175_cascade_ ));
    InMux I__211 (
            .O(N__1529),
            .I(N__1526));
    LocalMux I__210 (
            .O(N__1526),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_1 ));
    CascadeMux I__209 (
            .O(N__1523),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__208 (
            .O(N__1520),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_2_cascade_ ));
    InMux I__207 (
            .O(N__1517),
            .I(N__1512));
    InMux I__206 (
            .O(N__1516),
            .I(N__1509));
    InMux I__205 (
            .O(N__1515),
            .I(N__1503));
    LocalMux I__204 (
            .O(N__1512),
            .I(N__1500));
    LocalMux I__203 (
            .O(N__1509),
            .I(N__1497));
    InMux I__202 (
            .O(N__1508),
            .I(N__1494));
    InMux I__201 (
            .O(N__1507),
            .I(N__1489));
    InMux I__200 (
            .O(N__1506),
            .I(N__1489));
    LocalMux I__199 (
            .O(N__1503),
            .I(\uart.timer_Count_6_repZ0Z1 ));
    Odrv4 I__198 (
            .O(N__1500),
            .I(\uart.timer_Count_6_repZ0Z1 ));
    Odrv4 I__197 (
            .O(N__1497),
            .I(\uart.timer_Count_6_repZ0Z1 ));
    LocalMux I__196 (
            .O(N__1494),
            .I(\uart.timer_Count_6_repZ0Z1 ));
    LocalMux I__195 (
            .O(N__1489),
            .I(\uart.timer_Count_6_repZ0Z1 ));
    CascadeMux I__194 (
            .O(N__1478),
            .I(N__1473));
    InMux I__193 (
            .O(N__1477),
            .I(N__1470));
    InMux I__192 (
            .O(N__1476),
            .I(N__1467));
    InMux I__191 (
            .O(N__1473),
            .I(N__1464));
    LocalMux I__190 (
            .O(N__1470),
            .I(\uart.timer_Count_fastZ0Z_6 ));
    LocalMux I__189 (
            .O(N__1467),
            .I(\uart.timer_Count_fastZ0Z_6 ));
    LocalMux I__188 (
            .O(N__1464),
            .I(\uart.timer_Count_fastZ0Z_6 ));
    CascadeMux I__187 (
            .O(N__1457),
            .I(\uart.un1_state_4_0_a2_iso_cascade_ ));
    CEMux I__186 (
            .O(N__1454),
            .I(N__1451));
    LocalMux I__185 (
            .O(N__1451),
            .I(N__1448));
    Span4Mux_h I__184 (
            .O(N__1448),
            .I(N__1445));
    Odrv4 I__183 (
            .O(N__1445),
            .I(\uart.N_38_0 ));
    InMux I__182 (
            .O(N__1442),
            .I(N__1438));
    InMux I__181 (
            .O(N__1441),
            .I(N__1435));
    LocalMux I__180 (
            .O(N__1438),
            .I(\uart.N_165_1 ));
    LocalMux I__179 (
            .O(N__1435),
            .I(\uart.N_165_1 ));
    InMux I__178 (
            .O(N__1430),
            .I(N__1427));
    LocalMux I__177 (
            .O(N__1427),
            .I(\uart.timer_Count_RNIICSG1Z0Z_6 ));
    InMux I__176 (
            .O(N__1424),
            .I(N__1421));
    LocalMux I__175 (
            .O(N__1421),
            .I(\uart.state_RNO_0Z0Z_3 ));
    CascadeMux I__174 (
            .O(N__1418),
            .I(N__1415));
    InMux I__173 (
            .O(N__1415),
            .I(N__1412));
    LocalMux I__172 (
            .O(N__1412),
            .I(N__1409));
    Odrv4 I__171 (
            .O(N__1409),
            .I(\uart.state_RNO_1Z0Z_3 ));
    CascadeMux I__170 (
            .O(N__1406),
            .I(N__1403));
    InMux I__169 (
            .O(N__1403),
            .I(N__1399));
    InMux I__168 (
            .O(N__1402),
            .I(N__1396));
    LocalMux I__167 (
            .O(N__1399),
            .I(N__1393));
    LocalMux I__166 (
            .O(N__1396),
            .I(\uart.N_147_0 ));
    Odrv4 I__165 (
            .O(N__1393),
            .I(\uart.N_147_0 ));
    InMux I__164 (
            .O(N__1388),
            .I(N__1385));
    LocalMux I__163 (
            .O(N__1385),
            .I(N__1382));
    Odrv4 I__162 (
            .O(N__1382),
            .I(\uart.N_159 ));
    CascadeMux I__161 (
            .O(N__1379),
            .I(\uart.timer_Count_6_rep1_RNIRC5SZ0Z1_cascade_ ));
    CascadeMux I__160 (
            .O(N__1376),
            .I(\uart.un1_state_2_0_a3_0_cascade_ ));
    CascadeMux I__159 (
            .O(N__1373),
            .I(N__1367));
    InMux I__158 (
            .O(N__1372),
            .I(N__1361));
    InMux I__157 (
            .O(N__1371),
            .I(N__1356));
    InMux I__156 (
            .O(N__1370),
            .I(N__1356));
    InMux I__155 (
            .O(N__1367),
            .I(N__1350));
    InMux I__154 (
            .O(N__1366),
            .I(N__1350));
    InMux I__153 (
            .O(N__1365),
            .I(N__1345));
    InMux I__152 (
            .O(N__1364),
            .I(N__1345));
    LocalMux I__151 (
            .O(N__1361),
            .I(N__1340));
    LocalMux I__150 (
            .O(N__1356),
            .I(N__1340));
    InMux I__149 (
            .O(N__1355),
            .I(N__1337));
    LocalMux I__148 (
            .O(N__1350),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__147 (
            .O(N__1345),
            .I(\uart.timer_CountZ0Z_6 ));
    Odrv4 I__146 (
            .O(N__1340),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__145 (
            .O(N__1337),
            .I(\uart.timer_CountZ0Z_6 ));
    CEMux I__144 (
            .O(N__1328),
            .I(N__1325));
    LocalMux I__143 (
            .O(N__1325),
            .I(N__1322));
    Odrv4 I__142 (
            .O(N__1322),
            .I(\uart.N_44_0 ));
    CascadeMux I__141 (
            .O(N__1319),
            .I(\uart.N_147_0_cascade_ ));
    InMux I__140 (
            .O(N__1316),
            .I(N__1313));
    LocalMux I__139 (
            .O(N__1313),
            .I(\uart.timer_Count_RNITC202Z0Z_6 ));
    CascadeMux I__138 (
            .O(N__1310),
            .I(\uart.timer_Count_RNIGLM11Z0Z_6_cascade_ ));
    InMux I__137 (
            .O(N__1307),
            .I(N__1303));
    InMux I__136 (
            .O(N__1306),
            .I(N__1300));
    LocalMux I__135 (
            .O(N__1303),
            .I(\uart.un1_state_7_0_0 ));
    LocalMux I__134 (
            .O(N__1300),
            .I(\uart.un1_state_7_0_0 ));
    CascadeMux I__133 (
            .O(N__1295),
            .I(\uart.un1_state_7_0_0_cascade_ ));
    InMux I__132 (
            .O(N__1292),
            .I(N__1286));
    InMux I__131 (
            .O(N__1291),
            .I(N__1286));
    LocalMux I__130 (
            .O(N__1286),
            .I(\uart.N_177 ));
    InMux I__129 (
            .O(N__1283),
            .I(N__1280));
    LocalMux I__128 (
            .O(N__1280),
            .I(N__1277));
    Odrv4 I__127 (
            .O(N__1277),
            .I(\uart.un1_state_5 ));
    CascadeMux I__126 (
            .O(N__1274),
            .I(\uart.state_RNO_1Z0Z_2_cascade_ ));
    InMux I__125 (
            .O(N__1271),
            .I(N__1268));
    LocalMux I__124 (
            .O(N__1268),
            .I(\uart.state_RNO_2Z0Z_2 ));
    CascadeMux I__123 (
            .O(N__1265),
            .I(\uart.N_170_cascade_ ));
    CascadeMux I__122 (
            .O(N__1262),
            .I(N__1257));
    CascadeMux I__121 (
            .O(N__1261),
            .I(N__1254));
    InMux I__120 (
            .O(N__1260),
            .I(N__1244));
    InMux I__119 (
            .O(N__1257),
            .I(N__1244));
    InMux I__118 (
            .O(N__1254),
            .I(N__1244));
    InMux I__117 (
            .O(N__1253),
            .I(N__1244));
    LocalMux I__116 (
            .O(N__1244),
            .I(\uart.stateZ0Z_2 ));
    CascadeMux I__115 (
            .O(N__1241),
            .I(N__1237));
    InMux I__114 (
            .O(N__1240),
            .I(N__1229));
    InMux I__113 (
            .O(N__1237),
            .I(N__1229));
    InMux I__112 (
            .O(N__1236),
            .I(N__1229));
    LocalMux I__111 (
            .O(N__1229),
            .I(\uart.stateZ0Z_1 ));
    CascadeMux I__110 (
            .O(N__1226),
            .I(\uart.data_Aux_esr_RNO_0Z0Z_7_cascade_ ));
    CascadeMux I__109 (
            .O(N__1223),
            .I(\uart.CO0_0_cascade_ ));
    CascadeMux I__108 (
            .O(N__1220),
            .I(\uart.bit_Count_RNO_1Z0Z_2_cascade_ ));
    CascadeMux I__107 (
            .O(N__1217),
            .I(\uart.CO1_1_cascade_ ));
    InMux I__106 (
            .O(N__1214),
            .I(N__1211));
    LocalMux I__105 (
            .O(N__1211),
            .I(\uart.bit_Count_RNO_2Z0Z_2 ));
    InMux I__104 (
            .O(N__1208),
            .I(N__1205));
    LocalMux I__103 (
            .O(N__1205),
            .I(\uart.bit_Count_RNO_1Z0Z_1 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uart.bit_Count_RNO_0_1_LC_13_17_1 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_1_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_1_LC_13_17_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uart.bit_Count_RNO_0_1_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__1208),
            .in2(_gnd_net_),
            .in3(N__2586),
            .lcout(),
            .ltout(\uart.CO0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_1_LC_13_17_2 .C_ON=1'b0;
    defparam \uart.bit_Count_1_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_1_LC_13_17_2 .LUT_INIT=16'b0101011100100000;
    LogicCell40 \uart.bit_Count_1_LC_13_17_2  (
            .in0(N__1779),
            .in1(N__1307),
            .in2(N__1223),
            .in3(N__2114),
            .lcout(\uart.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2749),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_1_2_LC_13_18_2 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_1_2_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_1_2_LC_13_18_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uart.bit_Count_RNO_1_2_LC_13_18_2  (
            .in0(N__2202),
            .in1(N__2098),
            .in2(N__1931),
            .in3(N__2573),
            .lcout(),
            .ltout(\uart.bit_Count_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_0_2_LC_13_18_3 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_2_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_2_LC_13_18_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \uart.bit_Count_RNO_0_2_LC_13_18_3  (
            .in0(N__1615),
            .in1(N__1214),
            .in2(N__1220),
            .in3(N__1517),
            .lcout(),
            .ltout(\uart.CO1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_2_LC_13_18_4 .C_ON=1'b0;
    defparam \uart.bit_Count_2_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_2_LC_13_18_4 .LUT_INIT=16'b0101011100100000;
    LogicCell40 \uart.bit_Count_2_LC_13_18_4  (
            .in0(N__1780),
            .in1(N__1306),
            .in2(N__1217),
            .in3(N__2488),
            .lcout(\uart.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2746),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_2_2_LC_13_18_6 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_2_2_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_2_2_LC_13_18_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart.bit_Count_RNO_2_2_LC_13_18_6  (
            .in0(N__2200),
            .in1(N__2097),
            .in2(_gnd_net_),
            .in3(N__2572),
            .lcout(\uart.bit_Count_RNO_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_1_1_LC_13_18_7 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_1_1_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_1_1_LC_13_18_7 .LUT_INIT=16'b0000000010110011;
    LogicCell40 \uart.bit_Count_RNO_1_1_LC_13_18_7  (
            .in0(N__1372),
            .in1(N__1900),
            .in2(N__1616),
            .in3(N__2201),
            .lcout(\uart.bit_Count_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_1_3_LC_13_19_0 .C_ON=1'b0;
    defparam \uart.state_RNO_1_3_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_1_3_LC_13_19_0 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \uart.state_RNO_1_3_LC_13_19_0  (
            .in0(N__1933),
            .in1(N__1476),
            .in2(N__1261),
            .in3(N__1606),
            .lcout(\uart.state_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIB0BC_2_LC_13_19_1 .C_ON=1'b0;
    defparam \uart.state_RNIB0BC_2_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIB0BC_2_LC_13_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart.state_RNIB0BC_2_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__1253),
            .in2(_gnd_net_),
            .in3(N__1932),
            .lcout(\uart.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_2_2_LC_13_19_2 .C_ON=1'b0;
    defparam \uart.state_RNO_2_2_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_2_2_LC_13_19_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart.state_RNO_2_2_LC_13_19_2  (
            .in0(N__1364),
            .in1(N__1236),
            .in2(_gnd_net_),
            .in3(N__1604),
            .lcout(\uart.state_RNO_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_1_2_LC_13_19_3 .C_ON=1'b0;
    defparam \uart.state_RNO_1_2_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_1_2_LC_13_19_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uart.state_RNO_1_2_LC_13_19_3  (
            .in0(N__1605),
            .in1(N__1365),
            .in2(N__1241),
            .in3(N__1853),
            .lcout(),
            .ltout(\uart.state_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_2_LC_13_19_4 .C_ON=1'b0;
    defparam \uart.state_RNO_0_2_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_2_LC_13_19_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uart.state_RNO_0_2_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__1402),
            .in2(N__1274),
            .in3(N__1271),
            .lcout(),
            .ltout(\uart.N_170_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_2_LC_13_19_5 .C_ON=1'b0;
    defparam \uart.state_2_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \uart.state_2_LC_13_19_5 .LUT_INIT=16'b0000111100000010;
    LogicCell40 \uart.state_2_LC_13_19_5  (
            .in0(N__1240),
            .in1(N__2902),
            .in2(N__1265),
            .in3(N__1260),
            .lcout(\uart.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2743),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_1_LC_13_19_6 .C_ON=1'b0;
    defparam \uart.state_1_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \uart.state_1_LC_13_19_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart.state_1_LC_13_19_6  (
            .in0(N__1934),
            .in1(N__2901),
            .in2(N__1262),
            .in3(N__2210),
            .lcout(\uart.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2743),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_3_LC_13_19_7 .C_ON=1'b0;
    defparam \uart.state_RNO_0_3_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_3_LC_13_19_7 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \uart.state_RNO_0_3_LC_13_19_7  (
            .in0(N__2033),
            .in1(N__1985),
            .in2(N__1670),
            .in3(N__1852),
            .lcout(\uart.state_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_7_LC_14_17_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_7_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_7_LC_14_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_7_LC_14_17_0  (
            .in0(N__2130),
            .in1(N__2585),
            .in2(N__2489),
            .in3(N__2437),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_7_LC_14_17_1 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_7_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_7_LC_14_17_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_7_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1226),
            .in3(N__2645),
            .lcout(\uart.N_44_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_7_LC_14_17_2 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_7_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_7_LC_14_17_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_7_LC_14_17_2  (
            .in0(N__2856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2753),
            .ce(N__1328),
            .sr(N__2646));
    defparam \uart.timer_Count_RNIBAKE2_6_LC_14_18_0 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIBAKE2_6_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIBAKE2_6_LC_14_18_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart.timer_Count_RNIBAKE2_6_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__1291),
            .in2(_gnd_net_),
            .in3(N__1316),
            .lcout(\uart.N_165_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIQ1101_3_LC_14_18_1 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIQ1101_3_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIQ1101_3_LC_14_18_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.timer_Count_RNIQ1101_3_LC_14_18_1  (
            .in0(N__2022),
            .in1(N__1978),
            .in2(_gnd_net_),
            .in3(N__1657),
            .lcout(\uart.N_147_0 ),
            .ltout(\uart.N_147_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNITC202_6_LC_14_18_2 .C_ON=1'b0;
    defparam \uart.timer_Count_RNITC202_6_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNITC202_6_LC_14_18_2 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \uart.timer_Count_RNITC202_6_LC_14_18_2  (
            .in0(N__1609),
            .in1(N__1370),
            .in2(N__1319),
            .in3(N__1846),
            .lcout(\uart.timer_Count_RNITC202Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIGLM11_6_LC_14_18_3 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIGLM11_6_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIGLM11_6_LC_14_18_3 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart.timer_Count_RNIGLM11_6_LC_14_18_3  (
            .in0(N__1371),
            .in1(N__1610),
            .in2(N__1937),
            .in3(N__2203),
            .lcout(),
            .ltout(\uart.timer_Count_RNIGLM11Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIBLJS1_3_LC_14_18_4 .C_ON=1'b0;
    defparam \uart.state_RNIBLJS1_3_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIBLJS1_3_LC_14_18_4 .LUT_INIT=16'b1111000000010001;
    LogicCell40 \uart.state_RNIBLJS1_3_LC_14_18_4  (
            .in0(N__2204),
            .in1(N__1923),
            .in2(N__1310),
            .in3(N__1292),
            .lcout(\uart.un1_state_7_0_0 ),
            .ltout(\uart.un1_state_7_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_0_LC_14_18_5 .C_ON=1'b0;
    defparam \uart.bit_Count_0_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_0_LC_14_18_5 .LUT_INIT=16'b0010011000101010;
    LogicCell40 \uart.bit_Count_0_LC_14_18_5  (
            .in0(N__2571),
            .in1(N__1781),
            .in2(N__1295),
            .in3(N__1283),
            .lcout(\uart.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2750),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNIETHE_2_LC_14_18_6 .C_ON=1'b0;
    defparam \uart.bit_Count_RNIETHE_2_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNIETHE_2_LC_14_18_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.bit_Count_RNIETHE_2_LC_14_18_6  (
            .in0(N__2096),
            .in1(N__2468),
            .in2(_gnd_net_),
            .in3(N__2570),
            .lcout(\uart.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNO_0_0_LC_14_18_7 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_0_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_0_LC_14_18_7 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart.bit_Count_RNO_0_0_LC_14_18_7  (
            .in0(N__1516),
            .in1(N__1611),
            .in2(N__1938),
            .in3(N__2205),
            .lcout(\uart.un1_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNINU001_0_1_LC_14_19_0 .C_ON=1'b0;
    defparam \uart.timer_Count_RNINU001_0_1_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNINU001_0_1_LC_14_19_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.timer_Count_RNINU001_0_1_LC_14_19_0  (
            .in0(N__2023),
            .in1(N__1979),
            .in2(_gnd_net_),
            .in3(N__1724),
            .lcout(\uart.N_22_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_3_LC_14_19_1 .C_ON=1'b0;
    defparam \uart.state_3_LC_14_19_1 .SEQ_MODE=4'b1000;
    defparam \uart.state_3_LC_14_19_1 .LUT_INIT=16'b0011111100000101;
    LogicCell40 \uart.state_3_LC_14_19_1  (
            .in0(N__1424),
            .in1(N__1441),
            .in2(N__1418),
            .in3(N__1935),
            .lcout(\uart.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2747),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_6_rep1_RNIRC5S1_LC_14_19_2 .C_ON=1'b0;
    defparam \uart.timer_Count_6_rep1_RNIRC5S1_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_6_rep1_RNIRC5S1_LC_14_19_2 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \uart.timer_Count_6_rep1_RNIRC5S1_LC_14_19_2  (
            .in0(N__1832),
            .in1(N__1508),
            .in2(N__1406),
            .in3(N__1591),
            .lcout(),
            .ltout(\uart.timer_Count_6_rep1_RNIRC5SZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNILALH5_4_LC_14_19_3 .C_ON=1'b0;
    defparam \uart.state_RNILALH5_4_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNILALH5_4_LC_14_19_3 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \uart.state_RNILALH5_4_LC_14_19_3  (
            .in0(N__1388),
            .in1(N__2236),
            .in2(N__1379),
            .in3(N__2176),
            .lcout(\uart.un1_timer_Count_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIQ9BL_0_LC_14_19_4 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIQ9BL_0_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIQ9BL_0_LC_14_19_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \uart.timer_Count_RNIQ9BL_0_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1665),
            .in3(N__1747),
            .lcout(),
            .ltout(\uart.un1_state_2_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIICSG1_6_LC_14_19_5 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIICSG1_6_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIICSG1_6_LC_14_19_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uart.timer_Count_RNIICSG1_6_LC_14_19_5  (
            .in0(N__1355),
            .in1(N__2174),
            .in2(N__1376),
            .in3(N__1830),
            .lcout(\uart.timer_Count_RNIICSG1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIN6BL_0_LC_14_19_6 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIN6BL_0_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIN6BL_0_LC_14_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart.timer_Count_RNIN6BL_0_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__1725),
            .in2(_gnd_net_),
            .in3(N__1748),
            .lcout(\uart.un4_timer_Count_1_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_fast_RNI7MEA1_6_LC_14_19_7 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_RNI7MEA1_6_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_fast_RNI7MEA1_6_LC_14_19_7 .LUT_INIT=16'b0001010111111111;
    LogicCell40 \uart.timer_Count_fast_RNI7MEA1_6_LC_14_19_7  (
            .in0(N__1590),
            .in1(N__1831),
            .in2(N__1478),
            .in3(N__2175),
            .lcout(\uart.N_28_mux_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_7_LC_14_20_0 .C_ON=1'b0;
    defparam \uart.timer_Count_7_LC_14_20_0 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_7_LC_14_20_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uart.timer_Count_7_LC_14_20_0  (
            .in0(N__1842),
            .in1(N__2051),
            .in2(N__1373),
            .in3(N__1608),
            .lcout(\uart.timer_CountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2744),
            .ce(),
            .sr(N__1692));
    defparam \uart.timer_Count_6_LC_14_20_1 .C_ON=1'b0;
    defparam \uart.timer_Count_6_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_6_LC_14_20_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uart.timer_Count_6_LC_14_20_1  (
            .in0(N__2048),
            .in1(N__1366),
            .in2(_gnd_net_),
            .in3(N__1844),
            .lcout(\uart.timer_CountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2744),
            .ce(),
            .sr(N__1692));
    defparam \uart.timer_Count_fast_6_LC_14_20_2 .C_ON=1'b0;
    defparam \uart.timer_Count_fast_6_LC_14_20_2 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_fast_6_LC_14_20_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uart.timer_Count_fast_6_LC_14_20_2  (
            .in0(N__1843),
            .in1(N__2050),
            .in2(_gnd_net_),
            .in3(N__1477),
            .lcout(\uart.timer_Count_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2744),
            .ce(),
            .sr(N__1692));
    defparam \uart.timer_Count_6_rep1_LC_14_20_3 .C_ON=1'b0;
    defparam \uart.timer_Count_6_rep1_LC_14_20_3 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_6_rep1_LC_14_20_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uart.timer_Count_6_rep1_LC_14_20_3  (
            .in0(N__2049),
            .in1(N__1515),
            .in2(_gnd_net_),
            .in3(N__1845),
            .lcout(\uart.timer_Count_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2744),
            .ce(),
            .sr(N__1692));
    defparam \uart.timer_Count_0_LC_14_20_4 .C_ON=1'b0;
    defparam \uart.timer_Count_0_LC_14_20_4 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_0_LC_14_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart.timer_Count_0_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1751),
            .lcout(\uart.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2744),
            .ce(),
            .sr(N__1692));
    defparam \uart.data_Aux_esr_1_LC_15_16_2 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_1_LC_15_16_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_1_LC_15_16_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_1_LC_15_16_2  (
            .in0(N__2890),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2758),
            .ce(N__1454),
            .sr(N__2649));
    defparam \uart.data_Aux_esr_RNO_0_4_LC_15_17_1 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_4_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_4_LC_15_17_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_4_LC_15_17_1  (
            .in0(N__2581),
            .in1(N__2517),
            .in2(N__2438),
            .in3(N__2116),
            .lcout(\uart.data_Aux_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_0_LC_15_17_2 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_0_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_0_LC_15_17_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_0_LC_15_17_2  (
            .in0(N__2115),
            .in1(N__2580),
            .in2(N__2519),
            .in3(N__2429),
            .lcout(\uart.data_Aux_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNID2BC_3_LC_15_17_5 .C_ON=1'b0;
    defparam \uart.state_RNID2BC_3_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNID2BC_3_LC_15_17_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart.state_RNID2BC_3_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__1939),
            .in2(_gnd_net_),
            .in3(N__2177),
            .lcout(\uart.un1_state_4_0_a2_iso ),
            .ltout(\uart.un1_state_4_0_a2_iso_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_1_LC_15_17_6 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_1_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_1_LC_15_17_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_1_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1457),
            .in3(N__1529),
            .lcout(\uart.N_38_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_4_LC_15_18_1 .C_ON=1'b0;
    defparam \uart.state_4_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \uart.state_4_LC_15_18_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \uart.state_4_LC_15_18_1  (
            .in0(N__2235),
            .in1(N__1442),
            .in2(N__1940),
            .in3(N__2199),
            .lcout(\uart.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2754),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNI9BTG2_6_LC_15_18_2 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI9BTG2_6_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI9BTG2_6_LC_15_18_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart.timer_Count_RNI9BTG2_6_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__2248),
            .in2(_gnd_net_),
            .in3(N__1430),
            .lcout(\uart.N_175 ),
            .ltout(\uart.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_1_LC_15_18_3 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_1_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_1_LC_15_18_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_1_LC_15_18_3  (
            .in0(N__2131),
            .in1(N__2490),
            .in2(N__1532),
            .in3(N__2574),
            .lcout(\uart.data_Aux_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_3_LC_15_18_4 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_3_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_3_LC_15_18_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_3_LC_15_18_4  (
            .in0(N__2576),
            .in1(N__2133),
            .in2(N__2509),
            .in3(N__2435),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_3_LC_15_18_5 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_3_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_3_LC_15_18_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_3_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1523),
            .in3(N__2661),
            .lcout(\uart.N_40_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_2_LC_15_18_6 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_2_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_2_LC_15_18_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_2_LC_15_18_6  (
            .in0(N__2575),
            .in1(N__2132),
            .in2(N__2508),
            .in3(N__2434),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_2_LC_15_18_7 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_2_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_2_LC_15_18_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_2_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1520),
            .in3(N__2660),
            .lcout(\uart.N_39_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_4_LC_15_19_1 .C_ON=1'b0;
    defparam \uart.timer_Count_4_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_4_LC_15_19_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uart.timer_Count_4_LC_15_19_1  (
            .in0(N__1664),
            .in1(N__2068),
            .in2(N__2031),
            .in3(N__1977),
            .lcout(\uart.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2751),
            .ce(),
            .sr(N__1703));
    defparam \uart.timer_Count_6_rep1_RNI1B4S_LC_15_19_2 .C_ON=1'b0;
    defparam \uart.timer_Count_6_rep1_RNI1B4S_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_6_rep1_RNI1B4S_LC_15_19_2 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \uart.timer_Count_6_rep1_RNI1B4S_LC_15_19_2  (
            .in0(N__1589),
            .in1(N__1506),
            .in2(_gnd_net_),
            .in3(N__1828),
            .lcout(\uart.timer_Count_6_rep1_RNI1B4SZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_6_rep1_RNI02Q61_LC_15_19_4 .C_ON=1'b0;
    defparam \uart.timer_Count_6_rep1_RNI02Q61_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_6_rep1_RNI02Q61_LC_15_19_4 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart.timer_Count_6_rep1_RNI02Q61_LC_15_19_4  (
            .in0(N__1588),
            .in1(N__1507),
            .in2(N__1666),
            .in3(N__1829),
            .lcout(\uart.timer_Count_6_rep1_RNI02QZ0Z61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNINU001_1_LC_15_19_5 .C_ON=1'b0;
    defparam \uart.timer_Count_RNINU001_1_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNINU001_1_LC_15_19_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.timer_Count_RNINU001_1_LC_15_19_5  (
            .in0(N__2017),
            .in1(N__1974),
            .in2(_gnd_net_),
            .in3(N__1723),
            .lcout(\uart.N_145_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_3_LC_15_19_6 .C_ON=1'b0;
    defparam \uart.timer_Count_3_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_3_LC_15_19_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uart.timer_Count_3_LC_15_19_6  (
            .in0(N__1976),
            .in1(_gnd_net_),
            .in2(N__2069),
            .in3(N__2018),
            .lcout(\uart.timer_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2751),
            .ce(),
            .sr(N__1703));
    defparam \uart.timer_Count_2_LC_15_19_7 .C_ON=1'b0;
    defparam \uart.timer_Count_2_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_2_LC_15_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart.timer_Count_2_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__2064),
            .in2(_gnd_net_),
            .in3(N__1975),
            .lcout(\uart.timer_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2751),
            .ce(),
            .sr(N__1703));
    defparam \uart.timer_Count_RNIMLMA1_1_LC_15_20_0 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIMLMA1_1_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIMLMA1_1_LC_15_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart.timer_Count_RNIMLMA1_1_LC_15_20_0  (
            .in0(N__1980),
            .in1(N__1660),
            .in2(N__2032),
            .in3(N__1726),
            .lcout(),
            .ltout(\uart.timer_Count_RNIMLMA1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIH8CL1_0_LC_15_20_1 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIH8CL1_0_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIH8CL1_0_LC_15_20_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uart.timer_Count_RNIH8CL1_0_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2054),
            .in3(N__1749),
            .lcout(\uart.un4_timer_Count_1_c5 ),
            .ltout(\uart.un4_timer_Count_1_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_5_LC_15_20_2 .C_ON=1'b0;
    defparam \uart.timer_Count_5_LC_15_20_2 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_5_LC_15_20_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uart.timer_Count_5_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2036),
            .in3(N__1838),
            .lcout(\uart.timer_CountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2748),
            .ce(),
            .sr(N__1702));
    defparam \uart.timer_Count_RNIHJ661_3_LC_15_20_3 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIHJ661_3_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIHJ661_3_LC_15_20_3 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \uart.timer_Count_RNIHJ661_3_LC_15_20_3  (
            .in0(N__1836),
            .in1(N__2027),
            .in2(N__1936),
            .in3(N__1981),
            .lcout(),
            .ltout(\uart.timer_Count_RNIHJ661Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNI6JN12_4_LC_15_20_4 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI6JN12_4_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI6JN12_4_LC_15_20_4 .LUT_INIT=16'b1111001111010001;
    LogicCell40 \uart.timer_Count_RNI6JN12_4_LC_15_20_4  (
            .in0(N__1927),
            .in1(N__1659),
            .in2(N__1856),
            .in3(N__1837),
            .lcout(\uart.state_0_sqmuxa_1_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_1_LC_15_20_5 .C_ON=1'b0;
    defparam \uart.timer_Count_1_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_1_LC_15_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uart.timer_Count_1_LC_15_20_5  (
            .in0(N__1727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1750),
            .lcout(\uart.timer_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2748),
            .ce(),
            .sr(N__1702));
    defparam \uart.timer_Count_RNIV5RV2_4_LC_15_20_7 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIV5RV2_4_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIV5RV2_4_LC_15_20_7 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \uart.timer_Count_RNIV5RV2_4_LC_15_20_7  (
            .in0(N__1658),
            .in1(N__1607),
            .in2(N__1547),
            .in3(N__1538),
            .lcout(\uart.state_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_rdy_LC_15_21_3 .C_ON=1'b0;
    defparam \uart.data_rdy_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_rdy_LC_15_21_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart.data_rdy_LC_15_21_3  (
            .in0(N__2866),
            .in1(N__2237),
            .in2(_gnd_net_),
            .in3(N__2209),
            .lcout(data_rdy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2745),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_LC_16_16_2 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_LC_16_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart.data_Aux_esr_RNO_0_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__2647),
            .in2(_gnd_net_),
            .in3(N__2291),
            .lcout(\uart.N_37_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_4_LC_16_16_5 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_4_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_4_LC_16_16_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart.data_Aux_esr_RNO_4_LC_16_16_5  (
            .in0(N__2648),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2285),
            .lcout(\uart.N_41_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_2_LC_16_17_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_2_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_2_LC_16_17_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_2_LC_16_17_0  (
            .in0(N__2857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2759),
            .ce(N__2279),
            .sr(N__2650));
    defparam \uart.data_Aux_esr_3_LC_16_18_2 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_3_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_3_LC_16_18_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_3_LC_16_18_2  (
            .in0(N__2906),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2756),
            .ce(N__2270),
            .sr(N__2659));
    defparam \uart.data_Aux_esr_RNO_0_6_LC_16_18_7 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_6_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_6_LC_16_18_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_6_LC_16_18_7  (
            .in0(N__2134),
            .in1(N__2587),
            .in2(N__2510),
            .in3(N__2433),
            .lcout(\uart.data_Aux_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_6_rep1_RNIOBV23_LC_16_19_0 .C_ON=1'b0;
    defparam \uart.timer_Count_6_rep1_RNIOBV23_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_6_rep1_RNIOBV23_LC_16_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart.timer_Count_6_rep1_RNIOBV23_LC_16_19_0  (
            .in0(N__2261),
            .in1(N__2255),
            .in2(_gnd_net_),
            .in3(N__2249),
            .lcout(\uart.timer_Count28 ),
            .ltout(\uart.timer_Count28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIVF8I3_4_LC_16_19_1 .C_ON=1'b0;
    defparam \uart.state_RNIVF8I3_4_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIVF8I3_4_LC_16_19_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uart.state_RNIVF8I3_4_LC_16_19_1  (
            .in0(N__2909),
            .in1(_gnd_net_),
            .in2(N__2213),
            .in3(N__2178),
            .lcout(\uart.state_RNIVF8I3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_0_5_LC_16_19_2 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_0_5_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_0_5_LC_16_19_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uart.data_Aux_esr_RNO_0_5_LC_16_19_2  (
            .in0(N__2135),
            .in1(N__2591),
            .in2(N__2518),
            .in3(N__2436),
            .lcout(),
            .ltout(\uart.data_Aux_esr_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_5_LC_16_19_3 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_5_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_5_LC_16_19_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.data_Aux_esr_RNO_5_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2399),
            .in3(N__2662),
            .lcout(\uart.N_42_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_RNO_6_LC_16_19_6 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_RNO_6_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_esr_RNO_6_LC_16_19_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart.data_Aux_esr_RNO_6_LC_16_19_6  (
            .in0(N__2663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2396),
            .lcout(\uart.N_43_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIUL3I6_4_LC_16_19_7 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIUL3I6_4_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIUL3I6_4_LC_16_19_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart.timer_Count_RNIUL3I6_4_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__2390),
            .in2(_gnd_net_),
            .in3(N__2922),
            .lcout(\uart.state_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_esr_5_LC_16_20_3 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_5_LC_16_20_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_5_LC_16_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_Aux_esr_5_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2907),
            .lcout(\uart.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2752),
            .ce(N__2384),
            .sr(N__2683));
    defparam \uart.data_Aux_esr_4_LC_17_16_5 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_4_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_4_LC_17_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_4_LC_17_16_5  (
            .in0(N__2897),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2762),
            .ce(N__2378),
            .sr(N__2676));
    defparam \uart.data_Aux_esr_0_LC_17_17_1 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_0_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_0_LC_17_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_0_LC_17_17_1  (
            .in0(N__2858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2761),
            .ce(N__2369),
            .sr(N__2675));
    defparam \uart.data_esr_0_LC_17_18_0 .C_ON=1'b0;
    defparam \uart.data_esr_0_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_0_LC_17_18_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart.data_esr_0_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__2363),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2760),
            .ce(N__2954),
            .sr(N__2936));
    defparam \uart.data_esr_1_LC_17_18_1 .C_ON=1'b0;
    defparam \uart.data_esr_1_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_1_LC_17_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_esr_1_LC_17_18_1  (
            .in0(N__2342),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2760),
            .ce(N__2954),
            .sr(N__2936));
    defparam \uart.data_esr_2_LC_17_18_2 .C_ON=1'b0;
    defparam \uart.data_esr_2_LC_17_18_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_2_LC_17_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_2_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3113),
            .lcout(data_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2760),
            .ce(N__2954),
            .sr(N__2936));
    defparam \uart.data_esr_3_LC_17_18_3 .C_ON=1'b0;
    defparam \uart.data_esr_3_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_3_LC_17_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_3_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3086),
            .lcout(data_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2760),
            .ce(N__2954),
            .sr(N__2936));
    defparam \uart.data_esr_5_LC_17_18_5 .C_ON=1'b0;
    defparam \uart.data_esr_5_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_5_LC_17_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_5_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3056),
            .lcout(data_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2760),
            .ce(N__2954),
            .sr(N__2936));
    defparam \uart.data_esr_6_LC_17_18_6 .C_ON=1'b0;
    defparam \uart.data_esr_6_LC_17_18_6 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_6_LC_17_18_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_esr_6_LC_17_18_6  (
            .in0(N__2771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2760),
            .ce(N__2954),
            .sr(N__2936));
    defparam \uart.data_esr_7_LC_17_18_7 .C_ON=1'b0;
    defparam \uart.data_esr_7_LC_17_18_7 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_7_LC_17_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_7_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3011),
            .lcout(data_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2760),
            .ce(N__2954),
            .sr(N__2936));
    defparam \uart.data_esr_4_LC_17_19_5 .C_ON=1'b0;
    defparam \uart.data_esr_4_LC_17_19_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_4_LC_17_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_4_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2981),
            .lcout(data_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2757),
            .ce(N__2953),
            .sr(N__2929));
    defparam \uart.data_Aux_esr_6_LC_17_20_0 .C_ON=1'b0;
    defparam \uart.data_Aux_esr_6_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_esr_6_LC_17_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_Aux_esr_6_LC_17_20_0  (
            .in0(N__2908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2755),
            .ce(N__2696),
            .sr(N__2684));
endmodule // Pc2Drone
