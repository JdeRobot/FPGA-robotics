-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Apr 3 2019 22:10:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2drone
entity Pc2drone is
port (
    uart_input_drone : in std_logic;
    uart_data_rdy_debug : out std_logic;
    ppm_output : out std_logic;
    uart_input_pc : in std_logic;
    uart_input_debug : out std_logic;
    drone_frame_decoder_data_rdy_debug : out std_logic;
    clk_system : in std_logic);
end Pc2drone;

-- Architecture of Pc2drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2drone is

signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10124\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_2\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_5\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_4\ : std_logic;
signal \frame_dron_decoder_1.WDT_RNIMRG3Z0Z_4\ : std_logic;
signal \frame_dron_decoder_1.WDT_RNI6TFJ1Z0Z_10_cascade_\ : std_logic;
signal \frame_dron_decoder_1.WDT10lt14_0_cascade_\ : std_logic;
signal \frame_dron_decoder_1.WDT10lt14_0\ : std_logic;
signal \frame_dron_decoder_1.WDT10lto13_1\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_7\ : std_logic;
signal \frame_dron_decoder_1.state_ns_i_a2_0_2_0_cascade_\ : std_logic;
signal \frame_dron_decoder_1.state_ns_i_a3_1_0_cascade_\ : std_logic;
signal \frame_dron_decoder_1.N_229_cascade_\ : std_logic;
signal \frame_dron_decoder_1.state_ns_i_a2_0_2_0\ : std_logic;
signal \frame_dron_decoder_1.N_231\ : std_logic;
signal \frame_dron_decoder_1.state_ns_0_a3_0_0_1_cascade_\ : std_logic;
signal \frame_dron_decoder_1.state_ns_0_a3_0_3_1\ : std_logic;
signal \frame_dron_decoder_1.N_249\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_3\ : std_logic;
signal \frame_dron_decoder_1.WDT10_0_i\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_0\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_1\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_0\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_2\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_1\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_3\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_2\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_4\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_3\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_5\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_4\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_6\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_5\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_7\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_6\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_7\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_8\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_9\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_8\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_10\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_9\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_11\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_10\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_12\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_11\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_13\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_12\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_14\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_13\ : std_logic;
signal \frame_dron_decoder_1.un1_WDT_cry_14\ : std_logic;
signal \frame_dron_decoder_1.WDTZ0Z_15\ : std_logic;
signal \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_1\ : std_logic;
signal uart_drone_data_4 : std_logic;
signal \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3_cascade_\ : std_logic;
signal \frame_dron_decoder_1.state_ns_0_a3_0_3_3\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_0\ : std_logic;
signal \frame_dron_decoder_1.state_ns_i_a2_1_2_0\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.reset6_3_cascade_\ : std_logic;
signal \reset_module_System.reset6_13\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.reset6_17_cascade_\ : std_logic;
signal \reset_module_System.reset6_11\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.reset6_15_cascade_\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \frame_dron_decoder_1.stateZ0Z_6\ : std_logic;
signal drone_frame_decoder_data_rdy_debug_c : std_logic;
signal uart_drone_data_2 : std_logic;
signal \frame_dron_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_\ : std_logic;
signal \frame_dron_decoder_1.N_255\ : std_logic;
signal uart_data_rdy_debug_c : std_logic;
signal \frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal uart_drone_data_1 : std_logic;
signal uart_drone_data_3 : std_logic;
signal uart_drone_data_0 : std_logic;
signal uart_drone_data_5 : std_logic;
signal uart_drone_data_6 : std_logic;
signal uart_drone_data_7 : std_logic;
signal \uart_drone.state_1_sqmuxa_0\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_1\ : std_logic;
signal \uart_drone.data_AuxZ0Z_3\ : std_logic;
signal \uart_drone.data_Auxce_0_0_4_cascade_\ : std_logic;
signal \uart_drone.data_AuxZ0Z_4\ : std_logic;
signal \uart_drone.data_Auxce_0_0_0\ : std_logic;
signal \uart_drone.state_1_sqmuxa\ : std_logic;
signal \uart_drone.data_Auxce_0_1\ : std_logic;
signal \uart_drone.data_Auxce_0_3\ : std_logic;
signal \uart_drone.N_126_li_cascade_\ : std_logic;
signal \uart_drone.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_3\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_2\ : std_logic;
signal \uart_drone.timer_CountZ1Z_2\ : std_logic;
signal \uart_drone.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \reset_module_System.count_1_1_cascade_\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \uart_drone_sync.aux_3__0__0_0\ : std_logic;
signal \uart_pc.stateZ0Z_1\ : std_logic;
signal \uart_pc.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_pc.state_srsts_0_0_0\ : std_logic;
signal \uart_pc.stateZ0Z_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_7\ : std_logic;
signal \uart_drone.data_AuxZ0Z_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_6\ : std_logic;
signal \uart_drone.data_Auxce_0_5\ : std_logic;
signal \uart_drone.un1_state_2_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_5\ : std_logic;
signal \uart_drone.data_Auxce_0_6\ : std_logic;
signal \uart_drone.data_Auxce_0_0_2\ : std_logic;
signal \uart_drone.state_RNIOU0NZ0Z_4\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_4\ : std_logic;
signal \uart_drone.N_143_cascade_\ : std_logic;
signal \uart_drone.timer_CountZ0Z_0\ : std_logic;
signal \uart_drone.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_1_cascade_\ : std_logic;
signal \uart_drone.timer_CountZ1Z_1\ : std_logic;
signal \uart_drone.N_143\ : std_logic;
signal \uart_drone.N_144_1\ : std_logic;
signal \uart_drone.N_144_1_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_2\ : std_logic;
signal \uart_drone.N_145\ : std_logic;
signal \uart_drone.timer_CountZ1Z_3\ : std_logic;
signal \uart_drone.stateZ0Z_3\ : std_logic;
signal \uart_drone.N_152\ : std_logic;
signal uart_input_debug_c : std_logic;
signal \uart_drone.timer_CountZ0Z_4\ : std_logic;
signal \uart_drone.N_126_li\ : std_logic;
signal \uart_drone.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_4\ : std_logic;
signal \uart_drone.stateZ0Z_0\ : std_logic;
signal \uart_drone.un1_state_4_0\ : std_logic;
signal \uart_drone.bit_CountZ0Z_0\ : std_logic;
signal \uart_drone.CO0\ : std_logic;
signal \uart_drone.un1_state_7_0\ : std_logic;
signal \uart_drone.bit_CountZ0Z_1\ : std_logic;
signal \uart_drone.bit_CountZ0Z_2\ : std_logic;
signal \uart_drone_sync.aux_2__0__0_0\ : std_logic;
signal \uart_pc.data_Auxce_0_6\ : std_logic;
signal \uart_pc.data_Auxce_0_1\ : std_logic;
signal \uart_pc.state_RNIEAGSZ0Z_4\ : std_logic;
signal \uart_pc.data_Auxce_0_0_2\ : std_logic;
signal \uart_pc.data_Auxce_0_3\ : std_logic;
signal \uart_pc.data_Auxce_0_5\ : std_logic;
signal \uart_pc.data_Auxce_0_0_4\ : std_logic;
signal \uart_pc.data_Auxce_0_0_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_2\ : std_logic;
signal \uart_pc.un1_state_4_0_cascade_\ : std_logic;
signal \uart_pc.CO0\ : std_logic;
signal \uart_pc.un1_state_7_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_1\ : std_logic;
signal \uart_pc.un1_state_4_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_0\ : std_logic;
signal \uart_pc.N_145_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_2\ : std_logic;
signal \uart_pc.N_152\ : std_logic;
signal \uart_pc.N_144_1\ : std_logic;
signal \uart_pc.stateZ0Z_3\ : std_logic;
signal \uart_pc.un1_state_2_0\ : std_logic;
signal \uart_pc.N_126_li\ : std_logic;
signal \uart_pc.stateZ0Z_4\ : std_logic;
signal \uart_pc.N_126_li_cascade_\ : std_logic;
signal \uart_pc.N_143_cascade_\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_1\ : std_logic;
signal \uart_pc.timer_CountZ1Z_1\ : std_logic;
signal \uart_pc.timer_CountZ0Z_0\ : std_logic;
signal \uart_pc.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \uart_pc.timer_CountZ0Z_4\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_2\ : std_logic;
signal \uart_pc.timer_CountZ1Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_3\ : std_logic;
signal \uart_pc.N_143\ : std_logic;
signal \uart_pc.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_pc.timer_CountZ1Z_3\ : std_logic;
signal uart_input_drone_c : std_logic;
signal \uart_drone_sync.aux_0__0__0_0\ : std_logic;
signal \uart_drone_sync.aux_1__0__0_0\ : std_logic;
signal \uart_pc.data_AuxZ0Z_1\ : std_logic;
signal \uart_pc.data_AuxZ0Z_0\ : std_logic;
signal \uart_pc.data_AuxZ0Z_4\ : std_logic;
signal \uart_pc.data_AuxZ0Z_2\ : std_logic;
signal \uart_pc.data_AuxZ0Z_3\ : std_logic;
signal \uart_pc.data_AuxZ0Z_5\ : std_logic;
signal \uart_pc.data_AuxZ0Z_7\ : std_logic;
signal \uart_frame_decoder.source_offset2data_1_sqmuxa_cascade_\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \uart_frame_decoder.source_offset1data_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_2\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\ : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_4\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_7\ : std_logic;
signal \bfn_7_27_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_11\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_15\ : std_logic;
signal \bfn_7_28_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_16\ : std_logic;
signal uart_input_pc_c : std_logic;
signal \uart_pc_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_1__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_3__0_Z0Z_0\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_RNO_3Z0Z_0_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\ : std_logic;
signal \uart_frame_decoder.N_138_4\ : std_logic;
signal \uart_frame_decoder.N_138_4_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_1\ : std_logic;
signal \uart_frame_decoder.state_1_RNO_2Z0Z_0\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_\ : std_logic;
signal \uart_frame_decoder.N_85_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_6\ : std_logic;
signal \uart_frame_decoder.source_offset1data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_7\ : std_logic;
signal \uart_frame_decoder.source_offset2data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_8\ : std_logic;
signal \uart_frame_decoder.source_offset3data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.source_offset2data_1_sqmuxa_0\ : std_logic;
signal \uart_frame_decoder.source_offset3data_1_sqmuxa_0\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_\ : std_logic;
signal \uart_frame_decoder.WDT8lto13_1\ : std_logic;
signal \uart_frame_decoder.WDT8lt14_0\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \uart_frame_decoder.WDT8lt14_0_cascade_\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \uart_frame_decoder.WDT8_0_i\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \uart_frame_decoder.WDT_RNIQAB11Z0Z_4\ : std_logic;
signal \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \frame_decoder_CH1data_1\ : std_logic;
signal \frame_decoder_OFF1data_1\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH1data_2\ : std_logic;
signal \frame_decoder_OFF1data_2\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH1data_3\ : std_logic;
signal \frame_decoder_OFF1data_3\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH1data_4\ : std_logic;
signal \frame_decoder_OFF1data_4\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH1data_5\ : std_logic;
signal \frame_decoder_OFF1data_5\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH1data_6\ : std_logic;
signal \frame_decoder_OFF1data_6\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_1.un3_source_data_0_axb_7\ : std_logic;
signal \frame_decoder_CH1data_7\ : std_logic;
signal \frame_decoder_OFF1data_7\ : std_logic;
signal \scaler_1.N_508_i_l_ofxZ0\ : std_logic;
signal \uart_frame_decoder.count_RNIHJ501Z0Z_0\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \uart_frame_decoder.count8_axb_1\ : std_logic;
signal \uart_frame_decoder.count8_cry_0\ : std_logic;
signal \uart_frame_decoder.count_i_2\ : std_logic;
signal \uart_frame_decoder.count8_cry_1\ : std_logic;
signal \uart_frame_decoder.count8\ : std_logic;
signal \uart_frame_decoder.source_CH1data_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_10\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\ : std_logic;
signal \ppm_encoder_1.N_299\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_1\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_62_d_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_0_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_2_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_4\ : std_logic;
signal \uart_pc.data_AuxZ0Z_6\ : std_logic;
signal \uart_pc.state_1_sqmuxa_0\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2\ : std_logic;
signal \uart_frame_decoder.state_1_ns_i_i_0_0\ : std_logic;
signal \uart_frame_decoder.N_39_i_1\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_0\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_9\ : std_logic;
signal \uart_frame_decoder.source_offset4data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.source_offset4data_1_sqmuxa_cascade_\ : std_logic;
signal \uart_frame_decoder.countZ0Z_2\ : std_logic;
signal \uart_frame_decoder.countZ0Z_1\ : std_logic;
signal \uart_frame_decoder.state_1_RNINMHJZ0Z_10_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_o2_0_10\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \frame_decoder_CH2data_1\ : std_logic;
signal \frame_decoder_OFF2data_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH2data_2\ : std_logic;
signal \frame_decoder_OFF2data_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH2data_3\ : std_logic;
signal \frame_decoder_OFF2data_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH2data_4\ : std_logic;
signal \frame_decoder_OFF2data_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH2data_5\ : std_logic;
signal \frame_decoder_OFF2data_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH2data_6\ : std_logic;
signal \frame_decoder_OFF2data_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_3\ : std_logic;
signal \uart_frame_decoder.source_CH2data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.source_CH2data_1_sqmuxa_cascade_\ : std_logic;
signal \scaler_2.N_520_i_l_ofxZ0\ : std_logic;
signal scaler_1_data_5 : std_logic;
signal scaler_3_data_5 : std_logic;
signal scaler_1_data_4 : std_logic;
signal \frame_decoder_OFF2data_0\ : std_logic;
signal \frame_decoder_CH2data_0\ : std_logic;
signal scaler_2_data_4 : std_logic;
signal scaler_3_data_4 : std_logic;
signal scaler_4_data_4 : std_logic;
signal \uart_frame_decoder.state_1Z0Z_10\ : std_logic;
signal \uart_frame_decoder.count8_THRU_CO\ : std_logic;
signal uart_input_pc_sync : std_logic;
signal \uart_pc.state_1_sqmuxa\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_11\ : std_logic;
signal \ppm_encoder_1.N_306_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_8\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_9\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_4\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_4\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_5\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_5\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_5\ : std_logic;
signal \ppm_encoder_1.N_300_cascade_\ : std_logic;
signal scaler_2_data_5 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_1\ : std_logic;
signal \ppm_encoder_1.throttle_RNIALN65Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_2\ : std_logic;
signal \ppm_encoder_1.throttle_RNI5V123Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_3\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI60223Z0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_4\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNI8CGI5Z0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_3\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNIDHGI5Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_7\ : std_logic;
signal \ppm_encoder_1.throttle_RNIONI96Z0Z_8\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \ppm_encoder_1.throttle_RNITSI96Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_11\ : std_logic;
signal \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_13\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_16\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_18\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_17\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_15\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_15\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_162_d\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_18\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_16\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1_c_RNO_0\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \scaler_2.un2_source_data_0\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1_c_RNILSPH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_9\ : std_logic;
signal scaler_4_data_5 : std_logic;
signal \frame_decoder_OFF3data_0\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \frame_decoder_OFF3data_1\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_OFF3data_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_OFF3data_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_OFF3data_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_OFF3data_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_OFF3data_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8\ : std_logic;
signal \uart_frame_decoder.count8_0_i\ : std_logic;
signal \frame_decoder_OFF3data_7\ : std_logic;
signal \scaler_3.N_532_i_l_ofxZ0\ : std_logic;
signal \uart_frame_decoder.state_1_RNINMHJZ0Z_10\ : std_logic;
signal \uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61\ : std_logic;
signal \uart_frame_decoder.count8_0\ : std_logic;
signal \frame_decoder_OFF1data_0\ : std_logic;
signal \frame_decoder_CH1data_0\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \scaler_1.un2_source_data_0\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_1_c_RNIISC11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_9\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_11\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_11\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_8\ : std_logic;
signal \ppm_encoder_1.N_303_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_12\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_12\ : std_logic;
signal \ppm_encoder_1.N_307\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_12\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_12\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIJII96Z0Z_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_7\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_7\ : std_logic;
signal \ppm_encoder_1.N_302\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_7\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_6\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_6\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_10\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_10\ : std_logic;
signal \ppm_encoder_1.N_305_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_10\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_13\ : std_logic;
signal \ppm_encoder_1.N_308_cascade_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_13\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_9\ : std_logic;
signal \bfn_10_27_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_4\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_7\ : std_logic;
signal \bfn_10_28_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_9\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_16\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_17\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_10\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_11\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \frame_decoder_CH4data_1\ : std_logic;
signal \frame_decoder_OFF4data_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH4data_2\ : std_logic;
signal \frame_decoder_OFF4data_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH4data_3\ : std_logic;
signal \frame_decoder_OFF4data_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH4data_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH4data_5\ : std_logic;
signal \frame_decoder_OFF4data_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH4data_6\ : std_logic;
signal \frame_decoder_OFF4data_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8\ : std_logic;
signal \uart_frame_decoder.source_CH4data_1_sqmuxa_0\ : std_logic;
signal \frame_decoder_CH4data_0\ : std_logic;
signal \frame_decoder_OFF4data_0\ : std_logic;
signal \scaler_4.N_544_i_l_ofxZ0\ : std_logic;
signal \frame_decoder_OFF2data_7\ : std_logic;
signal \scaler_2.un3_source_data_0_axb_7\ : std_logic;
signal \frame_decoder_CH2data_7\ : std_logic;
signal \uart_frame_decoder.source_CH2data_1_sqmuxa_0\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_5\ : std_logic;
signal \uart_frame_decoder.source_CH4data_1_sqmuxa\ : std_logic;
signal \frame_decoder_OFF4data_7\ : std_logic;
signal \frame_decoder_CH4data_7\ : std_logic;
signal \scaler_4.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1_c_RNO_1\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \scaler_3.un2_source_data_0\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2_c_RNIR08I\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3_c_RNIU49I\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4_c_RNI19AI\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_9\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_13\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal scaler_3_data_6 : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal scaler_3_data_7 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6\ : std_logic;
signal scaler_3_data_8 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7\ : std_logic;
signal scaler_3_data_9 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8\ : std_logic;
signal scaler_3_data_10 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9\ : std_logic;
signal scaler_3_data_11 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10\ : std_logic;
signal scaler_3_data_12 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11\ : std_logic;
signal scaler_3_data_13 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_13\ : std_logic;
signal scaler_3_data_14 : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_14\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_2_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_14\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_9\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_7\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_4\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_4\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_8\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_5\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_7\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_7\ : std_logic;
signal scaler_2_data_6 : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal scaler_2_data_7 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6\ : std_logic;
signal scaler_2_data_8 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7\ : std_logic;
signal scaler_2_data_9 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8\ : std_logic;
signal scaler_2_data_10 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9\ : std_logic;
signal scaler_2_data_11 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10\ : std_logic;
signal scaler_2_data_12 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_13\ : std_logic;
signal scaler_2_data_14 : std_logic;
signal \bfn_11_25_0_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_13\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_0\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_3\ : std_logic;
signal \ppm_encoder_1.N_614_i\ : std_logic;
signal \bfn_11_28_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_7\ : std_logic;
signal \bfn_11_29_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_15\ : std_logic;
signal \bfn_11_30_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_17\ : std_logic;
signal \ppm_encoder_1.N_228_g\ : std_logic;
signal pc_frame_decoder_dv : std_logic;
signal pc_frame_decoder_dv_0 : std_logic;
signal \frame_decoder_OFF4data_4\ : std_logic;
signal \uart_frame_decoder.source_offset4data_1_sqmuxa_0\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1_c_RNO_2\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \scaler_4.un2_source_data_0\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI\ : std_logic;
signal scaler_4_data_7 : std_logic;
signal \scaler_4.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI\ : std_logic;
signal scaler_4_data_8 : std_logic;
signal \scaler_4.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3_c_RNI15MI\ : std_logic;
signal scaler_4_data_9 : std_logic;
signal \scaler_4.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4_c_RNI49NI\ : std_logic;
signal scaler_4_data_10 : std_logic;
signal \scaler_4.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8_c_RNIS918\ : std_logic;
signal scaler_4_data_13 : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_9\ : std_logic;
signal scaler_4_data_14 : std_logic;
signal pc_frame_decoder_dv_0_g : std_logic;
signal uart_pc_data_0 : std_logic;
signal \frame_decoder_CH3data_0\ : std_logic;
signal uart_pc_data_1 : std_logic;
signal \frame_decoder_CH3data_1\ : std_logic;
signal uart_pc_data_2 : std_logic;
signal \frame_decoder_CH3data_2\ : std_logic;
signal uart_pc_data_3 : std_logic;
signal \frame_decoder_CH3data_3\ : std_logic;
signal uart_pc_data_4 : std_logic;
signal \frame_decoder_CH3data_4\ : std_logic;
signal uart_pc_data_6 : std_logic;
signal \frame_decoder_CH3data_6\ : std_logic;
signal uart_pc_data_7 : std_logic;
signal \frame_decoder_CH3data_7\ : std_logic;
signal \uart_frame_decoder.source_CH1data_1_sqmuxa\ : std_logic;
signal scaler_1_data_6 : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal scaler_1_data_7 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9\ : std_logic;
signal scaler_1_data_11 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10\ : std_logic;
signal scaler_1_data_12 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11\ : std_logic;
signal scaler_1_data_13 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_13\ : std_logic;
signal scaler_1_data_14 : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_14\ : std_logic;
signal \ppm_encoder_1.scaler_1_dv_0\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\ : std_logic;
signal scaler_1_data_8 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_8\ : std_logic;
signal scaler_4_data_11 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\ : std_logic;
signal scaler_1_data_10 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_10\ : std_logic;
signal scaler_4_data_12 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.N_143_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_1\ : std_logic;
signal ppm_output_c : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\ : std_logic;
signal scaler_1_data_9 : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_7_cascade_\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_14\ : std_logic;
signal \ppm_encoder_1.N_309\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_14\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_5\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_10\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12\ : std_logic;
signal \ppm_encoder_1.N_301\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_6\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_11\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_11\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_12\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_323_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_13\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\ : std_logic;
signal \ppm_encoder_1.N_322\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_6\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_62_d\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_7\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_6\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_5\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_4\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_17\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_16\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_15\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_14\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_13\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_8\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_148_17_cascade_\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\ : std_logic;
signal \ppm_encoder_1.N_148_17\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\ : std_logic;
signal \ppm_encoder_1.N_148\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_10\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_9\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_11\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\ : std_logic;
signal \ppm_encoder_1.N_241\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2_THRU_CO\ : std_logic;
signal reset_system : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_2\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\ : std_logic;
signal \uart_frame_decoder.N_85\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_2\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_4\ : std_logic;
signal uart_pc_data_rdy : std_logic;
signal \uart_frame_decoder.source_CH3data_1_sqmuxa\ : std_logic;
signal uart_pc_data_5 : std_logic;
signal \frame_decoder_CH3data_5\ : std_logic;
signal \uart_frame_decoder.source_CH3data_1_sqmuxa_0\ : std_logic;
signal scaler_4_data_6 : std_logic;
signal \ppm_encoder_1.rudderZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_14\ : std_logic;
signal \ppm_encoder_1.N_614_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\ : std_logic;
signal \ppm_encoder_1.N_230\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_11_mux\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_9\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_304\ : std_logic;
signal scaler_2_data_13 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\ : std_logic;
signal scaler_1_dv : std_logic;
signal \ppm_encoder_1.aileronZ0Z_13\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_system_c_g : std_logic;
signal reset_system_g : std_logic;

signal clk_system_wire : std_logic;
signal uart_input_drone_wire : std_logic;
signal uart_input_pc_wire : std_logic;
signal ppm_output_wire : std_logic;
signal drone_frame_decoder_data_rdy_debug_wire : std_logic;
signal uart_input_debug_wire : std_logic;
signal uart_data_rdy_debug_wire : std_logic;

begin
    clk_system_wire <= clk_system;
    uart_input_drone_wire <= uart_input_drone;
    uart_input_pc_wire <= uart_input_pc;
    ppm_output <= ppm_output_wire;
    drone_frame_decoder_data_rdy_debug <= drone_frame_decoder_data_rdy_debug_wire;
    uart_input_debug <= uart_input_debug_wire;
    uart_data_rdy_debug <= uart_data_rdy_debug_wire;

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__26454\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26456\,
            DIN => \N__26455\,
            DOUT => \N__26454\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__26456\,
            PADOUT => \N__26455\,
            PADIN => \N__26454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_drone_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26445\,
            DIN => \N__26444\,
            DOUT => \N__26443\,
            PACKAGEPIN => uart_input_drone_wire
        );

    \uart_input_drone_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__26445\,
            PADOUT => \N__26444\,
            PADIN => \N__26443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_drone_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_pc_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26436\,
            DIN => \N__26435\,
            DOUT => \N__26434\,
            PACKAGEPIN => uart_input_pc_wire
        );

    \uart_input_pc_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__26436\,
            PADOUT => \N__26435\,
            PADIN => \N__26434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_pc_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ppm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26427\,
            DIN => \N__26426\,
            DOUT => \N__26425\,
            PACKAGEPIN => ppm_output_wire
        );

    \ppm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26427\,
            PADOUT => \N__26426\,
            PADIN => \N__26425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21440\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \drone_frame_decoder_data_rdy_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26418\,
            DIN => \N__26417\,
            DOUT => \N__26416\,
            PACKAGEPIN => drone_frame_decoder_data_rdy_debug_wire
        );

    \drone_frame_decoder_data_rdy_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26418\,
            PADOUT => \N__26417\,
            PADIN => \N__26416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26409\,
            DIN => \N__26408\,
            DOUT => \N__26407\,
            PACKAGEPIN => uart_input_debug_wire
        );

    \uart_input_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26409\,
            PADOUT => \N__26408\,
            PADIN => \N__26407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12055\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_data_rdy_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26400\,
            DIN => \N__26399\,
            DOUT => \N__26398\,
            PACKAGEPIN => uart_data_rdy_debug_wire
        );

    \uart_data_rdy_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26400\,
            PADOUT => \N__26399\,
            PADIN => \N__26398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__6282\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26378\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__6280\ : Span4Mux_h
    port map (
            O => \N__26375\,
            I => \N__26371\
        );

    \I__6279\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26368\
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__26371\,
            I => \uart_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__26368\,
            I => \uart_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__6276\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26356\
        );

    \I__6275\ : InMux
    port map (
            O => \N__26362\,
            I => \N__26352\
        );

    \I__6274\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26349\
        );

    \I__6273\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26346\
        );

    \I__6272\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26343\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__26356\,
            I => \N__26339\
        );

    \I__6270\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26336\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__26352\,
            I => \N__26333\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__26349\,
            I => \N__26325\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26325\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__26343\,
            I => \N__26325\
        );

    \I__6265\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26322\
        );

    \I__6264\ : Span4Mux_v
    port map (
            O => \N__26339\,
            I => \N__26317\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__26336\,
            I => \N__26317\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__26333\,
            I => \N__26314\
        );

    \I__6261\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26311\
        );

    \I__6260\ : Span4Mux_v
    port map (
            O => \N__26325\,
            I => \N__26304\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__26322\,
            I => \N__26304\
        );

    \I__6258\ : Span4Mux_h
    port map (
            O => \N__26317\,
            I => \N__26301\
        );

    \I__6257\ : Sp12to4
    port map (
            O => \N__26314\,
            I => \N__26296\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__26311\,
            I => \N__26296\
        );

    \I__6255\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26293\
        );

    \I__6254\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26290\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__26304\,
            I => uart_pc_data_5
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__26301\,
            I => uart_pc_data_5
        );

    \I__6251\ : Odrv12
    port map (
            O => \N__26296\,
            I => uart_pc_data_5
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__26293\,
            I => uart_pc_data_5
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__26290\,
            I => uart_pc_data_5
        );

    \I__6248\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__26273\,
            I => \frame_decoder_CH3data_5\
        );

    \I__6245\ : CEMux
    port map (
            O => \N__26270\,
            I => \N__26266\
        );

    \I__6244\ : CEMux
    port map (
            O => \N__26269\,
            I => \N__26263\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__26266\,
            I => \uart_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__26263\,
            I => \uart_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6241\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26254\
        );

    \I__6240\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26251\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26248\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__26251\,
            I => \N__26245\
        );

    \I__6237\ : Span4Mux_v
    port map (
            O => \N__26248\,
            I => \N__26242\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__26245\,
            I => \N__26239\
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__26242\,
            I => scaler_4_data_6
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__26239\,
            I => scaler_4_data_6
        );

    \I__6233\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26230\
        );

    \I__6232\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26227\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26223\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__26227\,
            I => \N__26220\
        );

    \I__6229\ : InMux
    port map (
            O => \N__26226\,
            I => \N__26217\
        );

    \I__6228\ : Span4Mux_v
    port map (
            O => \N__26223\,
            I => \N__26214\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__26220\,
            I => \N__26211\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__26217\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__26214\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__6224\ : Odrv4
    port map (
            O => \N__26211\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__6223\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26201\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__26201\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\
        );

    \I__6221\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26195\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__26195\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\
        );

    \I__6219\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26189\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__26189\,
            I => \N__26186\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__26186\,
            I => \N__26183\
        );

    \I__6216\ : Span4Mux_v
    port map (
            O => \N__26183\,
            I => \N__26180\
        );

    \I__6215\ : Odrv4
    port map (
            O => \N__26180\,
            I => \ppm_encoder_1.pulses2countZ0Z_14\
        );

    \I__6214\ : CEMux
    port map (
            O => \N__26177\,
            I => \N__26172\
        );

    \I__6213\ : CEMux
    port map (
            O => \N__26176\,
            I => \N__26168\
        );

    \I__6212\ : CEMux
    port map (
            O => \N__26175\,
            I => \N__26164\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26161\
        );

    \I__6210\ : CEMux
    port map (
            O => \N__26171\,
            I => \N__26157\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__26168\,
            I => \N__26154\
        );

    \I__6208\ : CEMux
    port map (
            O => \N__26167\,
            I => \N__26151\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__26164\,
            I => \N__26148\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__26161\,
            I => \N__26145\
        );

    \I__6205\ : CEMux
    port map (
            O => \N__26160\,
            I => \N__26142\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26139\
        );

    \I__6203\ : Span4Mux_h
    port map (
            O => \N__26154\,
            I => \N__26136\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__26151\,
            I => \N__26133\
        );

    \I__6201\ : Span4Mux_v
    port map (
            O => \N__26148\,
            I => \N__26130\
        );

    \I__6200\ : Span4Mux_s1_v
    port map (
            O => \N__26145\,
            I => \N__26127\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__26142\,
            I => \N__26124\
        );

    \I__6198\ : Span4Mux_h
    port map (
            O => \N__26139\,
            I => \N__26121\
        );

    \I__6197\ : Span4Mux_h
    port map (
            O => \N__26136\,
            I => \N__26118\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__26133\,
            I => \N__26111\
        );

    \I__6195\ : Span4Mux_v
    port map (
            O => \N__26130\,
            I => \N__26111\
        );

    \I__6194\ : Span4Mux_v
    port map (
            O => \N__26127\,
            I => \N__26111\
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__26124\,
            I => \ppm_encoder_1.N_614_0\
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__26121\,
            I => \ppm_encoder_1.N_614_0\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__26118\,
            I => \ppm_encoder_1.N_614_0\
        );

    \I__6190\ : Odrv4
    port map (
            O => \N__26111\,
            I => \ppm_encoder_1.N_614_0\
        );

    \I__6189\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26096\
        );

    \I__6188\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26093\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__26100\,
            I => \N__26087\
        );

    \I__6186\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26084\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__26096\,
            I => \N__26079\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26079\
        );

    \I__6183\ : InMux
    port map (
            O => \N__26092\,
            I => \N__26074\
        );

    \I__6182\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26074\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__26090\,
            I => \N__26068\
        );

    \I__6180\ : InMux
    port map (
            O => \N__26087\,
            I => \N__26059\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__26084\,
            I => \N__26052\
        );

    \I__6178\ : Span4Mux_h
    port map (
            O => \N__26079\,
            I => \N__26052\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__26074\,
            I => \N__26052\
        );

    \I__6176\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26049\
        );

    \I__6175\ : InMux
    port map (
            O => \N__26072\,
            I => \N__26043\
        );

    \I__6174\ : InMux
    port map (
            O => \N__26071\,
            I => \N__26043\
        );

    \I__6173\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26040\
        );

    \I__6172\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26035\
        );

    \I__6171\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26035\
        );

    \I__6170\ : CascadeMux
    port map (
            O => \N__26065\,
            I => \N__26032\
        );

    \I__6169\ : InMux
    port map (
            O => \N__26064\,
            I => \N__26028\
        );

    \I__6168\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26025\
        );

    \I__6167\ : InMux
    port map (
            O => \N__26062\,
            I => \N__26022\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__26059\,
            I => \N__26015\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__26052\,
            I => \N__26015\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__26049\,
            I => \N__26015\
        );

    \I__6163\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26012\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__26043\,
            I => \N__26008\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__26040\,
            I => \N__26005\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__26035\,
            I => \N__26002\
        );

    \I__6159\ : InMux
    port map (
            O => \N__26032\,
            I => \N__25997\
        );

    \I__6158\ : InMux
    port map (
            O => \N__26031\,
            I => \N__25997\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__26028\,
            I => \N__25994\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__26025\,
            I => \N__25991\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__26022\,
            I => \N__25988\
        );

    \I__6154\ : Span4Mux_v
    port map (
            O => \N__26015\,
            I => \N__25983\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__25983\
        );

    \I__6152\ : InMux
    port map (
            O => \N__26011\,
            I => \N__25980\
        );

    \I__6151\ : Span12Mux_v
    port map (
            O => \N__26008\,
            I => \N__25975\
        );

    \I__6150\ : Span4Mux_h
    port map (
            O => \N__26005\,
            I => \N__25968\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__26002\,
            I => \N__25968\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25968\
        );

    \I__6147\ : Span4Mux_v
    port map (
            O => \N__25994\,
            I => \N__25957\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__25991\,
            I => \N__25957\
        );

    \I__6145\ : Span4Mux_v
    port map (
            O => \N__25988\,
            I => \N__25957\
        );

    \I__6144\ : Span4Mux_v
    port map (
            O => \N__25983\,
            I => \N__25957\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__25980\,
            I => \N__25957\
        );

    \I__6142\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25952\
        );

    \I__6141\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25952\
        );

    \I__6140\ : Odrv12
    port map (
            O => \N__25975\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6139\ : Odrv4
    port map (
            O => \N__25968\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6138\ : Odrv4
    port map (
            O => \N__25957\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__25952\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6136\ : InMux
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__25940\,
            I => \N__25937\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__25937\,
            I => \N__25933\
        );

    \I__6133\ : CascadeMux
    port map (
            O => \N__25936\,
            I => \N__25926\
        );

    \I__6132\ : Span4Mux_v
    port map (
            O => \N__25933\,
            I => \N__25923\
        );

    \I__6131\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25920\
        );

    \I__6130\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25917\
        );

    \I__6129\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25914\
        );

    \I__6128\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25909\
        );

    \I__6127\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25909\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__25923\,
            I => \ppm_encoder_1.N_230\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__25920\,
            I => \ppm_encoder_1.N_230\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__25917\,
            I => \ppm_encoder_1.N_230\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__25914\,
            I => \ppm_encoder_1.N_230\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__25909\,
            I => \ppm_encoder_1.N_230\
        );

    \I__6121\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25886\
        );

    \I__6120\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25886\
        );

    \I__6119\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25880\
        );

    \I__6118\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25873\
        );

    \I__6117\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25873\
        );

    \I__6116\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25873\
        );

    \I__6115\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25870\
        );

    \I__6114\ : InMux
    port map (
            O => \N__25891\,
            I => \N__25867\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__25886\,
            I => \N__25864\
        );

    \I__6112\ : InMux
    port map (
            O => \N__25885\,
            I => \N__25854\
        );

    \I__6111\ : InMux
    port map (
            O => \N__25884\,
            I => \N__25854\
        );

    \I__6110\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25854\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__25880\,
            I => \N__25851\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__25873\,
            I => \N__25848\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__25870\,
            I => \N__25843\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__25867\,
            I => \N__25843\
        );

    \I__6105\ : Span4Mux_v
    port map (
            O => \N__25864\,
            I => \N__25840\
        );

    \I__6104\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25835\
        );

    \I__6103\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25835\
        );

    \I__6102\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25832\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__25854\,
            I => \N__25829\
        );

    \I__6100\ : Span4Mux_v
    port map (
            O => \N__25851\,
            I => \N__25824\
        );

    \I__6099\ : Span4Mux_h
    port map (
            O => \N__25848\,
            I => \N__25824\
        );

    \I__6098\ : Span4Mux_h
    port map (
            O => \N__25843\,
            I => \N__25819\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__25840\,
            I => \N__25819\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__25835\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__25832\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__25829\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__25824\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__6092\ : Odrv4
    port map (
            O => \N__25819\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__6091\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25801\
        );

    \I__6090\ : CascadeMux
    port map (
            O => \N__25807\,
            I => \N__25797\
        );

    \I__6089\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25791\
        );

    \I__6088\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25788\
        );

    \I__6087\ : CascadeMux
    port map (
            O => \N__25804\,
            I => \N__25782\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__25801\,
            I => \N__25778\
        );

    \I__6085\ : InMux
    port map (
            O => \N__25800\,
            I => \N__25774\
        );

    \I__6084\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25771\
        );

    \I__6083\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25768\
        );

    \I__6082\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25765\
        );

    \I__6081\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25762\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__25791\,
            I => \N__25757\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__25788\,
            I => \N__25757\
        );

    \I__6078\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25754\
        );

    \I__6077\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25751\
        );

    \I__6076\ : InMux
    port map (
            O => \N__25785\,
            I => \N__25748\
        );

    \I__6075\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25742\
        );

    \I__6074\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25742\
        );

    \I__6073\ : Span4Mux_v
    port map (
            O => \N__25778\,
            I => \N__25739\
        );

    \I__6072\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25736\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__25774\,
            I => \N__25727\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__25771\,
            I => \N__25727\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25724\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__25765\,
            I => \N__25721\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__25762\,
            I => \N__25714\
        );

    \I__6066\ : Span4Mux_v
    port map (
            O => \N__25757\,
            I => \N__25714\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__25754\,
            I => \N__25714\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__25751\,
            I => \N__25709\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__25748\,
            I => \N__25709\
        );

    \I__6062\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25706\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__25742\,
            I => \N__25703\
        );

    \I__6060\ : Span4Mux_v
    port map (
            O => \N__25739\,
            I => \N__25698\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25698\
        );

    \I__6058\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25695\
        );

    \I__6057\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25692\
        );

    \I__6056\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25687\
        );

    \I__6055\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25687\
        );

    \I__6054\ : Span4Mux_h
    port map (
            O => \N__25727\,
            I => \N__25674\
        );

    \I__6053\ : Span4Mux_v
    port map (
            O => \N__25724\,
            I => \N__25674\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__25721\,
            I => \N__25674\
        );

    \I__6051\ : Span4Mux_v
    port map (
            O => \N__25714\,
            I => \N__25674\
        );

    \I__6050\ : Span4Mux_v
    port map (
            O => \N__25709\,
            I => \N__25674\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__25706\,
            I => \N__25674\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__25703\,
            I => \N__25669\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__25698\,
            I => \N__25669\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__25695\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__25692\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__25687\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__25674\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6042\ : Odrv4
    port map (
            O => \N__25669\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6041\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25653\
        );

    \I__6040\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25650\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__25656\,
            I => \N__25647\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__25653\,
            I => \N__25642\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__25650\,
            I => \N__25642\
        );

    \I__6036\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25639\
        );

    \I__6035\ : Odrv12
    port map (
            O => \N__25642\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__25639\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__6033\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25629\
        );

    \I__6032\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25626\
        );

    \I__6031\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25623\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__25629\,
            I => \N__25620\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__25626\,
            I => \N__25617\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__25623\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__25620\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__25617\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__6025\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25607\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__25607\,
            I => \N__25604\
        );

    \I__6023\ : Span4Mux_h
    port map (
            O => \N__25604\,
            I => \N__25601\
        );

    \I__6022\ : Odrv4
    port map (
            O => \N__25601\,
            I => \ppm_encoder_1.N_304\
        );

    \I__6021\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25595\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__25595\,
            I => \N__25592\
        );

    \I__6019\ : Span4Mux_v
    port map (
            O => \N__25592\,
            I => \N__25588\
        );

    \I__6018\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25585\
        );

    \I__6017\ : Span4Mux_h
    port map (
            O => \N__25588\,
            I => \N__25580\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__25585\,
            I => \N__25580\
        );

    \I__6015\ : Span4Mux_v
    port map (
            O => \N__25580\,
            I => \N__25577\
        );

    \I__6014\ : Span4Mux_v
    port map (
            O => \N__25577\,
            I => \N__25574\
        );

    \I__6013\ : Odrv4
    port map (
            O => \N__25574\,
            I => scaler_2_data_13
        );

    \I__6012\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__25562\,
            I => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__25559\,
            I => \N__25555\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__25558\,
            I => \N__25551\
        );

    \I__6006\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25537\
        );

    \I__6005\ : InMux
    port map (
            O => \N__25554\,
            I => \N__25537\
        );

    \I__6004\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25534\
        );

    \I__6003\ : CascadeMux
    port map (
            O => \N__25550\,
            I => \N__25530\
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__25549\,
            I => \N__25525\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__25548\,
            I => \N__25517\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__25547\,
            I => \N__25513\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__25546\,
            I => \N__25509\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__25545\,
            I => \N__25506\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__25544\,
            I => \N__25502\
        );

    \I__5996\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25497\
        );

    \I__5995\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25497\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__25537\,
            I => \N__25491\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__25534\,
            I => \N__25488\
        );

    \I__5992\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25485\
        );

    \I__5991\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25482\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__25529\,
            I => \N__25478\
        );

    \I__5989\ : CascadeMux
    port map (
            O => \N__25528\,
            I => \N__25474\
        );

    \I__5988\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25468\
        );

    \I__5987\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25468\
        );

    \I__5986\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25461\
        );

    \I__5985\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25461\
        );

    \I__5984\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25461\
        );

    \I__5983\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25454\
        );

    \I__5982\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25454\
        );

    \I__5981\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25454\
        );

    \I__5980\ : InMux
    port map (
            O => \N__25513\,
            I => \N__25451\
        );

    \I__5979\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25448\
        );

    \I__5978\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25443\
        );

    \I__5977\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25443\
        );

    \I__5976\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25438\
        );

    \I__5975\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25438\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__25497\,
            I => \N__25435\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__25496\,
            I => \N__25431\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__25495\,
            I => \N__25426\
        );

    \I__5971\ : CascadeMux
    port map (
            O => \N__25494\,
            I => \N__25421\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__25491\,
            I => \N__25418\
        );

    \I__5969\ : Span4Mux_v
    port map (
            O => \N__25488\,
            I => \N__25411\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__25485\,
            I => \N__25411\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__25482\,
            I => \N__25411\
        );

    \I__5966\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25404\
        );

    \I__5965\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25404\
        );

    \I__5964\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25404\
        );

    \I__5963\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25401\
        );

    \I__5962\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25398\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__25468\,
            I => \N__25391\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__25461\,
            I => \N__25391\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__25454\,
            I => \N__25391\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25386\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__25448\,
            I => \N__25386\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25381\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__25438\,
            I => \N__25381\
        );

    \I__5954\ : Span4Mux_v
    port map (
            O => \N__25435\,
            I => \N__25378\
        );

    \I__5953\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25362\
        );

    \I__5952\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25362\
        );

    \I__5951\ : InMux
    port map (
            O => \N__25430\,
            I => \N__25362\
        );

    \I__5950\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25362\
        );

    \I__5949\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25362\
        );

    \I__5948\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25362\
        );

    \I__5947\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25362\
        );

    \I__5946\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25359\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__25418\,
            I => \N__25346\
        );

    \I__5944\ : Span4Mux_h
    port map (
            O => \N__25411\,
            I => \N__25346\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__25404\,
            I => \N__25346\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__25401\,
            I => \N__25346\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__25398\,
            I => \N__25346\
        );

    \I__5940\ : Span4Mux_v
    port map (
            O => \N__25391\,
            I => \N__25346\
        );

    \I__5939\ : Span4Mux_h
    port map (
            O => \N__25386\,
            I => \N__25343\
        );

    \I__5938\ : Span4Mux_v
    port map (
            O => \N__25381\,
            I => \N__25338\
        );

    \I__5937\ : Span4Mux_v
    port map (
            O => \N__25378\,
            I => \N__25338\
        );

    \I__5936\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25335\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__25362\,
            I => scaler_1_dv
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__25359\,
            I => scaler_1_dv
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__25346\,
            I => scaler_1_dv
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__25343\,
            I => scaler_1_dv
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__25338\,
            I => scaler_1_dv
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__25335\,
            I => scaler_1_dv
        );

    \I__5929\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25315\
        );

    \I__5928\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25315\
        );

    \I__5927\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25312\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__25315\,
            I => \N__25309\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__25312\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__5924\ : Odrv12
    port map (
            O => \N__25309\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__5923\ : ClkMux
    port map (
            O => \N__25304\,
            I => \N__24938\
        );

    \I__5922\ : ClkMux
    port map (
            O => \N__25303\,
            I => \N__24938\
        );

    \I__5921\ : ClkMux
    port map (
            O => \N__25302\,
            I => \N__24938\
        );

    \I__5920\ : ClkMux
    port map (
            O => \N__25301\,
            I => \N__24938\
        );

    \I__5919\ : ClkMux
    port map (
            O => \N__25300\,
            I => \N__24938\
        );

    \I__5918\ : ClkMux
    port map (
            O => \N__25299\,
            I => \N__24938\
        );

    \I__5917\ : ClkMux
    port map (
            O => \N__25298\,
            I => \N__24938\
        );

    \I__5916\ : ClkMux
    port map (
            O => \N__25297\,
            I => \N__24938\
        );

    \I__5915\ : ClkMux
    port map (
            O => \N__25296\,
            I => \N__24938\
        );

    \I__5914\ : ClkMux
    port map (
            O => \N__25295\,
            I => \N__24938\
        );

    \I__5913\ : ClkMux
    port map (
            O => \N__25294\,
            I => \N__24938\
        );

    \I__5912\ : ClkMux
    port map (
            O => \N__25293\,
            I => \N__24938\
        );

    \I__5911\ : ClkMux
    port map (
            O => \N__25292\,
            I => \N__24938\
        );

    \I__5910\ : ClkMux
    port map (
            O => \N__25291\,
            I => \N__24938\
        );

    \I__5909\ : ClkMux
    port map (
            O => \N__25290\,
            I => \N__24938\
        );

    \I__5908\ : ClkMux
    port map (
            O => \N__25289\,
            I => \N__24938\
        );

    \I__5907\ : ClkMux
    port map (
            O => \N__25288\,
            I => \N__24938\
        );

    \I__5906\ : ClkMux
    port map (
            O => \N__25287\,
            I => \N__24938\
        );

    \I__5905\ : ClkMux
    port map (
            O => \N__25286\,
            I => \N__24938\
        );

    \I__5904\ : ClkMux
    port map (
            O => \N__25285\,
            I => \N__24938\
        );

    \I__5903\ : ClkMux
    port map (
            O => \N__25284\,
            I => \N__24938\
        );

    \I__5902\ : ClkMux
    port map (
            O => \N__25283\,
            I => \N__24938\
        );

    \I__5901\ : ClkMux
    port map (
            O => \N__25282\,
            I => \N__24938\
        );

    \I__5900\ : ClkMux
    port map (
            O => \N__25281\,
            I => \N__24938\
        );

    \I__5899\ : ClkMux
    port map (
            O => \N__25280\,
            I => \N__24938\
        );

    \I__5898\ : ClkMux
    port map (
            O => \N__25279\,
            I => \N__24938\
        );

    \I__5897\ : ClkMux
    port map (
            O => \N__25278\,
            I => \N__24938\
        );

    \I__5896\ : ClkMux
    port map (
            O => \N__25277\,
            I => \N__24938\
        );

    \I__5895\ : ClkMux
    port map (
            O => \N__25276\,
            I => \N__24938\
        );

    \I__5894\ : ClkMux
    port map (
            O => \N__25275\,
            I => \N__24938\
        );

    \I__5893\ : ClkMux
    port map (
            O => \N__25274\,
            I => \N__24938\
        );

    \I__5892\ : ClkMux
    port map (
            O => \N__25273\,
            I => \N__24938\
        );

    \I__5891\ : ClkMux
    port map (
            O => \N__25272\,
            I => \N__24938\
        );

    \I__5890\ : ClkMux
    port map (
            O => \N__25271\,
            I => \N__24938\
        );

    \I__5889\ : ClkMux
    port map (
            O => \N__25270\,
            I => \N__24938\
        );

    \I__5888\ : ClkMux
    port map (
            O => \N__25269\,
            I => \N__24938\
        );

    \I__5887\ : ClkMux
    port map (
            O => \N__25268\,
            I => \N__24938\
        );

    \I__5886\ : ClkMux
    port map (
            O => \N__25267\,
            I => \N__24938\
        );

    \I__5885\ : ClkMux
    port map (
            O => \N__25266\,
            I => \N__24938\
        );

    \I__5884\ : ClkMux
    port map (
            O => \N__25265\,
            I => \N__24938\
        );

    \I__5883\ : ClkMux
    port map (
            O => \N__25264\,
            I => \N__24938\
        );

    \I__5882\ : ClkMux
    port map (
            O => \N__25263\,
            I => \N__24938\
        );

    \I__5881\ : ClkMux
    port map (
            O => \N__25262\,
            I => \N__24938\
        );

    \I__5880\ : ClkMux
    port map (
            O => \N__25261\,
            I => \N__24938\
        );

    \I__5879\ : ClkMux
    port map (
            O => \N__25260\,
            I => \N__24938\
        );

    \I__5878\ : ClkMux
    port map (
            O => \N__25259\,
            I => \N__24938\
        );

    \I__5877\ : ClkMux
    port map (
            O => \N__25258\,
            I => \N__24938\
        );

    \I__5876\ : ClkMux
    port map (
            O => \N__25257\,
            I => \N__24938\
        );

    \I__5875\ : ClkMux
    port map (
            O => \N__25256\,
            I => \N__24938\
        );

    \I__5874\ : ClkMux
    port map (
            O => \N__25255\,
            I => \N__24938\
        );

    \I__5873\ : ClkMux
    port map (
            O => \N__25254\,
            I => \N__24938\
        );

    \I__5872\ : ClkMux
    port map (
            O => \N__25253\,
            I => \N__24938\
        );

    \I__5871\ : ClkMux
    port map (
            O => \N__25252\,
            I => \N__24938\
        );

    \I__5870\ : ClkMux
    port map (
            O => \N__25251\,
            I => \N__24938\
        );

    \I__5869\ : ClkMux
    port map (
            O => \N__25250\,
            I => \N__24938\
        );

    \I__5868\ : ClkMux
    port map (
            O => \N__25249\,
            I => \N__24938\
        );

    \I__5867\ : ClkMux
    port map (
            O => \N__25248\,
            I => \N__24938\
        );

    \I__5866\ : ClkMux
    port map (
            O => \N__25247\,
            I => \N__24938\
        );

    \I__5865\ : ClkMux
    port map (
            O => \N__25246\,
            I => \N__24938\
        );

    \I__5864\ : ClkMux
    port map (
            O => \N__25245\,
            I => \N__24938\
        );

    \I__5863\ : ClkMux
    port map (
            O => \N__25244\,
            I => \N__24938\
        );

    \I__5862\ : ClkMux
    port map (
            O => \N__25243\,
            I => \N__24938\
        );

    \I__5861\ : ClkMux
    port map (
            O => \N__25242\,
            I => \N__24938\
        );

    \I__5860\ : ClkMux
    port map (
            O => \N__25241\,
            I => \N__24938\
        );

    \I__5859\ : ClkMux
    port map (
            O => \N__25240\,
            I => \N__24938\
        );

    \I__5858\ : ClkMux
    port map (
            O => \N__25239\,
            I => \N__24938\
        );

    \I__5857\ : ClkMux
    port map (
            O => \N__25238\,
            I => \N__24938\
        );

    \I__5856\ : ClkMux
    port map (
            O => \N__25237\,
            I => \N__24938\
        );

    \I__5855\ : ClkMux
    port map (
            O => \N__25236\,
            I => \N__24938\
        );

    \I__5854\ : ClkMux
    port map (
            O => \N__25235\,
            I => \N__24938\
        );

    \I__5853\ : ClkMux
    port map (
            O => \N__25234\,
            I => \N__24938\
        );

    \I__5852\ : ClkMux
    port map (
            O => \N__25233\,
            I => \N__24938\
        );

    \I__5851\ : ClkMux
    port map (
            O => \N__25232\,
            I => \N__24938\
        );

    \I__5850\ : ClkMux
    port map (
            O => \N__25231\,
            I => \N__24938\
        );

    \I__5849\ : ClkMux
    port map (
            O => \N__25230\,
            I => \N__24938\
        );

    \I__5848\ : ClkMux
    port map (
            O => \N__25229\,
            I => \N__24938\
        );

    \I__5847\ : ClkMux
    port map (
            O => \N__25228\,
            I => \N__24938\
        );

    \I__5846\ : ClkMux
    port map (
            O => \N__25227\,
            I => \N__24938\
        );

    \I__5845\ : ClkMux
    port map (
            O => \N__25226\,
            I => \N__24938\
        );

    \I__5844\ : ClkMux
    port map (
            O => \N__25225\,
            I => \N__24938\
        );

    \I__5843\ : ClkMux
    port map (
            O => \N__25224\,
            I => \N__24938\
        );

    \I__5842\ : ClkMux
    port map (
            O => \N__25223\,
            I => \N__24938\
        );

    \I__5841\ : ClkMux
    port map (
            O => \N__25222\,
            I => \N__24938\
        );

    \I__5840\ : ClkMux
    port map (
            O => \N__25221\,
            I => \N__24938\
        );

    \I__5839\ : ClkMux
    port map (
            O => \N__25220\,
            I => \N__24938\
        );

    \I__5838\ : ClkMux
    port map (
            O => \N__25219\,
            I => \N__24938\
        );

    \I__5837\ : ClkMux
    port map (
            O => \N__25218\,
            I => \N__24938\
        );

    \I__5836\ : ClkMux
    port map (
            O => \N__25217\,
            I => \N__24938\
        );

    \I__5835\ : ClkMux
    port map (
            O => \N__25216\,
            I => \N__24938\
        );

    \I__5834\ : ClkMux
    port map (
            O => \N__25215\,
            I => \N__24938\
        );

    \I__5833\ : ClkMux
    port map (
            O => \N__25214\,
            I => \N__24938\
        );

    \I__5832\ : ClkMux
    port map (
            O => \N__25213\,
            I => \N__24938\
        );

    \I__5831\ : ClkMux
    port map (
            O => \N__25212\,
            I => \N__24938\
        );

    \I__5830\ : ClkMux
    port map (
            O => \N__25211\,
            I => \N__24938\
        );

    \I__5829\ : ClkMux
    port map (
            O => \N__25210\,
            I => \N__24938\
        );

    \I__5828\ : ClkMux
    port map (
            O => \N__25209\,
            I => \N__24938\
        );

    \I__5827\ : ClkMux
    port map (
            O => \N__25208\,
            I => \N__24938\
        );

    \I__5826\ : ClkMux
    port map (
            O => \N__25207\,
            I => \N__24938\
        );

    \I__5825\ : ClkMux
    port map (
            O => \N__25206\,
            I => \N__24938\
        );

    \I__5824\ : ClkMux
    port map (
            O => \N__25205\,
            I => \N__24938\
        );

    \I__5823\ : ClkMux
    port map (
            O => \N__25204\,
            I => \N__24938\
        );

    \I__5822\ : ClkMux
    port map (
            O => \N__25203\,
            I => \N__24938\
        );

    \I__5821\ : ClkMux
    port map (
            O => \N__25202\,
            I => \N__24938\
        );

    \I__5820\ : ClkMux
    port map (
            O => \N__25201\,
            I => \N__24938\
        );

    \I__5819\ : ClkMux
    port map (
            O => \N__25200\,
            I => \N__24938\
        );

    \I__5818\ : ClkMux
    port map (
            O => \N__25199\,
            I => \N__24938\
        );

    \I__5817\ : ClkMux
    port map (
            O => \N__25198\,
            I => \N__24938\
        );

    \I__5816\ : ClkMux
    port map (
            O => \N__25197\,
            I => \N__24938\
        );

    \I__5815\ : ClkMux
    port map (
            O => \N__25196\,
            I => \N__24938\
        );

    \I__5814\ : ClkMux
    port map (
            O => \N__25195\,
            I => \N__24938\
        );

    \I__5813\ : ClkMux
    port map (
            O => \N__25194\,
            I => \N__24938\
        );

    \I__5812\ : ClkMux
    port map (
            O => \N__25193\,
            I => \N__24938\
        );

    \I__5811\ : ClkMux
    port map (
            O => \N__25192\,
            I => \N__24938\
        );

    \I__5810\ : ClkMux
    port map (
            O => \N__25191\,
            I => \N__24938\
        );

    \I__5809\ : ClkMux
    port map (
            O => \N__25190\,
            I => \N__24938\
        );

    \I__5808\ : ClkMux
    port map (
            O => \N__25189\,
            I => \N__24938\
        );

    \I__5807\ : ClkMux
    port map (
            O => \N__25188\,
            I => \N__24938\
        );

    \I__5806\ : ClkMux
    port map (
            O => \N__25187\,
            I => \N__24938\
        );

    \I__5805\ : ClkMux
    port map (
            O => \N__25186\,
            I => \N__24938\
        );

    \I__5804\ : ClkMux
    port map (
            O => \N__25185\,
            I => \N__24938\
        );

    \I__5803\ : ClkMux
    port map (
            O => \N__25184\,
            I => \N__24938\
        );

    \I__5802\ : ClkMux
    port map (
            O => \N__25183\,
            I => \N__24938\
        );

    \I__5801\ : GlobalMux
    port map (
            O => \N__24938\,
            I => \N__24935\
        );

    \I__5800\ : gio2CtrlBuf
    port map (
            O => \N__24935\,
            I => clk_system_c_g
        );

    \I__5799\ : CascadeMux
    port map (
            O => \N__24932\,
            I => \N__24924\
        );

    \I__5798\ : CascadeMux
    port map (
            O => \N__24931\,
            I => \N__24921\
        );

    \I__5797\ : CascadeMux
    port map (
            O => \N__24930\,
            I => \N__24913\
        );

    \I__5796\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24892\
        );

    \I__5795\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24889\
        );

    \I__5794\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24886\
        );

    \I__5793\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24881\
        );

    \I__5792\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24881\
        );

    \I__5791\ : InMux
    port map (
            O => \N__24920\,
            I => \N__24878\
        );

    \I__5790\ : InMux
    port map (
            O => \N__24919\,
            I => \N__24875\
        );

    \I__5789\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24872\
        );

    \I__5788\ : InMux
    port map (
            O => \N__24917\,
            I => \N__24869\
        );

    \I__5787\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24862\
        );

    \I__5786\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24862\
        );

    \I__5785\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24862\
        );

    \I__5784\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24859\
        );

    \I__5783\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24856\
        );

    \I__5782\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24853\
        );

    \I__5781\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24850\
        );

    \I__5780\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24847\
        );

    \I__5779\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24842\
        );

    \I__5778\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24842\
        );

    \I__5777\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24839\
        );

    \I__5776\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24836\
        );

    \I__5775\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24833\
        );

    \I__5774\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24830\
        );

    \I__5773\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24827\
        );

    \I__5772\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24824\
        );

    \I__5771\ : InMux
    port map (
            O => \N__24898\,
            I => \N__24821\
        );

    \I__5770\ : InMux
    port map (
            O => \N__24897\,
            I => \N__24816\
        );

    \I__5769\ : InMux
    port map (
            O => \N__24896\,
            I => \N__24816\
        );

    \I__5768\ : InMux
    port map (
            O => \N__24895\,
            I => \N__24813\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__24892\,
            I => \N__24737\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__24889\,
            I => \N__24734\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__24886\,
            I => \N__24731\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__24881\,
            I => \N__24728\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__24878\,
            I => \N__24725\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__24875\,
            I => \N__24722\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__24872\,
            I => \N__24719\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__24869\,
            I => \N__24716\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__24862\,
            I => \N__24713\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__24859\,
            I => \N__24710\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__24856\,
            I => \N__24707\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__24853\,
            I => \N__24704\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__24850\,
            I => \N__24701\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__24847\,
            I => \N__24698\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__24842\,
            I => \N__24695\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__24839\,
            I => \N__24692\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__24836\,
            I => \N__24689\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__24833\,
            I => \N__24686\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__24830\,
            I => \N__24683\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__24827\,
            I => \N__24680\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__24824\,
            I => \N__24677\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__24821\,
            I => \N__24674\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__24816\,
            I => \N__24671\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__24813\,
            I => \N__24668\
        );

    \I__5743\ : SRMux
    port map (
            O => \N__24812\,
            I => \N__24473\
        );

    \I__5742\ : SRMux
    port map (
            O => \N__24811\,
            I => \N__24473\
        );

    \I__5741\ : SRMux
    port map (
            O => \N__24810\,
            I => \N__24473\
        );

    \I__5740\ : SRMux
    port map (
            O => \N__24809\,
            I => \N__24473\
        );

    \I__5739\ : SRMux
    port map (
            O => \N__24808\,
            I => \N__24473\
        );

    \I__5738\ : SRMux
    port map (
            O => \N__24807\,
            I => \N__24473\
        );

    \I__5737\ : SRMux
    port map (
            O => \N__24806\,
            I => \N__24473\
        );

    \I__5736\ : SRMux
    port map (
            O => \N__24805\,
            I => \N__24473\
        );

    \I__5735\ : SRMux
    port map (
            O => \N__24804\,
            I => \N__24473\
        );

    \I__5734\ : SRMux
    port map (
            O => \N__24803\,
            I => \N__24473\
        );

    \I__5733\ : SRMux
    port map (
            O => \N__24802\,
            I => \N__24473\
        );

    \I__5732\ : SRMux
    port map (
            O => \N__24801\,
            I => \N__24473\
        );

    \I__5731\ : SRMux
    port map (
            O => \N__24800\,
            I => \N__24473\
        );

    \I__5730\ : SRMux
    port map (
            O => \N__24799\,
            I => \N__24473\
        );

    \I__5729\ : SRMux
    port map (
            O => \N__24798\,
            I => \N__24473\
        );

    \I__5728\ : SRMux
    port map (
            O => \N__24797\,
            I => \N__24473\
        );

    \I__5727\ : SRMux
    port map (
            O => \N__24796\,
            I => \N__24473\
        );

    \I__5726\ : SRMux
    port map (
            O => \N__24795\,
            I => \N__24473\
        );

    \I__5725\ : SRMux
    port map (
            O => \N__24794\,
            I => \N__24473\
        );

    \I__5724\ : SRMux
    port map (
            O => \N__24793\,
            I => \N__24473\
        );

    \I__5723\ : SRMux
    port map (
            O => \N__24792\,
            I => \N__24473\
        );

    \I__5722\ : SRMux
    port map (
            O => \N__24791\,
            I => \N__24473\
        );

    \I__5721\ : SRMux
    port map (
            O => \N__24790\,
            I => \N__24473\
        );

    \I__5720\ : SRMux
    port map (
            O => \N__24789\,
            I => \N__24473\
        );

    \I__5719\ : SRMux
    port map (
            O => \N__24788\,
            I => \N__24473\
        );

    \I__5718\ : SRMux
    port map (
            O => \N__24787\,
            I => \N__24473\
        );

    \I__5717\ : SRMux
    port map (
            O => \N__24786\,
            I => \N__24473\
        );

    \I__5716\ : SRMux
    port map (
            O => \N__24785\,
            I => \N__24473\
        );

    \I__5715\ : SRMux
    port map (
            O => \N__24784\,
            I => \N__24473\
        );

    \I__5714\ : SRMux
    port map (
            O => \N__24783\,
            I => \N__24473\
        );

    \I__5713\ : SRMux
    port map (
            O => \N__24782\,
            I => \N__24473\
        );

    \I__5712\ : SRMux
    port map (
            O => \N__24781\,
            I => \N__24473\
        );

    \I__5711\ : SRMux
    port map (
            O => \N__24780\,
            I => \N__24473\
        );

    \I__5710\ : SRMux
    port map (
            O => \N__24779\,
            I => \N__24473\
        );

    \I__5709\ : SRMux
    port map (
            O => \N__24778\,
            I => \N__24473\
        );

    \I__5708\ : SRMux
    port map (
            O => \N__24777\,
            I => \N__24473\
        );

    \I__5707\ : SRMux
    port map (
            O => \N__24776\,
            I => \N__24473\
        );

    \I__5706\ : SRMux
    port map (
            O => \N__24775\,
            I => \N__24473\
        );

    \I__5705\ : SRMux
    port map (
            O => \N__24774\,
            I => \N__24473\
        );

    \I__5704\ : SRMux
    port map (
            O => \N__24773\,
            I => \N__24473\
        );

    \I__5703\ : SRMux
    port map (
            O => \N__24772\,
            I => \N__24473\
        );

    \I__5702\ : SRMux
    port map (
            O => \N__24771\,
            I => \N__24473\
        );

    \I__5701\ : SRMux
    port map (
            O => \N__24770\,
            I => \N__24473\
        );

    \I__5700\ : SRMux
    port map (
            O => \N__24769\,
            I => \N__24473\
        );

    \I__5699\ : SRMux
    port map (
            O => \N__24768\,
            I => \N__24473\
        );

    \I__5698\ : SRMux
    port map (
            O => \N__24767\,
            I => \N__24473\
        );

    \I__5697\ : SRMux
    port map (
            O => \N__24766\,
            I => \N__24473\
        );

    \I__5696\ : SRMux
    port map (
            O => \N__24765\,
            I => \N__24473\
        );

    \I__5695\ : SRMux
    port map (
            O => \N__24764\,
            I => \N__24473\
        );

    \I__5694\ : SRMux
    port map (
            O => \N__24763\,
            I => \N__24473\
        );

    \I__5693\ : SRMux
    port map (
            O => \N__24762\,
            I => \N__24473\
        );

    \I__5692\ : SRMux
    port map (
            O => \N__24761\,
            I => \N__24473\
        );

    \I__5691\ : SRMux
    port map (
            O => \N__24760\,
            I => \N__24473\
        );

    \I__5690\ : SRMux
    port map (
            O => \N__24759\,
            I => \N__24473\
        );

    \I__5689\ : SRMux
    port map (
            O => \N__24758\,
            I => \N__24473\
        );

    \I__5688\ : SRMux
    port map (
            O => \N__24757\,
            I => \N__24473\
        );

    \I__5687\ : SRMux
    port map (
            O => \N__24756\,
            I => \N__24473\
        );

    \I__5686\ : SRMux
    port map (
            O => \N__24755\,
            I => \N__24473\
        );

    \I__5685\ : SRMux
    port map (
            O => \N__24754\,
            I => \N__24473\
        );

    \I__5684\ : SRMux
    port map (
            O => \N__24753\,
            I => \N__24473\
        );

    \I__5683\ : SRMux
    port map (
            O => \N__24752\,
            I => \N__24473\
        );

    \I__5682\ : SRMux
    port map (
            O => \N__24751\,
            I => \N__24473\
        );

    \I__5681\ : SRMux
    port map (
            O => \N__24750\,
            I => \N__24473\
        );

    \I__5680\ : SRMux
    port map (
            O => \N__24749\,
            I => \N__24473\
        );

    \I__5679\ : SRMux
    port map (
            O => \N__24748\,
            I => \N__24473\
        );

    \I__5678\ : SRMux
    port map (
            O => \N__24747\,
            I => \N__24473\
        );

    \I__5677\ : SRMux
    port map (
            O => \N__24746\,
            I => \N__24473\
        );

    \I__5676\ : SRMux
    port map (
            O => \N__24745\,
            I => \N__24473\
        );

    \I__5675\ : SRMux
    port map (
            O => \N__24744\,
            I => \N__24473\
        );

    \I__5674\ : SRMux
    port map (
            O => \N__24743\,
            I => \N__24473\
        );

    \I__5673\ : SRMux
    port map (
            O => \N__24742\,
            I => \N__24473\
        );

    \I__5672\ : SRMux
    port map (
            O => \N__24741\,
            I => \N__24473\
        );

    \I__5671\ : SRMux
    port map (
            O => \N__24740\,
            I => \N__24473\
        );

    \I__5670\ : Glb2LocalMux
    port map (
            O => \N__24737\,
            I => \N__24473\
        );

    \I__5669\ : Glb2LocalMux
    port map (
            O => \N__24734\,
            I => \N__24473\
        );

    \I__5668\ : Glb2LocalMux
    port map (
            O => \N__24731\,
            I => \N__24473\
        );

    \I__5667\ : Glb2LocalMux
    port map (
            O => \N__24728\,
            I => \N__24473\
        );

    \I__5666\ : Glb2LocalMux
    port map (
            O => \N__24725\,
            I => \N__24473\
        );

    \I__5665\ : Glb2LocalMux
    port map (
            O => \N__24722\,
            I => \N__24473\
        );

    \I__5664\ : Glb2LocalMux
    port map (
            O => \N__24719\,
            I => \N__24473\
        );

    \I__5663\ : Glb2LocalMux
    port map (
            O => \N__24716\,
            I => \N__24473\
        );

    \I__5662\ : Glb2LocalMux
    port map (
            O => \N__24713\,
            I => \N__24473\
        );

    \I__5661\ : Glb2LocalMux
    port map (
            O => \N__24710\,
            I => \N__24473\
        );

    \I__5660\ : Glb2LocalMux
    port map (
            O => \N__24707\,
            I => \N__24473\
        );

    \I__5659\ : Glb2LocalMux
    port map (
            O => \N__24704\,
            I => \N__24473\
        );

    \I__5658\ : Glb2LocalMux
    port map (
            O => \N__24701\,
            I => \N__24473\
        );

    \I__5657\ : Glb2LocalMux
    port map (
            O => \N__24698\,
            I => \N__24473\
        );

    \I__5656\ : Glb2LocalMux
    port map (
            O => \N__24695\,
            I => \N__24473\
        );

    \I__5655\ : Glb2LocalMux
    port map (
            O => \N__24692\,
            I => \N__24473\
        );

    \I__5654\ : Glb2LocalMux
    port map (
            O => \N__24689\,
            I => \N__24473\
        );

    \I__5653\ : Glb2LocalMux
    port map (
            O => \N__24686\,
            I => \N__24473\
        );

    \I__5652\ : Glb2LocalMux
    port map (
            O => \N__24683\,
            I => \N__24473\
        );

    \I__5651\ : Glb2LocalMux
    port map (
            O => \N__24680\,
            I => \N__24473\
        );

    \I__5650\ : Glb2LocalMux
    port map (
            O => \N__24677\,
            I => \N__24473\
        );

    \I__5649\ : Glb2LocalMux
    port map (
            O => \N__24674\,
            I => \N__24473\
        );

    \I__5648\ : Glb2LocalMux
    port map (
            O => \N__24671\,
            I => \N__24473\
        );

    \I__5647\ : Glb2LocalMux
    port map (
            O => \N__24668\,
            I => \N__24473\
        );

    \I__5646\ : GlobalMux
    port map (
            O => \N__24473\,
            I => \N__24470\
        );

    \I__5645\ : gio2CtrlBuf
    port map (
            O => \N__24470\,
            I => reset_system_g
        );

    \I__5644\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__24464\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\
        );

    \I__5642\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24456\
        );

    \I__5641\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24453\
        );

    \I__5640\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24450\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__24456\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__24453\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__24450\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__24443\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_\
        );

    \I__5635\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24435\
        );

    \I__5634\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24432\
        );

    \I__5633\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24429\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__24435\,
            I => \N__24426\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__24432\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__24429\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5629\ : Odrv4
    port map (
            O => \N__24426\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__24419\,
            I => \ppm_encoder_1.N_148_17_cascade_\
        );

    \I__5627\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24413\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__5625\ : Odrv12
    port map (
            O => \N__24410\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\
        );

    \I__5624\ : InMux
    port map (
            O => \N__24407\,
            I => \N__24401\
        );

    \I__5623\ : InMux
    port map (
            O => \N__24406\,
            I => \N__24401\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__24401\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\
        );

    \I__5621\ : InMux
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__24395\,
            I => \ppm_encoder_1.N_148_17\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__24392\,
            I => \N__24389\
        );

    \I__5618\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__24386\,
            I => \N__24383\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__24383\,
            I => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\
        );

    \I__5615\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24377\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__24377\,
            I => \N__24374\
        );

    \I__5613\ : Span12Mux_v
    port map (
            O => \N__24374\,
            I => \N__24371\
        );

    \I__5612\ : Odrv12
    port map (
            O => \N__24371\,
            I => \ppm_encoder_1.N_148\
        );

    \I__5611\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24363\
        );

    \I__5610\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24360\
        );

    \I__5609\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24357\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__24363\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__24360\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__24357\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5605\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24345\
        );

    \I__5604\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24342\
        );

    \I__5603\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24339\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__24345\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__24342\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__24339\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5599\ : CascadeMux
    port map (
            O => \N__24332\,
            I => \N__24328\
        );

    \I__5598\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24324\
        );

    \I__5597\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24321\
        );

    \I__5596\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24318\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__24324\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__24321\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__24318\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5592\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24306\
        );

    \I__5591\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24303\
        );

    \I__5590\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24300\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__24306\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__24303\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__24300\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5586\ : InMux
    port map (
            O => \N__24293\,
            I => \N__24287\
        );

    \I__5585\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24287\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__24287\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__24284\,
            I => \N__24281\
        );

    \I__5582\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24275\
        );

    \I__5581\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24275\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__5578\ : Span4Mux_v
    port map (
            O => \N__24269\,
            I => \N__24265\
        );

    \I__5577\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24262\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__24265\,
            I => \ppm_encoder_1.N_241\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__24262\,
            I => \ppm_encoder_1.N_241\
        );

    \I__5574\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24253\
        );

    \I__5573\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24249\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__24253\,
            I => \N__24246\
        );

    \I__5571\ : InMux
    port map (
            O => \N__24252\,
            I => \N__24243\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__24249\,
            I => \N__24240\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__24246\,
            I => \N__24236\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__24243\,
            I => \N__24233\
        );

    \I__5567\ : Span4Mux_v
    port map (
            O => \N__24240\,
            I => \N__24230\
        );

    \I__5566\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24227\
        );

    \I__5565\ : Span4Mux_v
    port map (
            O => \N__24236\,
            I => \N__24222\
        );

    \I__5564\ : Span4Mux_s2_v
    port map (
            O => \N__24233\,
            I => \N__24222\
        );

    \I__5563\ : Odrv4
    port map (
            O => \N__24230\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__24227\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__24222\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5560\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24207\
        );

    \I__5559\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24204\
        );

    \I__5558\ : IoInMux
    port map (
            O => \N__24213\,
            I => \N__24200\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__24212\,
            I => \N__24196\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__24211\,
            I => \N__24188\
        );

    \I__5555\ : CascadeMux
    port map (
            O => \N__24210\,
            I => \N__24185\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__24207\,
            I => \N__24181\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__24204\,
            I => \N__24178\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__24203\,
            I => \N__24174\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__24200\,
            I => \N__24170\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__24199\,
            I => \N__24165\
        );

    \I__5549\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24160\
        );

    \I__5548\ : InMux
    port map (
            O => \N__24195\,
            I => \N__24160\
        );

    \I__5547\ : InMux
    port map (
            O => \N__24194\,
            I => \N__24157\
        );

    \I__5546\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24154\
        );

    \I__5545\ : InMux
    port map (
            O => \N__24192\,
            I => \N__24151\
        );

    \I__5544\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24148\
        );

    \I__5543\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24141\
        );

    \I__5542\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24141\
        );

    \I__5541\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24141\
        );

    \I__5540\ : Span4Mux_v
    port map (
            O => \N__24181\,
            I => \N__24136\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__24178\,
            I => \N__24136\
        );

    \I__5538\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24133\
        );

    \I__5537\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24130\
        );

    \I__5536\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24127\
        );

    \I__5535\ : IoSpan4Mux
    port map (
            O => \N__24170\,
            I => \N__24124\
        );

    \I__5534\ : CascadeMux
    port map (
            O => \N__24169\,
            I => \N__24121\
        );

    \I__5533\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24111\
        );

    \I__5532\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24111\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__24160\,
            I => \N__24106\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__24157\,
            I => \N__24106\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24101\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__24151\,
            I => \N__24101\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__24148\,
            I => \N__24098\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__24141\,
            I => \N__24091\
        );

    \I__5525\ : Sp12to4
    port map (
            O => \N__24136\,
            I => \N__24091\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__24133\,
            I => \N__24091\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24088\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24085\
        );

    \I__5521\ : Sp12to4
    port map (
            O => \N__24124\,
            I => \N__24082\
        );

    \I__5520\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24077\
        );

    \I__5519\ : InMux
    port map (
            O => \N__24120\,
            I => \N__24077\
        );

    \I__5518\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24072\
        );

    \I__5517\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24072\
        );

    \I__5516\ : InMux
    port map (
            O => \N__24117\,
            I => \N__24067\
        );

    \I__5515\ : InMux
    port map (
            O => \N__24116\,
            I => \N__24067\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__24111\,
            I => \N__24064\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__24106\,
            I => \N__24061\
        );

    \I__5512\ : Span4Mux_h
    port map (
            O => \N__24101\,
            I => \N__24056\
        );

    \I__5511\ : Span4Mux_s3_h
    port map (
            O => \N__24098\,
            I => \N__24056\
        );

    \I__5510\ : Span12Mux_h
    port map (
            O => \N__24091\,
            I => \N__24051\
        );

    \I__5509\ : Span12Mux_h
    port map (
            O => \N__24088\,
            I => \N__24051\
        );

    \I__5508\ : Span12Mux_h
    port map (
            O => \N__24085\,
            I => \N__24046\
        );

    \I__5507\ : Span12Mux_s9_v
    port map (
            O => \N__24082\,
            I => \N__24046\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__24077\,
            I => reset_system
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__24072\,
            I => reset_system
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__24067\,
            I => reset_system
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__24064\,
            I => reset_system
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__24061\,
            I => reset_system
        );

    \I__5501\ : Odrv4
    port map (
            O => \N__24056\,
            I => reset_system
        );

    \I__5500\ : Odrv12
    port map (
            O => \N__24051\,
            I => reset_system
        );

    \I__5499\ : Odrv12
    port map (
            O => \N__24046\,
            I => reset_system
        );

    \I__5498\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24024\
        );

    \I__5497\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24020\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__24027\,
            I => \N__24016\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__24024\,
            I => \N__24013\
        );

    \I__5494\ : InMux
    port map (
            O => \N__24023\,
            I => \N__24010\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__24007\
        );

    \I__5492\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24002\
        );

    \I__5491\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24002\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__24013\,
            I => \N__23999\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__24010\,
            I => \N__23996\
        );

    \I__5488\ : Span4Mux_h
    port map (
            O => \N__24007\,
            I => \N__23991\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23986\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__23999\,
            I => \N__23986\
        );

    \I__5485\ : Span12Mux_s7_v
    port map (
            O => \N__23996\,
            I => \N__23983\
        );

    \I__5484\ : InMux
    port map (
            O => \N__23995\,
            I => \N__23978\
        );

    \I__5483\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23978\
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__23991\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5481\ : Odrv4
    port map (
            O => \N__23986\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5480\ : Odrv12
    port map (
            O => \N__23983\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__23978\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5478\ : IoInMux
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__23966\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\
        );

    \I__5476\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23960\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__23960\,
            I => \N__23957\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__23954\,
            I => \N__23950\
        );

    \I__5472\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23947\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__23950\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_2\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__23947\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_2\
        );

    \I__5469\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23939\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__5467\ : Span4Mux_h
    port map (
            O => \N__23936\,
            I => \N__23933\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__23933\,
            I => \N__23928\
        );

    \I__5465\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23925\
        );

    \I__5464\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23922\
        );

    \I__5463\ : Odrv4
    port map (
            O => \N__23928\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__23925\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__23922\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\
        );

    \I__5460\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23910\
        );

    \I__5459\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23905\
        );

    \I__5458\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23905\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23895\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__23905\,
            I => \N__23892\
        );

    \I__5455\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23889\
        );

    \I__5454\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23876\
        );

    \I__5453\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23876\
        );

    \I__5452\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23876\
        );

    \I__5451\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23876\
        );

    \I__5450\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23876\
        );

    \I__5449\ : InMux
    port map (
            O => \N__23898\,
            I => \N__23876\
        );

    \I__5448\ : Odrv12
    port map (
            O => \N__23895\,
            I => \uart_frame_decoder.N_85\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__23892\,
            I => \uart_frame_decoder.N_85\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__23889\,
            I => \uart_frame_decoder.N_85\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__23876\,
            I => \uart_frame_decoder.N_85\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__23867\,
            I => \N__23863\
        );

    \I__5443\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23860\
        );

    \I__5442\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23854\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__23857\,
            I => \N__23849\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__23854\,
            I => \N__23849\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__23849\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__5437\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23842\
        );

    \I__5436\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__23842\,
            I => \N__23836\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__23839\,
            I => \uart_frame_decoder.state_1Z0Z_4\
        );

    \I__5433\ : Odrv12
    port map (
            O => \N__23836\,
            I => \uart_frame_decoder.state_1Z0Z_4\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__23831\,
            I => \N__23828\
        );

    \I__5431\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23813\
        );

    \I__5430\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23808\
        );

    \I__5429\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23808\
        );

    \I__5428\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23801\
        );

    \I__5427\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23801\
        );

    \I__5426\ : InMux
    port map (
            O => \N__23823\,
            I => \N__23801\
        );

    \I__5425\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23798\
        );

    \I__5424\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23793\
        );

    \I__5423\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23793\
        );

    \I__5422\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23789\
        );

    \I__5421\ : CascadeMux
    port map (
            O => \N__23818\,
            I => \N__23784\
        );

    \I__5420\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23779\
        );

    \I__5419\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23779\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__23813\,
            I => \N__23772\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__23808\,
            I => \N__23772\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23772\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23769\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__23793\,
            I => \N__23766\
        );

    \I__5413\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23763\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__23789\,
            I => \N__23760\
        );

    \I__5411\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23757\
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__23787\,
            I => \N__23754\
        );

    \I__5409\ : InMux
    port map (
            O => \N__23784\,
            I => \N__23751\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__23779\,
            I => \N__23744\
        );

    \I__5407\ : Span4Mux_v
    port map (
            O => \N__23772\,
            I => \N__23744\
        );

    \I__5406\ : Span4Mux_h
    port map (
            O => \N__23769\,
            I => \N__23744\
        );

    \I__5405\ : Span4Mux_h
    port map (
            O => \N__23766\,
            I => \N__23739\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__23763\,
            I => \N__23739\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__23760\,
            I => \N__23734\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__23757\,
            I => \N__23734\
        );

    \I__5401\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23731\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__23751\,
            I => \N__23726\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__23744\,
            I => \N__23726\
        );

    \I__5398\ : Span4Mux_v
    port map (
            O => \N__23739\,
            I => \N__23721\
        );

    \I__5397\ : Span4Mux_h
    port map (
            O => \N__23734\,
            I => \N__23721\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__23731\,
            I => uart_pc_data_rdy
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__23726\,
            I => uart_pc_data_rdy
        );

    \I__5394\ : Odrv4
    port map (
            O => \N__23721\,
            I => uart_pc_data_rdy
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__23714\,
            I => \N__23702\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__23713\,
            I => \N__23695\
        );

    \I__5391\ : InMux
    port map (
            O => \N__23712\,
            I => \N__23664\
        );

    \I__5390\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23664\
        );

    \I__5389\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23664\
        );

    \I__5388\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23664\
        );

    \I__5387\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23664\
        );

    \I__5386\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23657\
        );

    \I__5385\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23657\
        );

    \I__5384\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23657\
        );

    \I__5383\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23644\
        );

    \I__5382\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23644\
        );

    \I__5381\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23644\
        );

    \I__5380\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23644\
        );

    \I__5379\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23641\
        );

    \I__5378\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23638\
        );

    \I__5377\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23635\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__23693\,
            I => \N__23632\
        );

    \I__5375\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23618\
        );

    \I__5374\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23618\
        );

    \I__5373\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23618\
        );

    \I__5372\ : InMux
    port map (
            O => \N__23689\,
            I => \N__23618\
        );

    \I__5371\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23607\
        );

    \I__5370\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23607\
        );

    \I__5369\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23607\
        );

    \I__5368\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23607\
        );

    \I__5367\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23607\
        );

    \I__5366\ : InMux
    port map (
            O => \N__23683\,
            I => \N__23602\
        );

    \I__5365\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23602\
        );

    \I__5364\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23595\
        );

    \I__5363\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23595\
        );

    \I__5362\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23595\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__23678\,
            I => \N__23585\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__23677\,
            I => \N__23582\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__23676\,
            I => \N__23579\
        );

    \I__5358\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23576\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__23664\,
            I => \N__23573\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23569\
        );

    \I__5355\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23560\
        );

    \I__5354\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23560\
        );

    \I__5353\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23560\
        );

    \I__5352\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23560\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__23644\,
            I => \N__23557\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__23641\,
            I => \N__23550\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23545\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__23635\,
            I => \N__23545\
        );

    \I__5347\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23540\
        );

    \I__5346\ : InMux
    port map (
            O => \N__23631\,
            I => \N__23540\
        );

    \I__5345\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23531\
        );

    \I__5344\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23531\
        );

    \I__5343\ : InMux
    port map (
            O => \N__23628\,
            I => \N__23531\
        );

    \I__5342\ : InMux
    port map (
            O => \N__23627\,
            I => \N__23531\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__23618\,
            I => \N__23522\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__23607\,
            I => \N__23522\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__23602\,
            I => \N__23522\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23522\
        );

    \I__5337\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23513\
        );

    \I__5336\ : InMux
    port map (
            O => \N__23593\,
            I => \N__23513\
        );

    \I__5335\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23513\
        );

    \I__5334\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23513\
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__23590\,
            I => \N__23500\
        );

    \I__5332\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23496\
        );

    \I__5331\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23493\
        );

    \I__5330\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23486\
        );

    \I__5329\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23486\
        );

    \I__5328\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23486\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__23576\,
            I => \N__23481\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__23573\,
            I => \N__23481\
        );

    \I__5325\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23478\
        );

    \I__5324\ : Span4Mux_v
    port map (
            O => \N__23569\,
            I => \N__23471\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__23560\,
            I => \N__23471\
        );

    \I__5322\ : Span4Mux_h
    port map (
            O => \N__23557\,
            I => \N__23471\
        );

    \I__5321\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23462\
        );

    \I__5320\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23462\
        );

    \I__5319\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23462\
        );

    \I__5318\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23462\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__23550\,
            I => \N__23455\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__23545\,
            I => \N__23455\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__23540\,
            I => \N__23455\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23448\
        );

    \I__5313\ : Span4Mux_v
    port map (
            O => \N__23522\,
            I => \N__23448\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__23513\,
            I => \N__23448\
        );

    \I__5311\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23443\
        );

    \I__5310\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23443\
        );

    \I__5309\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23430\
        );

    \I__5308\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23430\
        );

    \I__5307\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23430\
        );

    \I__5306\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23430\
        );

    \I__5305\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23430\
        );

    \I__5304\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23430\
        );

    \I__5303\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23421\
        );

    \I__5302\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23421\
        );

    \I__5301\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23421\
        );

    \I__5300\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23421\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__23496\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__23493\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__23486\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__23481\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__23478\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__23471\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__23462\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__23455\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__23448\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__23443\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__23430\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__23421\,
            I => \ppm_encoder_1.PPM_STATE_62_d\
        );

    \I__5287\ : InMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__5285\ : Span12Mux_s10_v
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__5284\ : Odrv12
    port map (
            O => \N__23387\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\
        );

    \I__5283\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__23375\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__23372\,
            I => \N__23369\
        );

    \I__5278\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23366\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__23366\,
            I => \ppm_encoder_1.pulses2countZ0Z_7\
        );

    \I__5276\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__5274\ : Odrv4
    port map (
            O => \N__23357\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\
        );

    \I__5273\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23351\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__23351\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\
        );

    \I__5271\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__23345\,
            I => \ppm_encoder_1.pulses2countZ0Z_6\
        );

    \I__5269\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23336\
        );

    \I__5267\ : Span4Mux_v
    port map (
            O => \N__23336\,
            I => \N__23333\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__5265\ : Sp12to4
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__5264\ : Odrv12
    port map (
            O => \N__23327\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\
        );

    \I__5263\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__23321\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\
        );

    \I__5261\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__23315\,
            I => \ppm_encoder_1.pulses2countZ0Z_12\
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__23312\,
            I => \N__23305\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__23311\,
            I => \N__23302\
        );

    \I__5257\ : InMux
    port map (
            O => \N__23310\,
            I => \N__23296\
        );

    \I__5256\ : InMux
    port map (
            O => \N__23309\,
            I => \N__23293\
        );

    \I__5255\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23290\
        );

    \I__5254\ : InMux
    port map (
            O => \N__23305\,
            I => \N__23281\
        );

    \I__5253\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23281\
        );

    \I__5252\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23281\
        );

    \I__5251\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23281\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__23299\,
            I => \N__23278\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__23296\,
            I => \N__23266\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__23293\,
            I => \N__23266\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__23290\,
            I => \N__23266\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__23281\,
            I => \N__23266\
        );

    \I__5245\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23263\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__23277\,
            I => \N__23260\
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__23276\,
            I => \N__23255\
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__23275\,
            I => \N__23252\
        );

    \I__5241\ : Span4Mux_v
    port map (
            O => \N__23266\,
            I => \N__23246\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__23263\,
            I => \N__23246\
        );

    \I__5239\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23237\
        );

    \I__5238\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23237\
        );

    \I__5237\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23237\
        );

    \I__5236\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23237\
        );

    \I__5235\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23232\
        );

    \I__5234\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23232\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__23246\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__23237\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__23232\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__5230\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23216\
        );

    \I__5229\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23213\
        );

    \I__5228\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23202\
        );

    \I__5227\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23193\
        );

    \I__5226\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23193\
        );

    \I__5225\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23193\
        );

    \I__5224\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23193\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__23216\,
            I => \N__23187\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__23213\,
            I => \N__23187\
        );

    \I__5221\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23184\
        );

    \I__5220\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23181\
        );

    \I__5219\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23172\
        );

    \I__5218\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23172\
        );

    \I__5217\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23172\
        );

    \I__5216\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23172\
        );

    \I__5215\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23167\
        );

    \I__5214\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23167\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23161\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__23193\,
            I => \N__23161\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__23192\,
            I => \N__23157\
        );

    \I__5210\ : Span4Mux_v
    port map (
            O => \N__23187\,
            I => \N__23145\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__23184\,
            I => \N__23145\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__23181\,
            I => \N__23145\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23145\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__23167\,
            I => \N__23145\
        );

    \I__5205\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23142\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__23161\,
            I => \N__23139\
        );

    \I__5203\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23132\
        );

    \I__5202\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23132\
        );

    \I__5201\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23132\
        );

    \I__5200\ : Span4Mux_v
    port map (
            O => \N__23145\,
            I => \N__23129\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__23142\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__23139\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__23132\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__23129\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__5194\ : InMux
    port map (
            O => \N__23117\,
            I => \N__23113\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__23116\,
            I => \N__23110\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__23113\,
            I => \N__23105\
        );

    \I__5191\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23098\
        );

    \I__5190\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23098\
        );

    \I__5189\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23098\
        );

    \I__5188\ : Span4Mux_v
    port map (
            O => \N__23105\,
            I => \N__23093\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__23093\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__23093\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__5185\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23087\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__23087\,
            I => \N__23083\
        );

    \I__5183\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23080\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__23083\,
            I => \N__23076\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__23073\
        );

    \I__5180\ : InMux
    port map (
            O => \N__23079\,
            I => \N__23070\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__23076\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__23073\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__23070\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__5176\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__23060\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\
        );

    \I__5174\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23052\
        );

    \I__5173\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23049\
        );

    \I__5172\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23046\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23043\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__23049\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__23046\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__23043\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5167\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23031\
        );

    \I__5166\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23028\
        );

    \I__5165\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23025\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__23031\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__23028\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__23025\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5161\ : CascadeMux
    port map (
            O => \N__23018\,
            I => \N__23013\
        );

    \I__5160\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23010\
        );

    \I__5159\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23007\
        );

    \I__5158\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23004\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__23010\,
            I => \N__23001\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__23007\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__23004\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__23001\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5153\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22989\
        );

    \I__5152\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22986\
        );

    \I__5151\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22983\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__22989\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__22986\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__22983\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__5147\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22971\
        );

    \I__5146\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22968\
        );

    \I__5145\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22965\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__22971\,
            I => \N__22962\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__22968\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__22965\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5141\ : Odrv4
    port map (
            O => \N__22962\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5140\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22950\
        );

    \I__5139\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22947\
        );

    \I__5138\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22944\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22941\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__22947\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__22944\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__22941\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__22934\,
            I => \N__22929\
        );

    \I__5132\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22926\
        );

    \I__5131\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22923\
        );

    \I__5130\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22920\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__22926\,
            I => \N__22917\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__22923\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__22920\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__22917\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5125\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22907\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__22907\,
            I => \N__22902\
        );

    \I__5123\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22899\
        );

    \I__5122\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22896\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__22902\,
            I => \N__22893\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__22899\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__22896\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5118\ : Odrv4
    port map (
            O => \N__22893\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5117\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22883\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__22883\,
            I => \N__22878\
        );

    \I__5115\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22875\
        );

    \I__5114\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22872\
        );

    \I__5113\ : Span4Mux_h
    port map (
            O => \N__22878\,
            I => \N__22869\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__22875\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__22872\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__22869\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__5109\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22857\
        );

    \I__5108\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22854\
        );

    \I__5107\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22851\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22848\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__22854\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__22851\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5103\ : Odrv4
    port map (
            O => \N__22848\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5102\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22834\
        );

    \I__5101\ : CascadeMux
    port map (
            O => \N__22840\,
            I => \N__22831\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__22839\,
            I => \N__22828\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__22838\,
            I => \N__22816\
        );

    \I__5098\ : InMux
    port map (
            O => \N__22837\,
            I => \N__22810\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__22834\,
            I => \N__22807\
        );

    \I__5096\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22800\
        );

    \I__5095\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22800\
        );

    \I__5094\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22800\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__22826\,
            I => \N__22797\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__22825\,
            I => \N__22793\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__22824\,
            I => \N__22788\
        );

    \I__5090\ : CascadeMux
    port map (
            O => \N__22823\,
            I => \N__22783\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__22822\,
            I => \N__22780\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__22821\,
            I => \N__22776\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__22820\,
            I => \N__22773\
        );

    \I__5086\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22761\
        );

    \I__5085\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22761\
        );

    \I__5084\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22761\
        );

    \I__5083\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22761\
        );

    \I__5082\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22756\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__22810\,
            I => \N__22753\
        );

    \I__5080\ : Span4Mux_v
    port map (
            O => \N__22807\,
            I => \N__22747\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__22800\,
            I => \N__22744\
        );

    \I__5078\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22735\
        );

    \I__5077\ : InMux
    port map (
            O => \N__22796\,
            I => \N__22735\
        );

    \I__5076\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22735\
        );

    \I__5075\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22735\
        );

    \I__5074\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22724\
        );

    \I__5073\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22724\
        );

    \I__5072\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22724\
        );

    \I__5071\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22724\
        );

    \I__5070\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22724\
        );

    \I__5069\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22719\
        );

    \I__5068\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22719\
        );

    \I__5067\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22712\
        );

    \I__5066\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22712\
        );

    \I__5065\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22712\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__22771\,
            I => \N__22709\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__22770\,
            I => \N__22706\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__22761\,
            I => \N__22701\
        );

    \I__5061\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22696\
        );

    \I__5060\ : InMux
    port map (
            O => \N__22759\,
            I => \N__22696\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__22756\,
            I => \N__22688\
        );

    \I__5058\ : Span4Mux_s3_v
    port map (
            O => \N__22753\,
            I => \N__22688\
        );

    \I__5057\ : CascadeMux
    port map (
            O => \N__22752\,
            I => \N__22684\
        );

    \I__5056\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22678\
        );

    \I__5055\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22678\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__22747\,
            I => \N__22665\
        );

    \I__5053\ : Span4Mux_s3_v
    port map (
            O => \N__22744\,
            I => \N__22665\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22665\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__22724\,
            I => \N__22665\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__22719\,
            I => \N__22665\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__22712\,
            I => \N__22665\
        );

    \I__5048\ : InMux
    port map (
            O => \N__22709\,
            I => \N__22656\
        );

    \I__5047\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22656\
        );

    \I__5046\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22656\
        );

    \I__5045\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22656\
        );

    \I__5044\ : Span4Mux_v
    port map (
            O => \N__22701\,
            I => \N__22651\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__22696\,
            I => \N__22651\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__22695\,
            I => \N__22646\
        );

    \I__5041\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22643\
        );

    \I__5040\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22640\
        );

    \I__5039\ : Span4Mux_v
    port map (
            O => \N__22688\,
            I => \N__22637\
        );

    \I__5038\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22634\
        );

    \I__5037\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22629\
        );

    \I__5036\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22629\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__22678\,
            I => \N__22622\
        );

    \I__5034\ : Span4Mux_v
    port map (
            O => \N__22665\,
            I => \N__22622\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22622\
        );

    \I__5032\ : Span4Mux_h
    port map (
            O => \N__22651\,
            I => \N__22619\
        );

    \I__5031\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22614\
        );

    \I__5030\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22614\
        );

    \I__5029\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22611\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__22643\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__22640\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5026\ : Odrv4
    port map (
            O => \N__22637\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__22634\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__22629\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__22622\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__22619\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__22614\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__22611\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__5019\ : InMux
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__5017\ : Span4Mux_h
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__22583\,
            I => \ppm_encoder_1.N_301\
        );

    \I__5015\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22577\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22574\
        );

    \I__5013\ : Sp12to4
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__5012\ : Span12Mux_s7_v
    port map (
            O => \N__22571\,
            I => \N__22566\
        );

    \I__5011\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22561\
        );

    \I__5010\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22561\
        );

    \I__5009\ : Odrv12
    port map (
            O => \N__22566\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__22561\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__5007\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__22550\,
            I => \N__22545\
        );

    \I__5004\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22540\
        );

    \I__5003\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22540\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__22545\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__22540\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__5000\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__22532\,
            I => \N__22527\
        );

    \I__4998\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22524\
        );

    \I__4997\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22521\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__22527\,
            I => \N__22516\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__22524\,
            I => \N__22516\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__22521\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__22516\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__4992\ : CascadeMux
    port map (
            O => \N__22511\,
            I => \N__22507\
        );

    \I__4991\ : CascadeMux
    port map (
            O => \N__22510\,
            I => \N__22504\
        );

    \I__4990\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22499\
        );

    \I__4989\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22494\
        );

    \I__4988\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22494\
        );

    \I__4987\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22491\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22486\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22486\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22483\
        );

    \I__4983\ : Span4Mux_h
    port map (
            O => \N__22486\,
            I => \N__22480\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__22483\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__22480\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__4980\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22472\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__4978\ : Span4Mux_h
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__22466\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\
        );

    \I__4976\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22455\
        );

    \I__4974\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22450\
        );

    \I__4973\ : InMux
    port map (
            O => \N__22458\,
            I => \N__22450\
        );

    \I__4972\ : Odrv12
    port map (
            O => \N__22455\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__22450\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__4970\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22440\
        );

    \I__4969\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22437\
        );

    \I__4968\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22434\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__22440\,
            I => \N__22431\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22428\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__22434\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__4964\ : Odrv12
    port map (
            O => \N__22431\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__22428\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \ppm_encoder_1.N_323_cascade_\
        );

    \I__4961\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22410\
        );

    \I__4959\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22405\
        );

    \I__4958\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22405\
        );

    \I__4957\ : Odrv12
    port map (
            O => \N__22410\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__22405\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4955\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22393\
        );

    \I__4953\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22390\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__22393\,
            I => \N__22384\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__22390\,
            I => \N__22384\
        );

    \I__4950\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22381\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__22384\,
            I => \N__22378\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__22381\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__22378\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4946\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__22370\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\
        );

    \I__4944\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__22364\,
            I => \ppm_encoder_1.N_322\
        );

    \I__4942\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__4940\ : Span4Mux_v
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__22352\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\
        );

    \I__4938\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22341\
        );

    \I__4936\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22336\
        );

    \I__4935\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22336\
        );

    \I__4934\ : Odrv12
    port map (
            O => \N__22341\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__22336\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4932\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22327\
        );

    \I__4931\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22324\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__22327\,
            I => \N__22321\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22318\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__22321\,
            I => \N__22314\
        );

    \I__4927\ : Span4Mux_v
    port map (
            O => \N__22318\,
            I => \N__22311\
        );

    \I__4926\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22308\
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__22314\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__22311\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__22308\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__22301\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7_cascade_\
        );

    \I__4921\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__22295\,
            I => \N__22291\
        );

    \I__4919\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__4918\ : Span4Mux_v
    port map (
            O => \N__22291\,
            I => \N__22285\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__22288\,
            I => \N__22282\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__22285\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__4915\ : Odrv12
    port map (
            O => \N__22282\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__4914\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__22274\,
            I => \ppm_encoder_1.N_309\
        );

    \I__4912\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22267\
        );

    \I__4911\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22264\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__22267\,
            I => \N__22261\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__22264\,
            I => \N__22258\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__22261\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__4907\ : Odrv4
    port map (
            O => \N__22258\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__4906\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22246\
        );

    \I__4904\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22243\
        );

    \I__4903\ : Span4Mux_v
    port map (
            O => \N__22246\,
            I => \N__22234\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__22243\,
            I => \N__22234\
        );

    \I__4901\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22230\
        );

    \I__4900\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22227\
        );

    \I__4899\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22224\
        );

    \I__4898\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22221\
        );

    \I__4897\ : Span4Mux_h
    port map (
            O => \N__22234\,
            I => \N__22218\
        );

    \I__4896\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22215\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__22230\,
            I => \N__22210\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22210\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__22224\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__22221\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__22218\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__22215\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__22210\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__4888\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__22196\,
            I => \N__22191\
        );

    \I__4886\ : CascadeMux
    port map (
            O => \N__22195\,
            I => \N__22185\
        );

    \I__4885\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22182\
        );

    \I__4884\ : Span4Mux_h
    port map (
            O => \N__22191\,
            I => \N__22179\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22176\
        );

    \I__4882\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22171\
        );

    \I__4881\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22171\
        );

    \I__4880\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22168\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__22182\,
            I => \N__22165\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__22179\,
            I => \N__22162\
        );

    \I__4877\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22159\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__22171\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__22168\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4874\ : Odrv12
    port map (
            O => \N__22165\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4873\ : Odrv4
    port map (
            O => \N__22162\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__22159\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__22148\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\
        );

    \I__4870\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__4868\ : Span4Mux_h
    port map (
            O => \N__22139\,
            I => \N__22133\
        );

    \I__4867\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22128\
        );

    \I__4866\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22128\
        );

    \I__4865\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22125\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__22133\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__22128\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__22125\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__4861\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__22115\,
            I => \N__22112\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__4858\ : Span4Mux_v
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__22106\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__22103\,
            I => \N__22099\
        );

    \I__4855\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22095\
        );

    \I__4854\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22090\
        );

    \I__4853\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22090\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__22095\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__22090\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__4850\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__22082\,
            I => \N__22078\
        );

    \I__4848\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22075\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__22078\,
            I => \N__22070\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__22075\,
            I => \N__22070\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__4844\ : Odrv4
    port map (
            O => \N__22067\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__4843\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__22058\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\
        );

    \I__4840\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22051\
        );

    \I__4839\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22048\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__22051\,
            I => \N__22043\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__22048\,
            I => \N__22043\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__22043\,
            I => \N__22039\
        );

    \I__4835\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22036\
        );

    \I__4834\ : Span4Mux_v
    port map (
            O => \N__22039\,
            I => \N__22033\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__22036\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__22033\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__4831\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__22025\,
            I => \N__22021\
        );

    \I__4829\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22018\
        );

    \I__4828\ : Span4Mux_h
    port map (
            O => \N__22021\,
            I => \N__22014\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__22011\
        );

    \I__4826\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22008\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__22014\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__4824\ : Odrv12
    port map (
            O => \N__22011\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__22008\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__4822\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__4820\ : Span4Mux_s2_v
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__21989\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\
        );

    \I__4817\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21982\
        );

    \I__4816\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21979\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__21982\,
            I => \N__21976\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__21979\,
            I => \N__21973\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__21976\,
            I => \N__21970\
        );

    \I__4812\ : Odrv12
    port map (
            O => \N__21973\,
            I => scaler_1_data_13
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__21970\,
            I => scaler_1_data_13
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__21965\,
            I => \N__21961\
        );

    \I__4809\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21956\
        );

    \I__4808\ : InMux
    port map (
            O => \N__21961\,
            I => \N__21956\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__21956\,
            I => \N__21945\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__21955\,
            I => \N__21942\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__21954\,
            I => \N__21939\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__21953\,
            I => \N__21936\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__21952\,
            I => \N__21933\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__21951\,
            I => \N__21930\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__21950\,
            I => \N__21927\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__21949\,
            I => \N__21924\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__21948\,
            I => \N__21917\
        );

    \I__4798\ : Span4Mux_v
    port map (
            O => \N__21945\,
            I => \N__21913\
        );

    \I__4797\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21904\
        );

    \I__4796\ : InMux
    port map (
            O => \N__21939\,
            I => \N__21904\
        );

    \I__4795\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21904\
        );

    \I__4794\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21904\
        );

    \I__4793\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21897\
        );

    \I__4792\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21897\
        );

    \I__4791\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21897\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__21923\,
            I => \N__21894\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__21922\,
            I => \N__21890\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__21921\,
            I => \N__21887\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__21920\,
            I => \N__21884\
        );

    \I__4786\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21881\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__21916\,
            I => \N__21878\
        );

    \I__4784\ : Span4Mux_s1_v
    port map (
            O => \N__21913\,
            I => \N__21871\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__21904\,
            I => \N__21871\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__21897\,
            I => \N__21871\
        );

    \I__4781\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21868\
        );

    \I__4780\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21863\
        );

    \I__4779\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21863\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21860\
        );

    \I__4777\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21857\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21854\
        );

    \I__4775\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21851\
        );

    \I__4774\ : Sp12to4
    port map (
            O => \N__21871\,
            I => \N__21843\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__21868\,
            I => \N__21843\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21840\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__21860\,
            I => \N__21835\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21835\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__21854\,
            I => \N__21830\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__21851\,
            I => \N__21830\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__21850\,
            I => \N__21827\
        );

    \I__4766\ : InMux
    port map (
            O => \N__21849\,
            I => \N__21824\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__21848\,
            I => \N__21821\
        );

    \I__4764\ : Span12Mux_s11_v
    port map (
            O => \N__21843\,
            I => \N__21818\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__21840\,
            I => \N__21815\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__21835\,
            I => \N__21810\
        );

    \I__4761\ : Span4Mux_v
    port map (
            O => \N__21830\,
            I => \N__21810\
        );

    \I__4760\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21807\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21804\
        );

    \I__4758\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21801\
        );

    \I__4757\ : Odrv12
    port map (
            O => \N__21818\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__21815\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__21810\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__21807\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4753\ : Odrv12
    port map (
            O => \N__21804\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__21801\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4751\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__21776\,
            I => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\
        );

    \I__4746\ : InMux
    port map (
            O => \N__21773\,
            I => \ppm_encoder_1.un1_throttle_cry_12\
        );

    \I__4745\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__21764\,
            I => scaler_1_data_14
        );

    \I__4742\ : InMux
    port map (
            O => \N__21761\,
            I => \bfn_12_18_0_\
        );

    \I__4741\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21754\
        );

    \I__4740\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21751\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__21754\,
            I => \N__21746\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__21751\,
            I => \N__21746\
        );

    \I__4737\ : Span4Mux_v
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__21743\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__4735\ : CEMux
    port map (
            O => \N__21740\,
            I => \N__21735\
        );

    \I__4734\ : CEMux
    port map (
            O => \N__21739\,
            I => \N__21732\
        );

    \I__4733\ : CEMux
    port map (
            O => \N__21738\,
            I => \N__21727\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21723\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__21732\,
            I => \N__21720\
        );

    \I__4730\ : CEMux
    port map (
            O => \N__21731\,
            I => \N__21717\
        );

    \I__4729\ : CEMux
    port map (
            O => \N__21730\,
            I => \N__21714\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21711\
        );

    \I__4727\ : CEMux
    port map (
            O => \N__21726\,
            I => \N__21708\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__21723\,
            I => \N__21700\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__21720\,
            I => \N__21700\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__21717\,
            I => \N__21700\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__21714\,
            I => \N__21697\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__21711\,
            I => \N__21694\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__21708\,
            I => \N__21691\
        );

    \I__4720\ : CEMux
    port map (
            O => \N__21707\,
            I => \N__21688\
        );

    \I__4719\ : Sp12to4
    port map (
            O => \N__21700\,
            I => \N__21685\
        );

    \I__4718\ : Span4Mux_h
    port map (
            O => \N__21697\,
            I => \N__21680\
        );

    \I__4717\ : Span4Mux_h
    port map (
            O => \N__21694\,
            I => \N__21680\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__21691\,
            I => \N__21675\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__21688\,
            I => \N__21675\
        );

    \I__4714\ : Odrv12
    port map (
            O => \N__21685\,
            I => \ppm_encoder_1.scaler_1_dv_0\
        );

    \I__4713\ : Odrv4
    port map (
            O => \N__21680\,
            I => \ppm_encoder_1.scaler_1_dv_0\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__21675\,
            I => \ppm_encoder_1.scaler_1_dv_0\
        );

    \I__4711\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__21662\,
            I => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\
        );

    \I__4708\ : InMux
    port map (
            O => \N__21659\,
            I => \N__21656\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__21656\,
            I => \N__21652\
        );

    \I__4706\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21649\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__21652\,
            I => \N__21644\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__21649\,
            I => \N__21644\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__21644\,
            I => scaler_1_data_8
        );

    \I__4702\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21637\
        );

    \I__4701\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21634\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__21637\,
            I => \N__21630\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__21634\,
            I => \N__21627\
        );

    \I__4698\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21624\
        );

    \I__4697\ : Span4Mux_h
    port map (
            O => \N__21630\,
            I => \N__21621\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__21627\,
            I => \N__21618\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__21624\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__21621\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__21618\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__4692\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__21608\,
            I => \N__21604\
        );

    \I__4690\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21601\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__21604\,
            I => \N__21596\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__21601\,
            I => \N__21596\
        );

    \I__4687\ : Span4Mux_v
    port map (
            O => \N__21596\,
            I => \N__21593\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__21593\,
            I => scaler_4_data_11
        );

    \I__4685\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__21584\,
            I => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\
        );

    \I__4682\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__21578\,
            I => \N__21575\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__21575\,
            I => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\
        );

    \I__4679\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21569\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21565\
        );

    \I__4677\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21562\
        );

    \I__4676\ : Span4Mux_h
    port map (
            O => \N__21565\,
            I => \N__21559\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21556\
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__21559\,
            I => scaler_1_data_10
        );

    \I__4673\ : Odrv12
    port map (
            O => \N__21556\,
            I => scaler_1_data_10
        );

    \I__4672\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21544\
        );

    \I__4671\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21544\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__21549\,
            I => \N__21541\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__21544\,
            I => \N__21538\
        );

    \I__4668\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21535\
        );

    \I__4667\ : Span4Mux_v
    port map (
            O => \N__21538\,
            I => \N__21532\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__21535\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__21532\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4664\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__21524\,
            I => \N__21520\
        );

    \I__4662\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__21520\,
            I => \N__21514\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__21517\,
            I => \N__21511\
        );

    \I__4659\ : Span4Mux_v
    port map (
            O => \N__21514\,
            I => \N__21506\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__21511\,
            I => \N__21506\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__21506\,
            I => scaler_4_data_12
        );

    \I__4656\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21500\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__4653\ : Odrv4
    port map (
            O => \N__21494\,
            I => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\
        );

    \I__4652\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__21488\,
            I => \ppm_encoder_1.N_143_0\
        );

    \I__4650\ : CascadeMux
    port map (
            O => \N__21485\,
            I => \N__21482\
        );

    \I__4649\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21478\
        );

    \I__4648\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21475\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__21478\,
            I => \N__21472\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__21475\,
            I => \N__21469\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__21472\,
            I => \N__21464\
        );

    \I__4644\ : Span4Mux_h
    port map (
            O => \N__21469\,
            I => \N__21461\
        );

    \I__4643\ : CascadeMux
    port map (
            O => \N__21468\,
            I => \N__21458\
        );

    \I__4642\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21455\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__21464\,
            I => \N__21450\
        );

    \I__4640\ : Span4Mux_v
    port map (
            O => \N__21461\,
            I => \N__21450\
        );

    \I__4639\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21447\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__21455\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__21450\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__21447\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__4635\ : IoInMux
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__21437\,
            I => \N__21434\
        );

    \I__4633\ : IoSpan4Mux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__4632\ : Span4Mux_s2_v
    port map (
            O => \N__21431\,
            I => \N__21428\
        );

    \I__4631\ : Sp12to4
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__4630\ : Span12Mux_s10_v
    port map (
            O => \N__21425\,
            I => \N__21421\
        );

    \I__4629\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21418\
        );

    \I__4628\ : Odrv12
    port map (
            O => \N__21421\,
            I => ppm_output_c
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__21418\,
            I => ppm_output_c
        );

    \I__4626\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__4624\ : Odrv12
    port map (
            O => \N__21407\,
            I => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\
        );

    \I__4623\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__21401\,
            I => \N__21397\
        );

    \I__4621\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21394\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__21397\,
            I => \N__21391\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__21394\,
            I => \N__21388\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__21391\,
            I => scaler_1_data_9
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__21388\,
            I => scaler_1_data_9
        );

    \I__4616\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21376\
        );

    \I__4614\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21373\
        );

    \I__4613\ : Span4Mux_h
    port map (
            O => \N__21376\,
            I => \N__21370\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__21373\,
            I => \N__21367\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__21370\,
            I => \frame_decoder_CH3data_7\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__21367\,
            I => \frame_decoder_CH3data_7\
        );

    \I__4609\ : InMux
    port map (
            O => \N__21362\,
            I => \N__21358\
        );

    \I__4608\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21355\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__21358\,
            I => \N__21352\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__21355\,
            I => \N__21349\
        );

    \I__4605\ : Span4Mux_v
    port map (
            O => \N__21352\,
            I => \N__21346\
        );

    \I__4604\ : Span4Mux_v
    port map (
            O => \N__21349\,
            I => \N__21343\
        );

    \I__4603\ : Span4Mux_h
    port map (
            O => \N__21346\,
            I => \N__21338\
        );

    \I__4602\ : Span4Mux_h
    port map (
            O => \N__21343\,
            I => \N__21338\
        );

    \I__4601\ : Odrv4
    port map (
            O => \N__21338\,
            I => \uart_frame_decoder.source_CH1data_1_sqmuxa\
        );

    \I__4600\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21331\
        );

    \I__4599\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21328\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__21331\,
            I => \N__21325\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21322\
        );

    \I__4596\ : Odrv12
    port map (
            O => \N__21325\,
            I => scaler_1_data_6
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__21322\,
            I => scaler_1_data_6
        );

    \I__4594\ : InMux
    port map (
            O => \N__21317\,
            I => \N__21313\
        );

    \I__4593\ : InMux
    port map (
            O => \N__21316\,
            I => \N__21310\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__21313\,
            I => \N__21307\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__21310\,
            I => \N__21304\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__21307\,
            I => scaler_1_data_7
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__21304\,
            I => scaler_1_data_7
        );

    \I__4588\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21296\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__21296\,
            I => \N__21293\
        );

    \I__4586\ : Span4Mux_h
    port map (
            O => \N__21293\,
            I => \N__21290\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__21290\,
            I => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\
        );

    \I__4584\ : InMux
    port map (
            O => \N__21287\,
            I => \ppm_encoder_1.un1_throttle_cry_6\
        );

    \I__4583\ : InMux
    port map (
            O => \N__21284\,
            I => \ppm_encoder_1.un1_throttle_cry_7\
        );

    \I__4582\ : InMux
    port map (
            O => \N__21281\,
            I => \ppm_encoder_1.un1_throttle_cry_8\
        );

    \I__4581\ : InMux
    port map (
            O => \N__21278\,
            I => \ppm_encoder_1.un1_throttle_cry_9\
        );

    \I__4580\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21271\
        );

    \I__4579\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21268\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__21271\,
            I => \N__21265\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21262\
        );

    \I__4576\ : Odrv12
    port map (
            O => \N__21265\,
            I => scaler_1_data_11
        );

    \I__4575\ : Odrv12
    port map (
            O => \N__21262\,
            I => scaler_1_data_11
        );

    \I__4574\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__21248\,
            I => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\
        );

    \I__4570\ : InMux
    port map (
            O => \N__21245\,
            I => \ppm_encoder_1.un1_throttle_cry_10\
        );

    \I__4569\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21235\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__21238\,
            I => \N__21232\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__21235\,
            I => \N__21229\
        );

    \I__4565\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__4564\ : Span4Mux_v
    port map (
            O => \N__21229\,
            I => \N__21221\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21221\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__21221\,
            I => scaler_1_data_12
        );

    \I__4561\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__21209\,
            I => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\
        );

    \I__4557\ : InMux
    port map (
            O => \N__21206\,
            I => \ppm_encoder_1.un1_throttle_cry_11\
        );

    \I__4556\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21199\
        );

    \I__4555\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21196\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__21199\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__21196\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__4551\ : InMux
    port map (
            O => \N__21188\,
            I => \N__21185\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__21185\,
            I => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\
        );

    \I__4549\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__21179\,
            I => \N__21175\
        );

    \I__4547\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21172\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__21175\,
            I => \N__21167\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__21172\,
            I => \N__21167\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__21164\,
            I => scaler_4_data_13
        );

    \I__4542\ : InMux
    port map (
            O => \N__21161\,
            I => \bfn_12_14_0_\
        );

    \I__4541\ : InMux
    port map (
            O => \N__21158\,
            I => \scaler_4.un2_source_data_0_cry_9\
        );

    \I__4540\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N__21149\
        );

    \I__4538\ : Span4Mux_v
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__21146\,
            I => scaler_4_data_14
        );

    \I__4536\ : CEMux
    port map (
            O => \N__21143\,
            I => \N__21116\
        );

    \I__4535\ : CEMux
    port map (
            O => \N__21142\,
            I => \N__21116\
        );

    \I__4534\ : CEMux
    port map (
            O => \N__21141\,
            I => \N__21116\
        );

    \I__4533\ : CEMux
    port map (
            O => \N__21140\,
            I => \N__21116\
        );

    \I__4532\ : CEMux
    port map (
            O => \N__21139\,
            I => \N__21116\
        );

    \I__4531\ : CEMux
    port map (
            O => \N__21138\,
            I => \N__21116\
        );

    \I__4530\ : CEMux
    port map (
            O => \N__21137\,
            I => \N__21116\
        );

    \I__4529\ : CEMux
    port map (
            O => \N__21136\,
            I => \N__21116\
        );

    \I__4528\ : CEMux
    port map (
            O => \N__21135\,
            I => \N__21116\
        );

    \I__4527\ : GlobalMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__4526\ : gio2CtrlBuf
    port map (
            O => \N__21113\,
            I => pc_frame_decoder_dv_0_g
        );

    \I__4525\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21104\
        );

    \I__4524\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21098\
        );

    \I__4523\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21095\
        );

    \I__4522\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21091\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21088\
        );

    \I__4520\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21085\
        );

    \I__4519\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21082\
        );

    \I__4518\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21079\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__21098\,
            I => \N__21076\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21073\
        );

    \I__4515\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21070\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__21091\,
            I => \N__21066\
        );

    \I__4513\ : Span4Mux_v
    port map (
            O => \N__21088\,
            I => \N__21056\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21056\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__21082\,
            I => \N__21056\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__21079\,
            I => \N__21056\
        );

    \I__4509\ : Span4Mux_v
    port map (
            O => \N__21076\,
            I => \N__21049\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__21073\,
            I => \N__21049\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__21070\,
            I => \N__21049\
        );

    \I__4506\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21046\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__21066\,
            I => \N__21043\
        );

    \I__4504\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21040\
        );

    \I__4503\ : Span4Mux_v
    port map (
            O => \N__21056\,
            I => \N__21033\
        );

    \I__4502\ : Span4Mux_h
    port map (
            O => \N__21049\,
            I => \N__21033\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__21046\,
            I => \N__21033\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__21043\,
            I => uart_pc_data_0
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__21040\,
            I => uart_pc_data_0
        );

    \I__4498\ : Odrv4
    port map (
            O => \N__21033\,
            I => uart_pc_data_0
        );

    \I__4497\ : InMux
    port map (
            O => \N__21026\,
            I => \N__21022\
        );

    \I__4496\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21019\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__21022\,
            I => \N__21012\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__21019\,
            I => \N__21012\
        );

    \I__4493\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21009\
        );

    \I__4492\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21006\
        );

    \I__4491\ : Span4Mux_v
    port map (
            O => \N__21012\,
            I => \N__21001\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__21009\,
            I => \N__21001\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__21006\,
            I => \N__20998\
        );

    \I__4488\ : Span4Mux_h
    port map (
            O => \N__21001\,
            I => \N__20995\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__20998\,
            I => \frame_decoder_CH3data_0\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__20995\,
            I => \frame_decoder_CH3data_0\
        );

    \I__4485\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20985\
        );

    \I__4484\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20982\
        );

    \I__4483\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20977\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__20985\,
            I => \N__20971\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__20982\,
            I => \N__20968\
        );

    \I__4480\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20965\
        );

    \I__4479\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20962\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__20977\,
            I => \N__20959\
        );

    \I__4477\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20956\
        );

    \I__4476\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20952\
        );

    \I__4475\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20949\
        );

    \I__4474\ : Span4Mux_v
    port map (
            O => \N__20971\,
            I => \N__20942\
        );

    \I__4473\ : Span4Mux_v
    port map (
            O => \N__20968\,
            I => \N__20942\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__20965\,
            I => \N__20942\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__20962\,
            I => \N__20935\
        );

    \I__4470\ : Span4Mux_h
    port map (
            O => \N__20959\,
            I => \N__20935\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20935\
        );

    \I__4468\ : InMux
    port map (
            O => \N__20955\,
            I => \N__20932\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20927\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20927\
        );

    \I__4465\ : Span4Mux_h
    port map (
            O => \N__20942\,
            I => \N__20924\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__20935\,
            I => \N__20921\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__20932\,
            I => \N__20918\
        );

    \I__4462\ : Odrv12
    port map (
            O => \N__20927\,
            I => uart_pc_data_1
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__20924\,
            I => uart_pc_data_1
        );

    \I__4460\ : Odrv4
    port map (
            O => \N__20921\,
            I => uart_pc_data_1
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__20918\,
            I => uart_pc_data_1
        );

    \I__4458\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__20903\,
            I => \frame_decoder_CH3data_1\
        );

    \I__4455\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20894\
        );

    \I__4454\ : InMux
    port map (
            O => \N__20899\,
            I => \N__20889\
        );

    \I__4453\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20886\
        );

    \I__4452\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20883\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20879\
        );

    \I__4450\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20876\
        );

    \I__4449\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20873\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20865\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__20886\,
            I => \N__20865\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__20883\,
            I => \N__20865\
        );

    \I__4445\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20862\
        );

    \I__4444\ : Span4Mux_h
    port map (
            O => \N__20879\,
            I => \N__20855\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__20876\,
            I => \N__20855\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20855\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20852\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__20865\,
            I => \N__20845\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__20862\,
            I => \N__20845\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__20855\,
            I => \N__20842\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__20852\,
            I => \N__20839\
        );

    \I__4436\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20836\
        );

    \I__4435\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20833\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__20845\,
            I => uart_pc_data_2
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__20842\,
            I => uart_pc_data_2
        );

    \I__4432\ : Odrv12
    port map (
            O => \N__20839\,
            I => uart_pc_data_2
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__20836\,
            I => uart_pc_data_2
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__20833\,
            I => uart_pc_data_2
        );

    \I__4429\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__20816\,
            I => \frame_decoder_CH3data_2\
        );

    \I__4426\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20805\
        );

    \I__4425\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20802\
        );

    \I__4424\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20799\
        );

    \I__4423\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20795\
        );

    \I__4422\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20792\
        );

    \I__4421\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20789\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20781\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__20802\,
            I => \N__20781\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20781\
        );

    \I__4417\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20778\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__20795\,
            I => \N__20773\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__20792\,
            I => \N__20773\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__20789\,
            I => \N__20770\
        );

    \I__4413\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20767\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__20781\,
            I => \N__20761\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20761\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__20773\,
            I => \N__20758\
        );

    \I__4409\ : Span12Mux_v
    port map (
            O => \N__20770\,
            I => \N__20753\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__20767\,
            I => \N__20753\
        );

    \I__4407\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20750\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__20761\,
            I => uart_pc_data_3
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__20758\,
            I => uart_pc_data_3
        );

    \I__4404\ : Odrv12
    port map (
            O => \N__20753\,
            I => uart_pc_data_3
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__20750\,
            I => uart_pc_data_3
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__4401\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__20732\,
            I => \frame_decoder_CH3data_3\
        );

    \I__4398\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20722\
        );

    \I__4397\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20717\
        );

    \I__4396\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20713\
        );

    \I__4395\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20710\
        );

    \I__4394\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20707\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20704\
        );

    \I__4392\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20701\
        );

    \I__4391\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20698\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__20717\,
            I => \N__20695\
        );

    \I__4389\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20692\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20685\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__20710\,
            I => \N__20685\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__20707\,
            I => \N__20685\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__20704\,
            I => \N__20682\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__20701\,
            I => \N__20679\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__20698\,
            I => \N__20674\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__20695\,
            I => \N__20674\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__20692\,
            I => \N__20670\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__20685\,
            I => \N__20667\
        );

    \I__4379\ : Span4Mux_h
    port map (
            O => \N__20682\,
            I => \N__20664\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__20679\,
            I => \N__20659\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__20674\,
            I => \N__20659\
        );

    \I__4376\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20656\
        );

    \I__4375\ : Odrv12
    port map (
            O => \N__20670\,
            I => uart_pc_data_4
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__20667\,
            I => uart_pc_data_4
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__20664\,
            I => uart_pc_data_4
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__20659\,
            I => uart_pc_data_4
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__20656\,
            I => uart_pc_data_4
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__4369\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20639\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__4367\ : Odrv4
    port map (
            O => \N__20636\,
            I => \frame_decoder_CH3data_4\
        );

    \I__4366\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20628\
        );

    \I__4365\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20625\
        );

    \I__4364\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20622\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__20628\,
            I => \N__20614\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__20625\,
            I => \N__20614\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20610\
        );

    \I__4360\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20607\
        );

    \I__4359\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20603\
        );

    \I__4358\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20600\
        );

    \I__4357\ : Span4Mux_v
    port map (
            O => \N__20614\,
            I => \N__20596\
        );

    \I__4356\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20593\
        );

    \I__4355\ : Span4Mux_v
    port map (
            O => \N__20610\,
            I => \N__20588\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20588\
        );

    \I__4353\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20585\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__20603\,
            I => \N__20580\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__20600\,
            I => \N__20580\
        );

    \I__4350\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20577\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__20596\,
            I => \N__20574\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__20593\,
            I => \N__20571\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__20588\,
            I => \N__20568\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20565\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__20580\,
            I => \N__20560\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20560\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__20574\,
            I => uart_pc_data_6
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__20571\,
            I => uart_pc_data_6
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__20568\,
            I => uart_pc_data_6
        );

    \I__4340\ : Odrv12
    port map (
            O => \N__20565\,
            I => uart_pc_data_6
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__20560\,
            I => uart_pc_data_6
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__4337\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20543\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__20543\,
            I => \N__20540\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__20540\,
            I => \frame_decoder_CH3data_6\
        );

    \I__4334\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20532\
        );

    \I__4333\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20528\
        );

    \I__4332\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20523\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__20532\,
            I => \N__20520\
        );

    \I__4330\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20517\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20514\
        );

    \I__4328\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20511\
        );

    \I__4327\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20508\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__20523\,
            I => \N__20502\
        );

    \I__4325\ : Span4Mux_v
    port map (
            O => \N__20520\,
            I => \N__20497\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__20517\,
            I => \N__20497\
        );

    \I__4323\ : Span4Mux_v
    port map (
            O => \N__20514\,
            I => \N__20490\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__20511\,
            I => \N__20490\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20490\
        );

    \I__4320\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20487\
        );

    \I__4319\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20484\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__20505\,
            I => \N__20480\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__20502\,
            I => \N__20477\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__20497\,
            I => \N__20470\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__20490\,
            I => \N__20470\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__20487\,
            I => \N__20470\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__20484\,
            I => \N__20467\
        );

    \I__4312\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20464\
        );

    \I__4311\ : InMux
    port map (
            O => \N__20480\,
            I => \N__20461\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__20477\,
            I => uart_pc_data_7
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__20470\,
            I => uart_pc_data_7
        );

    \I__4308\ : Odrv12
    port map (
            O => \N__20467\,
            I => uart_pc_data_7
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__20464\,
            I => uart_pc_data_7
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__20461\,
            I => uart_pc_data_7
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__4304\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__20444\,
            I => \scaler_4.un2_source_data_0_cry_1_c_RNO_2\
        );

    \I__4302\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20436\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__20440\,
            I => \N__20433\
        );

    \I__4300\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20429\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20426\
        );

    \I__4298\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20421\
        );

    \I__4297\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20421\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__20429\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__20426\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__20421\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__4293\ : InMux
    port map (
            O => \N__20414\,
            I => \scaler_4.un2_source_data_0_cry_1\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__4291\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20402\
        );

    \I__4290\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20402\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__20402\,
            I => \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__4287\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__20390\,
            I => \N__20386\
        );

    \I__4284\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20383\
        );

    \I__4283\ : Span4Mux_v
    port map (
            O => \N__20386\,
            I => \N__20380\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__20383\,
            I => \N__20377\
        );

    \I__4281\ : Span4Mux_v
    port map (
            O => \N__20380\,
            I => \N__20374\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__20377\,
            I => \N__20371\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__20374\,
            I => scaler_4_data_7
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__20371\,
            I => scaler_4_data_7
        );

    \I__4277\ : InMux
    port map (
            O => \N__20366\,
            I => \scaler_4.un2_source_data_0_cry_2\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__4275\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20354\
        );

    \I__4274\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20354\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__20354\,
            I => \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI\
        );

    \I__4272\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__20348\,
            I => \N__20344\
        );

    \I__4270\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20341\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__20344\,
            I => \N__20336\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__20341\,
            I => \N__20336\
        );

    \I__4267\ : Span4Mux_v
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__20333\,
            I => scaler_4_data_8
        );

    \I__4265\ : InMux
    port map (
            O => \N__20330\,
            I => \scaler_4.un2_source_data_0_cry_3\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__20327\,
            I => \N__20324\
        );

    \I__4263\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20318\
        );

    \I__4262\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20318\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__20318\,
            I => \scaler_4.un3_source_data_0_cry_3_c_RNI15MI\
        );

    \I__4260\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20308\
        );

    \I__4258\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20305\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__20308\,
            I => \N__20300\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__20305\,
            I => \N__20300\
        );

    \I__4255\ : Span4Mux_v
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__20297\,
            I => scaler_4_data_9
        );

    \I__4253\ : InMux
    port map (
            O => \N__20294\,
            I => \scaler_4.un2_source_data_0_cry_4\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__4251\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20282\
        );

    \I__4250\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20282\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__20282\,
            I => \scaler_4.un3_source_data_0_cry_4_c_RNI49NI\
        );

    \I__4248\ : InMux
    port map (
            O => \N__20279\,
            I => \N__20275\
        );

    \I__4247\ : InMux
    port map (
            O => \N__20278\,
            I => \N__20272\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__20275\,
            I => \N__20269\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__20272\,
            I => \N__20266\
        );

    \I__4244\ : Span12Mux_h
    port map (
            O => \N__20269\,
            I => \N__20263\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__20266\,
            I => \N__20260\
        );

    \I__4242\ : Odrv12
    port map (
            O => \N__20263\,
            I => scaler_4_data_10
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__20260\,
            I => scaler_4_data_10
        );

    \I__4240\ : InMux
    port map (
            O => \N__20255\,
            I => \scaler_4.un2_source_data_0_cry_5\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__4238\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20243\
        );

    \I__4237\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20243\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__20243\,
            I => \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI\
        );

    \I__4235\ : InMux
    port map (
            O => \N__20240\,
            I => \scaler_4.un2_source_data_0_cry_6\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__4233\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20228\
        );

    \I__4232\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20228\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__20228\,
            I => \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI\
        );

    \I__4230\ : InMux
    port map (
            O => \N__20225\,
            I => \scaler_4.un2_source_data_0_cry_7\
        );

    \I__4229\ : InMux
    port map (
            O => \N__20222\,
            I => \ppm_encoder_1.un1_counter_13_cry_11\
        );

    \I__4228\ : InMux
    port map (
            O => \N__20219\,
            I => \ppm_encoder_1.un1_counter_13_cry_12\
        );

    \I__4227\ : InMux
    port map (
            O => \N__20216\,
            I => \ppm_encoder_1.un1_counter_13_cry_13\
        );

    \I__4226\ : InMux
    port map (
            O => \N__20213\,
            I => \ppm_encoder_1.un1_counter_13_cry_14\
        );

    \I__4225\ : InMux
    port map (
            O => \N__20210\,
            I => \bfn_11_30_0_\
        );

    \I__4224\ : InMux
    port map (
            O => \N__20207\,
            I => \ppm_encoder_1.un1_counter_13_cry_16\
        );

    \I__4223\ : InMux
    port map (
            O => \N__20204\,
            I => \ppm_encoder_1.un1_counter_13_cry_17\
        );

    \I__4222\ : SRMux
    port map (
            O => \N__20201\,
            I => \N__20192\
        );

    \I__4221\ : SRMux
    port map (
            O => \N__20200\,
            I => \N__20192\
        );

    \I__4220\ : SRMux
    port map (
            O => \N__20199\,
            I => \N__20192\
        );

    \I__4219\ : GlobalMux
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__4218\ : gio2CtrlBuf
    port map (
            O => \N__20189\,
            I => \ppm_encoder_1.N_228_g\
        );

    \I__4217\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__4215\ : Span4Mux_s1_v
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__20177\,
            I => \N__20173\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__20176\,
            I => \N__20170\
        );

    \I__4212\ : Sp12to4
    port map (
            O => \N__20173\,
            I => \N__20162\
        );

    \I__4211\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20153\
        );

    \I__4210\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20153\
        );

    \I__4209\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20153\
        );

    \I__4208\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20153\
        );

    \I__4207\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20148\
        );

    \I__4206\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20148\
        );

    \I__4205\ : Span12Mux_s10_v
    port map (
            O => \N__20162\,
            I => \N__20145\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__20153\,
            I => pc_frame_decoder_dv
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__20148\,
            I => pc_frame_decoder_dv
        );

    \I__4202\ : Odrv12
    port map (
            O => \N__20145\,
            I => pc_frame_decoder_dv
        );

    \I__4201\ : IoInMux
    port map (
            O => \N__20138\,
            I => \N__20135\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__20135\,
            I => pc_frame_decoder_dv_0
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__4198\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__20126\,
            I => \frame_decoder_OFF4data_4\
        );

    \I__4196\ : CEMux
    port map (
            O => \N__20123\,
            I => \N__20120\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__20120\,
            I => \N__20116\
        );

    \I__4194\ : CEMux
    port map (
            O => \N__20119\,
            I => \N__20113\
        );

    \I__4193\ : Span4Mux_h
    port map (
            O => \N__20116\,
            I => \N__20110\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__20113\,
            I => \N__20107\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__20110\,
            I => \uart_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__20107\,
            I => \uart_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__20102\,
            I => \N__20097\
        );

    \I__4188\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20093\
        );

    \I__4187\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20088\
        );

    \I__4186\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20088\
        );

    \I__4185\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20085\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__20093\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__20088\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__20085\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4181\ : InMux
    port map (
            O => \N__20078\,
            I => \ppm_encoder_1.un1_counter_13_cry_2\
        );

    \I__4180\ : InMux
    port map (
            O => \N__20075\,
            I => \ppm_encoder_1.un1_counter_13_cry_3\
        );

    \I__4179\ : InMux
    port map (
            O => \N__20072\,
            I => \ppm_encoder_1.un1_counter_13_cry_4\
        );

    \I__4178\ : InMux
    port map (
            O => \N__20069\,
            I => \ppm_encoder_1.un1_counter_13_cry_5\
        );

    \I__4177\ : InMux
    port map (
            O => \N__20066\,
            I => \ppm_encoder_1.un1_counter_13_cry_6\
        );

    \I__4176\ : InMux
    port map (
            O => \N__20063\,
            I => \bfn_11_29_0_\
        );

    \I__4175\ : InMux
    port map (
            O => \N__20060\,
            I => \ppm_encoder_1.un1_counter_13_cry_8\
        );

    \I__4174\ : InMux
    port map (
            O => \N__20057\,
            I => \ppm_encoder_1.un1_counter_13_cry_9\
        );

    \I__4173\ : InMux
    port map (
            O => \N__20054\,
            I => \ppm_encoder_1.un1_counter_13_cry_10\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__20051\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1_cascade_\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__4170\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__20042\,
            I => \ppm_encoder_1.pulses2countZ0Z_1\
        );

    \I__4168\ : InMux
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__20036\,
            I => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\
        );

    \I__4166\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__4164\ : Span4Mux_v
    port map (
            O => \N__20027\,
            I => \N__20021\
        );

    \I__4163\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20014\
        );

    \I__4162\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20014\
        );

    \I__4161\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20014\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__20021\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__20014\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__4158\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20006\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__20006\,
            I => \ppm_encoder_1.pulses2countZ0Z_0\
        );

    \I__4156\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19999\
        );

    \I__4155\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19996\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__19999\,
            I => \N__19990\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__19996\,
            I => \N__19990\
        );

    \I__4152\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19985\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__19990\,
            I => \N__19982\
        );

    \I__4150\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19977\
        );

    \I__4149\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19977\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__19985\,
            I => \N__19974\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__19982\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__19977\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__19974\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__19967\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__4142\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__19958\,
            I => \ppm_encoder_1.pulses2countZ0Z_3\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__19955\,
            I => \N__19951\
        );

    \I__4139\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19948\
        );

    \I__4138\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19945\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19940\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__19945\,
            I => \N__19940\
        );

    \I__4135\ : Span12Mux_s8_v
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__4134\ : Odrv12
    port map (
            O => \N__19937\,
            I => \ppm_encoder_1.N_614_i\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__19934\,
            I => \N__19929\
        );

    \I__4132\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19926\
        );

    \I__4131\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19922\
        );

    \I__4130\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19919\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__19926\,
            I => \N__19916\
        );

    \I__4128\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19913\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__19922\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__19919\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__19916\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__19913\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__4123\ : InMux
    port map (
            O => \N__19904\,
            I => \ppm_encoder_1.un1_counter_13_cry_0\
        );

    \I__4122\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19895\
        );

    \I__4121\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19890\
        );

    \I__4120\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19890\
        );

    \I__4119\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19887\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__19895\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__19890\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__19887\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4115\ : InMux
    port map (
            O => \N__19880\,
            I => \ppm_encoder_1.un1_counter_13_cry_1\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__4113\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19870\
        );

    \I__4112\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19867\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19864\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__19867\,
            I => \N__19861\
        );

    \I__4109\ : Span12Mux_s10_v
    port map (
            O => \N__19864\,
            I => \N__19858\
        );

    \I__4108\ : Span12Mux_v
    port map (
            O => \N__19861\,
            I => \N__19855\
        );

    \I__4107\ : Odrv12
    port map (
            O => \N__19858\,
            I => scaler_2_data_12
        );

    \I__4106\ : Odrv12
    port map (
            O => \N__19855\,
            I => scaler_2_data_12
        );

    \I__4105\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__4103\ : Span4Mux_h
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__19841\,
            I => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\
        );

    \I__4101\ : InMux
    port map (
            O => \N__19838\,
            I => \ppm_encoder_1.un1_aileron_cry_11\
        );

    \I__4100\ : InMux
    port map (
            O => \N__19835\,
            I => \ppm_encoder_1.un1_aileron_cry_12\
        );

    \I__4099\ : InMux
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__4095\ : Span4Mux_v
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__19817\,
            I => scaler_2_data_14
        );

    \I__4093\ : InMux
    port map (
            O => \N__19814\,
            I => \bfn_11_25_0_\
        );

    \I__4092\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__4089\ : Span4Mux_h
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__4088\ : Odrv4
    port map (
            O => \N__19799\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\
        );

    \I__4087\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__4085\ : Span4Mux_v
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__19787\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\
        );

    \I__4083\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__19778\,
            I => \ppm_encoder_1.pulses2countZ0Z_4\
        );

    \I__4080\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4078\ : Span4Mux_h
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__19766\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__4075\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__4073\ : Span4Mux_s3_v
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__19751\,
            I => \ppm_encoder_1.pulses2countZ0Z_5\
        );

    \I__4071\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__19745\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__4068\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__19736\,
            I => \ppm_encoder_1.pulses2countZ0Z_13\
        );

    \I__4066\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__19730\,
            I => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\
        );

    \I__4064\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__19724\,
            I => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\
        );

    \I__4062\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__4060\ : Span4Mux_h
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__19709\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_5\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \N__19696\
        );

    \I__4056\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19687\
        );

    \I__4055\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19687\
        );

    \I__4054\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19684\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__19702\,
            I => \N__19681\
        );

    \I__4052\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19678\
        );

    \I__4051\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19673\
        );

    \I__4050\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19673\
        );

    \I__4049\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19663\
        );

    \I__4048\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19658\
        );

    \I__4047\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19658\
        );

    \I__4046\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19653\
        );

    \I__4045\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19653\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19648\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19648\
        );

    \I__4042\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19645\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__19678\,
            I => \N__19642\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__19673\,
            I => \N__19639\
        );

    \I__4039\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19634\
        );

    \I__4038\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19634\
        );

    \I__4037\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19629\
        );

    \I__4036\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19629\
        );

    \I__4035\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19622\
        );

    \I__4034\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19622\
        );

    \I__4033\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19622\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__19663\,
            I => \N__19613\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19613\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__19653\,
            I => \N__19613\
        );

    \I__4029\ : Span4Mux_h
    port map (
            O => \N__19648\,
            I => \N__19613\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__19645\,
            I => \N__19606\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__19642\,
            I => \N__19606\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__19639\,
            I => \N__19606\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__19634\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__19629\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__19622\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__19613\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__19606\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__4020\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__4018\ : Span4Mux_h
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__19586\,
            I => \ppm_encoder_1.un1_init_pulses_11_7\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__19583\,
            I => \N__19577\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__19582\,
            I => \N__19572\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__19581\,
            I => \N__19569\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__19580\,
            I => \N__19563\
        );

    \I__4012\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19558\
        );

    \I__4011\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19553\
        );

    \I__4010\ : InMux
    port map (
            O => \N__19575\,
            I => \N__19553\
        );

    \I__4009\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19544\
        );

    \I__4008\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19544\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \N__19541\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__19567\,
            I => \N__19538\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__19566\,
            I => \N__19535\
        );

    \I__4004\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19532\
        );

    \I__4003\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19527\
        );

    \I__4002\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19527\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19522\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19522\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__19552\,
            I => \N__19519\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__19551\,
            I => \N__19516\
        );

    \I__3997\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19512\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__19549\,
            I => \N__19509\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19506\
        );

    \I__3994\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19501\
        );

    \I__3993\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19501\
        );

    \I__3992\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19498\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__19532\,
            I => \N__19491\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__19527\,
            I => \N__19491\
        );

    \I__3989\ : Span4Mux_v
    port map (
            O => \N__19522\,
            I => \N__19488\
        );

    \I__3988\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19483\
        );

    \I__3987\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19483\
        );

    \I__3986\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19480\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__19512\,
            I => \N__19477\
        );

    \I__3984\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19474\
        );

    \I__3983\ : Span4Mux_v
    port map (
            O => \N__19506\,
            I => \N__19470\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__19501\,
            I => \N__19465\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__19498\,
            I => \N__19465\
        );

    \I__3980\ : InMux
    port map (
            O => \N__19497\,
            I => \N__19460\
        );

    \I__3979\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19460\
        );

    \I__3978\ : Span4Mux_v
    port map (
            O => \N__19491\,
            I => \N__19451\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__19488\,
            I => \N__19451\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19451\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__19480\,
            I => \N__19451\
        );

    \I__3974\ : Span4Mux_h
    port map (
            O => \N__19477\,
            I => \N__19446\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19446\
        );

    \I__3972\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19443\
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__19470\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3970\ : Odrv12
    port map (
            O => \N__19465\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__19460\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__19451\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__19446\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__19443\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3965\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__3963\ : Span4Mux_h
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__19421\,
            I => \ppm_encoder_1.un1_init_pulses_10_7\
        );

    \I__3961\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19412\
        );

    \I__3960\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19412\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__19412\,
            I => \N__19408\
        );

    \I__3958\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19405\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__19405\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__19402\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__3954\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19393\
        );

    \I__3953\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19390\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__19393\,
            I => \N__19387\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__19390\,
            I => \N__19384\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__19387\,
            I => \N__19381\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__19384\,
            I => \N__19378\
        );

    \I__3948\ : Span4Mux_v
    port map (
            O => \N__19381\,
            I => \N__19375\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__3946\ : Span4Mux_v
    port map (
            O => \N__19375\,
            I => \N__19369\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__19372\,
            I => scaler_2_data_6
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__19369\,
            I => scaler_2_data_6
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__3942\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19357\
        );

    \I__3941\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__19357\,
            I => \N__19351\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__19354\,
            I => \N__19348\
        );

    \I__3938\ : Span4Mux_v
    port map (
            O => \N__19351\,
            I => \N__19343\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__19348\,
            I => \N__19343\
        );

    \I__3936\ : Span4Mux_v
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__19340\,
            I => scaler_2_data_7
        );

    \I__3934\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__19331\,
            I => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\
        );

    \I__3931\ : InMux
    port map (
            O => \N__19328\,
            I => \ppm_encoder_1.un1_aileron_cry_6\
        );

    \I__3930\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19321\
        );

    \I__3929\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19318\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__19321\,
            I => \N__19315\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__19318\,
            I => \N__19312\
        );

    \I__3926\ : Sp12to4
    port map (
            O => \N__19315\,
            I => \N__19307\
        );

    \I__3925\ : Span12Mux_h
    port map (
            O => \N__19312\,
            I => \N__19307\
        );

    \I__3924\ : Odrv12
    port map (
            O => \N__19307\,
            I => scaler_2_data_8
        );

    \I__3923\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__3921\ : Span4Mux_h
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__19292\,
            I => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\
        );

    \I__3918\ : InMux
    port map (
            O => \N__19289\,
            I => \ppm_encoder_1.un1_aileron_cry_7\
        );

    \I__3917\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19282\
        );

    \I__3916\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19279\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__19282\,
            I => \N__19276\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__19279\,
            I => \N__19271\
        );

    \I__3913\ : Span4Mux_v
    port map (
            O => \N__19276\,
            I => \N__19271\
        );

    \I__3912\ : Span4Mux_v
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__19268\,
            I => scaler_2_data_9
        );

    \I__3910\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__19256\,
            I => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\
        );

    \I__3906\ : InMux
    port map (
            O => \N__19253\,
            I => \ppm_encoder_1.un1_aileron_cry_8\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__3904\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19243\
        );

    \I__3903\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19240\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__19243\,
            I => \N__19235\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__19240\,
            I => \N__19235\
        );

    \I__3900\ : Span4Mux_v
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__3899\ : Span4Mux_v
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__19229\,
            I => scaler_2_data_10
        );

    \I__3897\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__19223\,
            I => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\
        );

    \I__3895\ : InMux
    port map (
            O => \N__19220\,
            I => \ppm_encoder_1.un1_aileron_cry_9\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__3893\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19210\
        );

    \I__3892\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19207\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__19210\,
            I => \N__19204\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19201\
        );

    \I__3889\ : Span4Mux_h
    port map (
            O => \N__19204\,
            I => \N__19196\
        );

    \I__3888\ : Span4Mux_v
    port map (
            O => \N__19201\,
            I => \N__19196\
        );

    \I__3887\ : Span4Mux_v
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__19193\,
            I => scaler_2_data_11
        );

    \I__3885\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__19181\,
            I => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\
        );

    \I__3881\ : InMux
    port map (
            O => \N__19178\,
            I => \ppm_encoder_1.un1_aileron_cry_10\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__19175\,
            I => \N__19171\
        );

    \I__3879\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19168\
        );

    \I__3878\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19165\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__19168\,
            I => \N__19162\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__19165\,
            I => \N__19159\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__19162\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__19159\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__3873\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__3871\ : Span4Mux_h
    port map (
            O => \N__19148\,
            I => \N__19143\
        );

    \I__3870\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19138\
        );

    \I__3869\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19138\
        );

    \I__3868\ : Odrv4
    port map (
            O => \N__19143\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__19138\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__3866\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19128\
        );

    \I__3865\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19125\
        );

    \I__3864\ : InMux
    port map (
            O => \N__19131\,
            I => \N__19122\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__19128\,
            I => \N__19119\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__19125\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__19122\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__19119\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__3859\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__19103\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__3854\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__19094\,
            I => \N__19089\
        );

    \I__3852\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19084\
        );

    \I__3851\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19084\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__19089\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__19084\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__3848\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__3846\ : Span12Mux_v
    port map (
            O => \N__19073\,
            I => \N__19068\
        );

    \I__3845\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19063\
        );

    \I__3844\ : InMux
    port map (
            O => \N__19071\,
            I => \N__19063\
        );

    \I__3843\ : Odrv12
    port map (
            O => \N__19068\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__19063\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__3841\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__19055\,
            I => \N__19051\
        );

    \I__3839\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19048\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__19051\,
            I => \N__19043\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__19048\,
            I => \N__19043\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__19040\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__19037\,
            I => \N__19033\
        );

    \I__3833\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19029\
        );

    \I__3832\ : InMux
    port map (
            O => \N__19033\,
            I => \N__19026\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__19032\,
            I => \N__19023\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__19029\,
            I => \N__19020\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__19026\,
            I => \N__19017\
        );

    \I__3828\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19014\
        );

    \I__3827\ : Span4Mux_v
    port map (
            O => \N__19020\,
            I => \N__19011\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__19017\,
            I => \N__19008\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__19014\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__19011\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__19008\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__3821\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__3819\ : Span4Mux_h
    port map (
            O => \N__18992\,
            I => \N__18989\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__18989\,
            I => \N__18984\
        );

    \I__3817\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18979\
        );

    \I__3816\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18979\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__18984\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__18979\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__3813\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__18971\,
            I => \N__18968\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__18968\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\
        );

    \I__3810\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__18956\,
            I => \ppm_encoder_1.un1_init_pulses_11_3\
        );

    \I__3806\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__3804\ : Span4Mux_h
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__18944\,
            I => \ppm_encoder_1.un1_init_pulses_10_3\
        );

    \I__3802\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18938\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__18932\,
            I => \ppm_encoder_1.un1_init_pulses_11_5\
        );

    \I__3798\ : InMux
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__18926\,
            I => \N__18923\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__18920\,
            I => \ppm_encoder_1.un1_init_pulses_10_5\
        );

    \I__3794\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18913\
        );

    \I__3793\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18910\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__18913\,
            I => \N__18907\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__18910\,
            I => \N__18904\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__18907\,
            I => \N__18901\
        );

    \I__3789\ : Odrv12
    port map (
            O => \N__18904\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__18901\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__3787\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__18893\,
            I => \N__18889\
        );

    \I__3785\ : InMux
    port map (
            O => \N__18892\,
            I => \N__18886\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__18889\,
            I => \N__18883\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__18886\,
            I => \N__18880\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__18883\,
            I => scaler_3_data_12
        );

    \I__3781\ : Odrv12
    port map (
            O => \N__18880\,
            I => scaler_3_data_12
        );

    \I__3780\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__18869\,
            I => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\
        );

    \I__3777\ : InMux
    port map (
            O => \N__18866\,
            I => \ppm_encoder_1.un1_elevator_cry_11\
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__3775\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__18857\,
            I => \N__18853\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__3772\ : Sp12to4
    port map (
            O => \N__18853\,
            I => \N__18847\
        );

    \I__3771\ : InMux
    port map (
            O => \N__18850\,
            I => \N__18844\
        );

    \I__3770\ : Span12Mux_s6_v
    port map (
            O => \N__18847\,
            I => \N__18839\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__18844\,
            I => \N__18839\
        );

    \I__3768\ : Odrv12
    port map (
            O => \N__18839\,
            I => scaler_3_data_13
        );

    \I__3767\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__3765\ : Sp12to4
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__3764\ : Odrv12
    port map (
            O => \N__18827\,
            I => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\
        );

    \I__3763\ : InMux
    port map (
            O => \N__18824\,
            I => \ppm_encoder_1.un1_elevator_cry_12\
        );

    \I__3762\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__18812\,
            I => scaler_3_data_14
        );

    \I__3758\ : InMux
    port map (
            O => \N__18809\,
            I => \bfn_11_20_0_\
        );

    \I__3757\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__3755\ : Odrv12
    port map (
            O => \N__18800\,
            I => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__3753\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__3751\ : Odrv12
    port map (
            O => \N__18788\,
            I => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__3749\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18777\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__18781\,
            I => \N__18774\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__18780\,
            I => \N__18770\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18762\
        );

    \I__3745\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18759\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__18773\,
            I => \N__18756\
        );

    \I__3743\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18753\
        );

    \I__3742\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18750\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__18768\,
            I => \N__18747\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__18767\,
            I => \N__18743\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__18766\,
            I => \N__18740\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__18765\,
            I => \N__18737\
        );

    \I__3737\ : Span4Mux_h
    port map (
            O => \N__18762\,
            I => \N__18732\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__18759\,
            I => \N__18732\
        );

    \I__3735\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18729\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__18753\,
            I => \N__18726\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18723\
        );

    \I__3732\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18718\
        );

    \I__3731\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18718\
        );

    \I__3730\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18715\
        );

    \I__3729\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18712\
        );

    \I__3728\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18709\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__18732\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__18729\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__18726\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__18723\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__18718\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__18715\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__18712\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__18709\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__3719\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18684\
        );

    \I__3718\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18681\
        );

    \I__3717\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18678\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__18689\,
            I => \N__18675\
        );

    \I__3715\ : InMux
    port map (
            O => \N__18688\,
            I => \N__18669\
        );

    \I__3714\ : InMux
    port map (
            O => \N__18687\,
            I => \N__18666\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__18684\,
            I => \N__18660\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__18681\,
            I => \N__18660\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__18678\,
            I => \N__18657\
        );

    \I__3710\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18653\
        );

    \I__3709\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18648\
        );

    \I__3708\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18648\
        );

    \I__3707\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18645\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__18669\,
            I => \N__18638\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__18666\,
            I => \N__18638\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__18665\,
            I => \N__18634\
        );

    \I__3703\ : Span4Mux_v
    port map (
            O => \N__18660\,
            I => \N__18631\
        );

    \I__3702\ : Span4Mux_h
    port map (
            O => \N__18657\,
            I => \N__18628\
        );

    \I__3701\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18625\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__18653\,
            I => \N__18620\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__18648\,
            I => \N__18620\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__18645\,
            I => \N__18617\
        );

    \I__3697\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18614\
        );

    \I__3696\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18611\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__18638\,
            I => \N__18608\
        );

    \I__3694\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18603\
        );

    \I__3693\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18603\
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__18631\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__18628\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__18625\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__18620\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__18617\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__18614\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__18611\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__18608\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__18603\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3683\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__18581\,
            I => \N__18578\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__18578\,
            I => \N__18574\
        );

    \I__3680\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18571\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__18574\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__18571\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__18566\,
            I => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__3675\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__3673\ : Span4Mux_v
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__18551\,
            I => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__3670\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18540\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__18544\,
            I => \N__18537\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__18543\,
            I => \N__18532\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18527\
        );

    \I__3666\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18524\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__18536\,
            I => \N__18521\
        );

    \I__3664\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18518\
        );

    \I__3663\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18514\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__18531\,
            I => \N__18509\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__18530\,
            I => \N__18506\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__18527\,
            I => \N__18500\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__18524\,
            I => \N__18500\
        );

    \I__3658\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18497\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__18518\,
            I => \N__18494\
        );

    \I__3656\ : InMux
    port map (
            O => \N__18517\,
            I => \N__18491\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__18514\,
            I => \N__18488\
        );

    \I__3654\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18483\
        );

    \I__3653\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18483\
        );

    \I__3652\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18480\
        );

    \I__3651\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18477\
        );

    \I__3650\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18474\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__18500\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__18497\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__18494\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__18491\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__18488\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__18483\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__18480\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__18477\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__18474\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3640\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18448\
        );

    \I__3639\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18445\
        );

    \I__3638\ : InMux
    port map (
            O => \N__18453\,
            I => \N__18441\
        );

    \I__3637\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18437\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__18451\,
            I => \N__18432\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__18448\,
            I => \N__18424\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__18445\,
            I => \N__18424\
        );

    \I__3633\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18421\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__18441\,
            I => \N__18418\
        );

    \I__3631\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18415\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__18437\,
            I => \N__18412\
        );

    \I__3629\ : InMux
    port map (
            O => \N__18436\,
            I => \N__18409\
        );

    \I__3628\ : InMux
    port map (
            O => \N__18435\,
            I => \N__18404\
        );

    \I__3627\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18404\
        );

    \I__3626\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18401\
        );

    \I__3625\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18398\
        );

    \I__3624\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18395\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__18424\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__18421\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__18418\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__18415\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3619\ : Odrv4
    port map (
            O => \N__18412\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__18409\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__18404\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__18401\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__18398\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__18395\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3613\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__18371\,
            I => \ppm_encoder_1.un2_throttle_iv_1_14\
        );

    \I__3611\ : InMux
    port map (
            O => \N__18368\,
            I => \ppm_encoder_1.un1_rudder_cry_12\
        );

    \I__3610\ : InMux
    port map (
            O => \N__18365\,
            I => \bfn_11_18_0_\
        );

    \I__3609\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__18359\,
            I => \N__18355\
        );

    \I__3607\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18352\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__18355\,
            I => \N__18347\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18347\
        );

    \I__3604\ : Span4Mux_v
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__18344\,
            I => scaler_3_data_6
        );

    \I__3602\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__18338\,
            I => \N__18334\
        );

    \I__3600\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18331\
        );

    \I__3599\ : Span4Mux_v
    port map (
            O => \N__18334\,
            I => \N__18328\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__18331\,
            I => \N__18325\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__18328\,
            I => scaler_3_data_7
        );

    \I__3596\ : Odrv12
    port map (
            O => \N__18325\,
            I => scaler_3_data_7
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__18320\,
            I => \N__18317\
        );

    \I__3594\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18314\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__3592\ : Span4Mux_v
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__18308\,
            I => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\
        );

    \I__3590\ : InMux
    port map (
            O => \N__18305\,
            I => \ppm_encoder_1.un1_elevator_cry_6\
        );

    \I__3589\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18298\
        );

    \I__3588\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18295\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__18298\,
            I => \N__18290\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__18295\,
            I => \N__18290\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__18287\,
            I => scaler_3_data_8
        );

    \I__3583\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__18281\,
            I => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\
        );

    \I__3581\ : InMux
    port map (
            O => \N__18278\,
            I => \ppm_encoder_1.un1_elevator_cry_7\
        );

    \I__3580\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__3578\ : Span4Mux_h
    port map (
            O => \N__18269\,
            I => \N__18265\
        );

    \I__3577\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18262\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__18265\,
            I => \N__18259\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__18262\,
            I => \N__18256\
        );

    \I__3574\ : Odrv4
    port map (
            O => \N__18259\,
            I => scaler_3_data_9
        );

    \I__3573\ : Odrv12
    port map (
            O => \N__18256\,
            I => scaler_3_data_9
        );

    \I__3572\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__18248\,
            I => \N__18245\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__18242\,
            I => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\
        );

    \I__3568\ : InMux
    port map (
            O => \N__18239\,
            I => \ppm_encoder_1.un1_elevator_cry_8\
        );

    \I__3567\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__18230\,
            I => \N__18226\
        );

    \I__3564\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18223\
        );

    \I__3563\ : Span4Mux_v
    port map (
            O => \N__18226\,
            I => \N__18220\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__18223\,
            I => \N__18217\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__18220\,
            I => scaler_3_data_10
        );

    \I__3560\ : Odrv12
    port map (
            O => \N__18217\,
            I => scaler_3_data_10
        );

    \I__3559\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__3557\ : Span4Mux_v
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__18203\,
            I => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\
        );

    \I__3555\ : InMux
    port map (
            O => \N__18200\,
            I => \ppm_encoder_1.un1_elevator_cry_9\
        );

    \I__3554\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18193\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__18196\,
            I => \N__18190\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__18193\,
            I => \N__18187\
        );

    \I__3551\ : InMux
    port map (
            O => \N__18190\,
            I => \N__18184\
        );

    \I__3550\ : Sp12to4
    port map (
            O => \N__18187\,
            I => \N__18179\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__18184\,
            I => \N__18179\
        );

    \I__3548\ : Odrv12
    port map (
            O => \N__18179\,
            I => scaler_3_data_11
        );

    \I__3547\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__18173\,
            I => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\
        );

    \I__3545\ : InMux
    port map (
            O => \N__18170\,
            I => \ppm_encoder_1.un1_elevator_cry_10\
        );

    \I__3544\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18163\
        );

    \I__3543\ : InMux
    port map (
            O => \N__18166\,
            I => \N__18160\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__18163\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__18160\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__3539\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__18149\,
            I => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\
        );

    \I__3537\ : InMux
    port map (
            O => \N__18146\,
            I => \bfn_11_16_0_\
        );

    \I__3536\ : InMux
    port map (
            O => \N__18143\,
            I => \scaler_3.un2_source_data_0_cry_9\
        );

    \I__3535\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18137\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__18137\,
            I => \N__18134\
        );

    \I__3533\ : Span4Mux_v
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__18131\,
            I => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\
        );

    \I__3531\ : InMux
    port map (
            O => \N__18128\,
            I => \ppm_encoder_1.un1_rudder_cry_6\
        );

    \I__3530\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__18119\,
            I => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\
        );

    \I__3527\ : InMux
    port map (
            O => \N__18116\,
            I => \ppm_encoder_1.un1_rudder_cry_7\
        );

    \I__3526\ : InMux
    port map (
            O => \N__18113\,
            I => \ppm_encoder_1.un1_rudder_cry_8\
        );

    \I__3525\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__3522\ : Odrv4
    port map (
            O => \N__18101\,
            I => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\
        );

    \I__3521\ : InMux
    port map (
            O => \N__18098\,
            I => \ppm_encoder_1.un1_rudder_cry_9\
        );

    \I__3520\ : InMux
    port map (
            O => \N__18095\,
            I => \ppm_encoder_1.un1_rudder_cry_10\
        );

    \I__3519\ : InMux
    port map (
            O => \N__18092\,
            I => \ppm_encoder_1.un1_rudder_cry_11\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__3517\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18083\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__3515\ : Span4Mux_h
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__18077\,
            I => \scaler_3.un2_source_data_0_cry_1_c_RNO_1\
        );

    \I__3513\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18070\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__18073\,
            I => \N__18066\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__18070\,
            I => \N__18062\
        );

    \I__3510\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18059\
        );

    \I__3509\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18054\
        );

    \I__3508\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18054\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__18062\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__18059\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__18054\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__3504\ : InMux
    port map (
            O => \N__18047\,
            I => \scaler_3.un2_source_data_0_cry_1\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__3502\ : InMux
    port map (
            O => \N__18041\,
            I => \N__18035\
        );

    \I__3501\ : InMux
    port map (
            O => \N__18040\,
            I => \N__18035\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__18035\,
            I => \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I\
        );

    \I__3499\ : InMux
    port map (
            O => \N__18032\,
            I => \scaler_3.un2_source_data_0_cry_2\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__18029\,
            I => \N__18026\
        );

    \I__3497\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18020\
        );

    \I__3496\ : InMux
    port map (
            O => \N__18025\,
            I => \N__18020\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__18020\,
            I => \scaler_3.un3_source_data_0_cry_2_c_RNIR08I\
        );

    \I__3494\ : InMux
    port map (
            O => \N__18017\,
            I => \scaler_3.un2_source_data_0_cry_3\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__3492\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18005\
        );

    \I__3491\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18005\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__18005\,
            I => \scaler_3.un3_source_data_0_cry_3_c_RNIU49I\
        );

    \I__3489\ : InMux
    port map (
            O => \N__18002\,
            I => \scaler_3.un2_source_data_0_cry_4\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__3487\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17990\
        );

    \I__3486\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17990\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__17990\,
            I => \scaler_3.un3_source_data_0_cry_4_c_RNI19AI\
        );

    \I__3484\ : InMux
    port map (
            O => \N__17987\,
            I => \scaler_3.un2_source_data_0_cry_5\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__3482\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17975\
        );

    \I__3481\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17975\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__17975\,
            I => \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI\
        );

    \I__3479\ : InMux
    port map (
            O => \N__17972\,
            I => \scaler_3.un2_source_data_0_cry_6\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__3477\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17960\
        );

    \I__3476\ : InMux
    port map (
            O => \N__17965\,
            I => \N__17960\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__17960\,
            I => \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI\
        );

    \I__3474\ : InMux
    port map (
            O => \N__17957\,
            I => \scaler_3.un2_source_data_0_cry_7\
        );

    \I__3473\ : InMux
    port map (
            O => \N__17954\,
            I => \bfn_11_13_0_\
        );

    \I__3472\ : InMux
    port map (
            O => \N__17951\,
            I => \scaler_4.un3_source_data_0_cry_8\
        );

    \I__3471\ : CEMux
    port map (
            O => \N__17948\,
            I => \N__17945\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__3469\ : Sp12to4
    port map (
            O => \N__17942\,
            I => \N__17939\
        );

    \I__3468\ : Odrv12
    port map (
            O => \N__17939\,
            I => \uart_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__3467\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17932\
        );

    \I__3466\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17929\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__17932\,
            I => \N__17926\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__17929\,
            I => \N__17922\
        );

    \I__3463\ : Span4Mux_h
    port map (
            O => \N__17926\,
            I => \N__17919\
        );

    \I__3462\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17916\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__17922\,
            I => \N__17908\
        );

    \I__3460\ : Span4Mux_v
    port map (
            O => \N__17919\,
            I => \N__17908\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__17916\,
            I => \N__17908\
        );

    \I__3458\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17905\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__17908\,
            I => \frame_decoder_CH4data_0\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__17905\,
            I => \frame_decoder_CH4data_0\
        );

    \I__3455\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17892\
        );

    \I__3453\ : InMux
    port map (
            O => \N__17896\,
            I => \N__17889\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__17895\,
            I => \N__17885\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__17892\,
            I => \N__17880\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__17889\,
            I => \N__17880\
        );

    \I__3449\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17877\
        );

    \I__3448\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17874\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__17880\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__17877\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__17874\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__3444\ : InMux
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__17864\,
            I => \scaler_4.N_544_i_l_ofxZ0\
        );

    \I__3442\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17857\
        );

    \I__3441\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17854\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__17857\,
            I => \N__17851\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__17854\,
            I => \frame_decoder_OFF2data_7\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__17851\,
            I => \frame_decoder_OFF2data_7\
        );

    \I__3437\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__17843\,
            I => \N__17840\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__17840\,
            I => \scaler_2.un3_source_data_0_axb_7\
        );

    \I__3434\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__17831\,
            I => \N__17827\
        );

    \I__3431\ : InMux
    port map (
            O => \N__17830\,
            I => \N__17824\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__17827\,
            I => \frame_decoder_CH2data_7\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__17824\,
            I => \frame_decoder_CH2data_7\
        );

    \I__3428\ : CEMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17812\
        );

    \I__3426\ : CEMux
    port map (
            O => \N__17815\,
            I => \N__17809\
        );

    \I__3425\ : Span4Mux_h
    port map (
            O => \N__17812\,
            I => \N__17806\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__17809\,
            I => \N__17803\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__17806\,
            I => \uart_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__3422\ : Odrv12
    port map (
            O => \N__17803\,
            I => \uart_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__3421\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17795\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17791\
        );

    \I__3419\ : InMux
    port map (
            O => \N__17794\,
            I => \N__17788\
        );

    \I__3418\ : Span4Mux_h
    port map (
            O => \N__17791\,
            I => \N__17785\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__17788\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__17785\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__3415\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__17777\,
            I => \N__17774\
        );

    \I__3413\ : Span4Mux_v
    port map (
            O => \N__17774\,
            I => \N__17770\
        );

    \I__3412\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17767\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__17770\,
            I => \uart_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__17767\,
            I => \uart_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__3409\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17758\
        );

    \I__3408\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17755\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17752\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__17755\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__17752\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__3404\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17743\
        );

    \I__3403\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17740\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__17743\,
            I => \N__17735\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__17740\,
            I => \N__17735\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__17735\,
            I => \frame_decoder_CH4data_7\
        );

    \I__3399\ : InMux
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__17726\,
            I => \scaler_4.un3_source_data_0_axb_7\
        );

    \I__3396\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17720\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__17720\,
            I => \frame_decoder_CH4data_1\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__3393\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17711\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__17711\,
            I => \frame_decoder_OFF4data_1\
        );

    \I__3391\ : InMux
    port map (
            O => \N__17708\,
            I => \scaler_4.un3_source_data_0_cry_0\
        );

    \I__3390\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17702\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__17702\,
            I => \frame_decoder_CH4data_2\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__3387\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__17693\,
            I => \frame_decoder_OFF4data_2\
        );

    \I__3385\ : InMux
    port map (
            O => \N__17690\,
            I => \scaler_4.un3_source_data_0_cry_1\
        );

    \I__3384\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__17684\,
            I => \frame_decoder_CH4data_3\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__17681\,
            I => \N__17678\
        );

    \I__3381\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__17675\,
            I => \frame_decoder_OFF4data_3\
        );

    \I__3379\ : InMux
    port map (
            O => \N__17672\,
            I => \scaler_4.un3_source_data_0_cry_2\
        );

    \I__3378\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17666\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__17666\,
            I => \frame_decoder_CH4data_4\
        );

    \I__3376\ : InMux
    port map (
            O => \N__17663\,
            I => \scaler_4.un3_source_data_0_cry_3\
        );

    \I__3375\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__17657\,
            I => \frame_decoder_CH4data_5\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__17654\,
            I => \N__17651\
        );

    \I__3372\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17648\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__17648\,
            I => \frame_decoder_OFF4data_5\
        );

    \I__3370\ : InMux
    port map (
            O => \N__17645\,
            I => \scaler_4.un3_source_data_0_cry_4\
        );

    \I__3369\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17639\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__17639\,
            I => \frame_decoder_CH4data_6\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__17636\,
            I => \N__17633\
        );

    \I__3366\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17630\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__17630\,
            I => \frame_decoder_OFF4data_6\
        );

    \I__3364\ : InMux
    port map (
            O => \N__17627\,
            I => \scaler_4.un3_source_data_0_cry_5\
        );

    \I__3363\ : InMux
    port map (
            O => \N__17624\,
            I => \scaler_4.un3_source_data_0_cry_6\
        );

    \I__3362\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__17618\,
            I => \ppm_encoder_1.pulses2countZ0Z_10\
        );

    \I__3360\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17612\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__3358\ : Odrv4
    port map (
            O => \N__17609\,
            I => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\
        );

    \I__3357\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__17603\,
            I => \N__17600\
        );

    \I__3355\ : Span4Mux_s3_v
    port map (
            O => \N__17600\,
            I => \N__17597\
        );

    \I__3354\ : Span4Mux_v
    port map (
            O => \N__17597\,
            I => \N__17594\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__17594\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__3351\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__17585\,
            I => \ppm_encoder_1.pulses2countZ0Z_11\
        );

    \I__3349\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__17579\,
            I => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\
        );

    \I__3347\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__17573\,
            I => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\
        );

    \I__3345\ : InMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__17567\,
            I => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\
        );

    \I__3343\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17560\
        );

    \I__3342\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17557\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__17560\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__17557\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__17552\,
            I => \N__17548\
        );

    \I__3338\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17545\
        );

    \I__3337\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17542\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__17545\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__17542\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__3334\ : InMux
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__17534\,
            I => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\
        );

    \I__3332\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17527\
        );

    \I__3331\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17524\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__17527\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__17524\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__3327\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__17513\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\
        );

    \I__3325\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17507\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__17507\,
            I => \N__17504\
        );

    \I__3323\ : Span4Mux_s2_v
    port map (
            O => \N__17504\,
            I => \N__17501\
        );

    \I__3322\ : Span4Mux_v
    port map (
            O => \N__17501\,
            I => \N__17498\
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__17498\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\
        );

    \I__3320\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__17492\,
            I => \ppm_encoder_1.pulses2countZ0Z_2\
        );

    \I__3318\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17486\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__17486\,
            I => \N__17483\
        );

    \I__3316\ : Span4Mux_s3_v
    port map (
            O => \N__17483\,
            I => \N__17480\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__17480\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\
        );

    \I__3314\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17474\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__17474\,
            I => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\
        );

    \I__3312\ : InMux
    port map (
            O => \N__17471\,
            I => \ppm_encoder_1.counter24_0_N_2\
        );

    \I__3311\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__3309\ : Span4Mux_s3_v
    port map (
            O => \N__17462\,
            I => \N__17459\
        );

    \I__3308\ : Span4Mux_v
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__17456\,
            I => \ppm_encoder_1.pulses2countZ0Z_8\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__3305\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17444\
        );

    \I__3303\ : Odrv12
    port map (
            O => \N__17444\,
            I => \ppm_encoder_1.pulses2countZ0Z_9\
        );

    \I__3302\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17438\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3300\ : Span4Mux_v
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__17432\,
            I => \ppm_encoder_1.un1_init_pulses_11_8\
        );

    \I__3298\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__17426\,
            I => \ppm_encoder_1.un1_init_pulses_10_8\
        );

    \I__3296\ : InMux
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__17420\,
            I => \N__17416\
        );

    \I__3294\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17413\
        );

    \I__3293\ : Sp12to4
    port map (
            O => \N__17416\,
            I => \N__17410\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__17413\,
            I => \N__17407\
        );

    \I__3291\ : Odrv12
    port map (
            O => \N__17410\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__17407\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__3289\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__17393\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_8\
        );

    \I__3285\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__3283\ : Span4Mux_v
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__17381\,
            I => \ppm_encoder_1.un1_init_pulses_11_9\
        );

    \I__3281\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17375\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__17375\,
            I => \ppm_encoder_1.un1_init_pulses_10_9\
        );

    \I__3279\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__17369\,
            I => \N__17366\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__17366\,
            I => \N__17362\
        );

    \I__3276\ : InMux
    port map (
            O => \N__17365\,
            I => \N__17359\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__17362\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__17359\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__3273\ : InMux
    port map (
            O => \N__17354\,
            I => \N__17351\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__17351\,
            I => \N__17348\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__17348\,
            I => \N__17345\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__17345\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_9\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__17342\,
            I => \ppm_encoder_1.N_305_cascade_\
        );

    \I__3268\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17330\
        );

    \I__3267\ : InMux
    port map (
            O => \N__17338\,
            I => \N__17330\
        );

    \I__3266\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17330\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__17330\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__3264\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17318\
        );

    \I__3263\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17318\
        );

    \I__3262\ : InMux
    port map (
            O => \N__17325\,
            I => \N__17318\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__17318\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__3260\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17311\
        );

    \I__3259\ : InMux
    port map (
            O => \N__17314\,
            I => \N__17308\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__17311\,
            I => \N__17303\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__17308\,
            I => \N__17303\
        );

    \I__3256\ : Odrv12
    port map (
            O => \N__17303\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__17300\,
            I => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \N__17294\
        );

    \I__3253\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17291\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__17291\,
            I => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\
        );

    \I__3251\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17285\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__17285\,
            I => \ppm_encoder_1.un2_throttle_iv_1_13\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__17282\,
            I => \ppm_encoder_1.N_308_cascade_\
        );

    \I__3248\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17270\
        );

    \I__3247\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17270\
        );

    \I__3246\ : InMux
    port map (
            O => \N__17277\,
            I => \N__17270\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__17270\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__3244\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17258\
        );

    \I__3243\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17258\
        );

    \I__3242\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17258\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__17258\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__3240\ : InMux
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__17252\,
            I => \ppm_encoder_1.un2_throttle_iv_1_6\
        );

    \I__3238\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17240\
        );

    \I__3237\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17240\
        );

    \I__3236\ : InMux
    port map (
            O => \N__17247\,
            I => \N__17240\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__17240\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__3234\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17228\
        );

    \I__3233\ : InMux
    port map (
            O => \N__17236\,
            I => \N__17228\
        );

    \I__3232\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17228\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__17228\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__3230\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__17222\,
            I => \N__17218\
        );

    \I__3228\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17215\
        );

    \I__3227\ : Span4Mux_h
    port map (
            O => \N__17218\,
            I => \N__17210\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__17215\,
            I => \N__17210\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__17210\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__17207\,
            I => \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__17204\,
            I => \N__17201\
        );

    \I__3222\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__17198\,
            I => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\
        );

    \I__3220\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__17192\,
            I => \ppm_encoder_1.un2_throttle_iv_1_10\
        );

    \I__3218\ : InMux
    port map (
            O => \N__17189\,
            I => \N__17185\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__17188\,
            I => \N__17182\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__17185\,
            I => \N__17179\
        );

    \I__3215\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__17179\,
            I => \N__17171\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__17176\,
            I => \N__17171\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__17171\,
            I => \N__17168\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__17168\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__17165\,
            I => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\
        );

    \I__3209\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17159\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__17159\,
            I => \N__17156\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__17156\,
            I => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\
        );

    \I__3206\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17150\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__17150\,
            I => \ppm_encoder_1.un2_throttle_iv_1_7\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__17147\,
            I => \N__17142\
        );

    \I__3203\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17137\
        );

    \I__3202\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17137\
        );

    \I__3201\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17134\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__17134\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__17131\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__3197\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17120\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__17120\,
            I => \ppm_encoder_1.N_302\
        );

    \I__3194\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17112\
        );

    \I__3193\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17107\
        );

    \I__3192\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17107\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__17112\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__17107\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__3189\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17099\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__17099\,
            I => \N__17094\
        );

    \I__3187\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17089\
        );

    \I__3186\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17089\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__17094\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__17089\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__3183\ : InMux
    port map (
            O => \N__17084\,
            I => \N__17080\
        );

    \I__3182\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__17080\,
            I => \N__17074\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__17077\,
            I => \N__17071\
        );

    \I__3179\ : Span4Mux_v
    port map (
            O => \N__17074\,
            I => \N__17068\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__17071\,
            I => \N__17065\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__17068\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__17065\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__3173\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__17051\,
            I => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__17048\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__3170\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__17039\,
            I => \N__17035\
        );

    \I__3167\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17032\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__17035\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__17032\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__17027\,
            I => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__3162\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__3160\ : Span4Mux_v
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__17012\,
            I => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\
        );

    \I__3158\ : InMux
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__17006\,
            I => \ppm_encoder_1.un2_throttle_iv_1_12\
        );

    \I__3156\ : InMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__17000\,
            I => \N__16997\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__16997\,
            I => \ppm_encoder_1.N_307\
        );

    \I__3153\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16985\
        );

    \I__3152\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16985\
        );

    \I__3151\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16985\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__16985\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__3149\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__16976\,
            I => \N__16971\
        );

    \I__3146\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16966\
        );

    \I__3145\ : InMux
    port map (
            O => \N__16974\,
            I => \N__16966\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__16971\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__16966\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__16961\,
            I => \N__16957\
        );

    \I__3141\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16954\
        );

    \I__3140\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16950\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__16954\,
            I => \N__16947\
        );

    \I__3138\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16944\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__16950\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__16947\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__16944\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__3134\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16930\
        );

    \I__3133\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16930\
        );

    \I__3132\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16927\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__16930\,
            I => \N__16924\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__16927\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__16924\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__3128\ : InMux
    port map (
            O => \N__16919\,
            I => \N__16914\
        );

    \I__3127\ : InMux
    port map (
            O => \N__16918\,
            I => \N__16909\
        );

    \I__3126\ : InMux
    port map (
            O => \N__16917\,
            I => \N__16909\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__16914\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__16909\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__16904\,
            I => \N__16900\
        );

    \I__3122\ : InMux
    port map (
            O => \N__16903\,
            I => \N__16896\
        );

    \I__3121\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16893\
        );

    \I__3120\ : InMux
    port map (
            O => \N__16899\,
            I => \N__16890\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__16896\,
            I => \N__16887\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__16893\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__16890\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__16887\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__16877\,
            I => \N__16873\
        );

    \I__3113\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16869\
        );

    \I__3112\ : InMux
    port map (
            O => \N__16873\,
            I => \N__16866\
        );

    \I__3111\ : InMux
    port map (
            O => \N__16872\,
            I => \N__16863\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__16869\,
            I => \N__16860\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__16866\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__16863\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__16860\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__16853\,
            I => \ppm_encoder_1.N_303_cascade_\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__16850\,
            I => \N__16846\
        );

    \I__3104\ : InMux
    port map (
            O => \N__16849\,
            I => \N__16842\
        );

    \I__3103\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16839\
        );

    \I__3102\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16836\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__16842\,
            I => \N__16833\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__16839\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__16836\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__16833\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__3096\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16817\
        );

    \I__3095\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16817\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__16817\,
            I => \N__16814\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__16814\,
            I => \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11\
        );

    \I__3092\ : InMux
    port map (
            O => \N__16811\,
            I => \scaler_1.un2_source_data_0_cry_3\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__3090\ : InMux
    port map (
            O => \N__16805\,
            I => \N__16799\
        );

    \I__3089\ : InMux
    port map (
            O => \N__16804\,
            I => \N__16799\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__16796\,
            I => \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11\
        );

    \I__3086\ : InMux
    port map (
            O => \N__16793\,
            I => \scaler_1.un2_source_data_0_cry_4\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__3084\ : InMux
    port map (
            O => \N__16787\,
            I => \N__16781\
        );

    \I__3083\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16781\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__3081\ : Odrv12
    port map (
            O => \N__16778\,
            I => \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11\
        );

    \I__3080\ : InMux
    port map (
            O => \N__16775\,
            I => \scaler_1.un2_source_data_0_cry_5\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__3078\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16763\
        );

    \I__3077\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16763\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__3075\ : Odrv12
    port map (
            O => \N__16760\,
            I => \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11\
        );

    \I__3074\ : InMux
    port map (
            O => \N__16757\,
            I => \scaler_1.un2_source_data_0_cry_6\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__3072\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16745\
        );

    \I__3071\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16745\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3069\ : Odrv12
    port map (
            O => \N__16742\,
            I => \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11\
        );

    \I__3068\ : InMux
    port map (
            O => \N__16739\,
            I => \scaler_1.un2_source_data_0_cry_7\
        );

    \I__3067\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16732\
        );

    \I__3066\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16729\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__16732\,
            I => \N__16724\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__16729\,
            I => \N__16724\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__16724\,
            I => \N__16721\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__16721\,
            I => \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__3060\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__16709\,
            I => \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F\
        );

    \I__3057\ : InMux
    port map (
            O => \N__16706\,
            I => \bfn_10_18_0_\
        );

    \I__3056\ : InMux
    port map (
            O => \N__16703\,
            I => \scaler_1.un2_source_data_0_cry_9\
        );

    \I__3055\ : InMux
    port map (
            O => \N__16700\,
            I => \bfn_10_16_0_\
        );

    \I__3054\ : InMux
    port map (
            O => \N__16697\,
            I => \scaler_3.un3_source_data_0_cry_8\
        );

    \I__3053\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16691\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__16691\,
            I => \N__16687\
        );

    \I__3051\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16684\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__16687\,
            I => \N__16681\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__16684\,
            I => \uart_frame_decoder.count8_0_i\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__16681\,
            I => \uart_frame_decoder.count8_0_i\
        );

    \I__3047\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3045\ : Span4Mux_h
    port map (
            O => \N__16670\,
            I => \N__16666\
        );

    \I__3044\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16663\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__16666\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__16663\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__3041\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__16655\,
            I => \scaler_3.N_532_i_l_ofxZ0\
        );

    \I__3039\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__16643\,
            I => \uart_frame_decoder.state_1_RNINMHJZ0Z_10\
        );

    \I__3035\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16637\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__16637\,
            I => \N__16632\
        );

    \I__3033\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16627\
        );

    \I__3032\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16627\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__16632\,
            I => \uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__16627\,
            I => \uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61\
        );

    \I__3029\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__16619\,
            I => \N__16615\
        );

    \I__3027\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16612\
        );

    \I__3026\ : Span4Mux_h
    port map (
            O => \N__16615\,
            I => \N__16607\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__16612\,
            I => \N__16604\
        );

    \I__3024\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16599\
        );

    \I__3023\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16599\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__16607\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__16604\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__16599\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__3019\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16588\
        );

    \I__3018\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16584\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__16588\,
            I => \N__16580\
        );

    \I__3016\ : InMux
    port map (
            O => \N__16587\,
            I => \N__16577\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__16584\,
            I => \N__16574\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16571\
        );

    \I__3013\ : Span4Mux_v
    port map (
            O => \N__16580\,
            I => \N__16564\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__16577\,
            I => \N__16564\
        );

    \I__3011\ : Span4Mux_v
    port map (
            O => \N__16574\,
            I => \N__16564\
        );

    \I__3010\ : InMux
    port map (
            O => \N__16571\,
            I => \N__16561\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__16564\,
            I => \frame_decoder_OFF1data_0\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__16561\,
            I => \frame_decoder_OFF1data_0\
        );

    \I__3007\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16551\
        );

    \I__3006\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16548\
        );

    \I__3005\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16545\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16542\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16537\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__16545\,
            I => \N__16537\
        );

    \I__3001\ : Span4Mux_v
    port map (
            O => \N__16542\,
            I => \N__16533\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__16537\,
            I => \N__16530\
        );

    \I__2999\ : InMux
    port map (
            O => \N__16536\,
            I => \N__16527\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__16533\,
            I => \frame_decoder_CH1data_0\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__16530\,
            I => \frame_decoder_CH1data_0\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__16527\,
            I => \frame_decoder_CH1data_0\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__2994\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__16514\,
            I => \scaler_1.un2_source_data_0_cry_1_c_RNOZ0\
        );

    \I__2992\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16507\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__16510\,
            I => \N__16504\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__16507\,
            I => \N__16499\
        );

    \I__2989\ : InMux
    port map (
            O => \N__16504\,
            I => \N__16494\
        );

    \I__2988\ : InMux
    port map (
            O => \N__16503\,
            I => \N__16494\
        );

    \I__2987\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16491\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__16499\,
            I => \N__16486\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16486\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__16491\,
            I => \scaler_1.un2_source_data_0\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__16486\,
            I => \scaler_1.un2_source_data_0\
        );

    \I__2982\ : InMux
    port map (
            O => \N__16481\,
            I => \scaler_1.un2_source_data_0_cry_1\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__2980\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16469\
        );

    \I__2979\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16469\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__16466\,
            I => \scaler_1.un3_source_data_0_cry_1_c_RNIISC11\
        );

    \I__2976\ : InMux
    port map (
            O => \N__16463\,
            I => \scaler_1.un2_source_data_0_cry_2\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__16460\,
            I => \N__16456\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__16459\,
            I => \N__16452\
        );

    \I__2973\ : InMux
    port map (
            O => \N__16456\,
            I => \N__16446\
        );

    \I__2972\ : InMux
    port map (
            O => \N__16455\,
            I => \N__16446\
        );

    \I__2971\ : InMux
    port map (
            O => \N__16452\,
            I => \N__16443\
        );

    \I__2970\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16440\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__16446\,
            I => \N__16437\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__16443\,
            I => \N__16434\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__16440\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__16437\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__16434\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__16427\,
            I => \N__16424\
        );

    \I__2963\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16421\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__16421\,
            I => \N__16418\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__16418\,
            I => \frame_decoder_OFF3data_1\
        );

    \I__2960\ : InMux
    port map (
            O => \N__16415\,
            I => \scaler_3.un3_source_data_0_cry_0\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__16412\,
            I => \N__16409\
        );

    \I__2958\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__16403\,
            I => \frame_decoder_OFF3data_2\
        );

    \I__2955\ : InMux
    port map (
            O => \N__16400\,
            I => \scaler_3.un3_source_data_0_cry_1\
        );

    \I__2954\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__16394\,
            I => \N__16391\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__16391\,
            I => \frame_decoder_OFF3data_3\
        );

    \I__2951\ : InMux
    port map (
            O => \N__16388\,
            I => \scaler_3.un3_source_data_0_cry_2\
        );

    \I__2950\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__16382\,
            I => \N__16379\
        );

    \I__2948\ : Odrv4
    port map (
            O => \N__16379\,
            I => \frame_decoder_OFF3data_4\
        );

    \I__2947\ : InMux
    port map (
            O => \N__16376\,
            I => \scaler_3.un3_source_data_0_cry_3\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__2945\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16367\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__16367\,
            I => \N__16364\
        );

    \I__2943\ : Span4Mux_h
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__16361\,
            I => \frame_decoder_OFF3data_5\
        );

    \I__2941\ : InMux
    port map (
            O => \N__16358\,
            I => \scaler_3.un3_source_data_0_cry_4\
        );

    \I__2940\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__16352\,
            I => \N__16349\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__16349\,
            I => \frame_decoder_OFF3data_6\
        );

    \I__2937\ : InMux
    port map (
            O => \N__16346\,
            I => \scaler_3.un3_source_data_0_cry_5\
        );

    \I__2936\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16340\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__16340\,
            I => \scaler_3.un3_source_data_0_axb_7\
        );

    \I__2934\ : InMux
    port map (
            O => \N__16337\,
            I => \scaler_3.un3_source_data_0_cry_6\
        );

    \I__2933\ : InMux
    port map (
            O => \N__16334\,
            I => \scaler_2.un2_source_data_0_cry_2\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__2931\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16322\
        );

    \I__2930\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16322\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__16322\,
            I => \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH\
        );

    \I__2928\ : InMux
    port map (
            O => \N__16319\,
            I => \scaler_2.un2_source_data_0_cry_3\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__16316\,
            I => \N__16313\
        );

    \I__2926\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16307\
        );

    \I__2925\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16307\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__16307\,
            I => \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH\
        );

    \I__2923\ : InMux
    port map (
            O => \N__16304\,
            I => \scaler_2.un2_source_data_0_cry_4\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__16301\,
            I => \N__16298\
        );

    \I__2921\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16292\
        );

    \I__2920\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16292\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__16292\,
            I => \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH\
        );

    \I__2918\ : InMux
    port map (
            O => \N__16289\,
            I => \scaler_2.un2_source_data_0_cry_5\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__16286\,
            I => \N__16283\
        );

    \I__2916\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16277\
        );

    \I__2915\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16277\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__16277\,
            I => \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH\
        );

    \I__2913\ : InMux
    port map (
            O => \N__16274\,
            I => \scaler_2.un2_source_data_0_cry_6\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__16271\,
            I => \N__16268\
        );

    \I__2911\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16262\
        );

    \I__2910\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16262\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__16262\,
            I => \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH\
        );

    \I__2908\ : InMux
    port map (
            O => \N__16259\,
            I => \scaler_2.un2_source_data_0_cry_7\
        );

    \I__2907\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16252\
        );

    \I__2906\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16249\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__16252\,
            I => \N__16246\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__16249\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__16246\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__16241\,
            I => \N__16238\
        );

    \I__2901\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16235\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__16235\,
            I => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\
        );

    \I__2899\ : InMux
    port map (
            O => \N__16232\,
            I => \bfn_10_14_0_\
        );

    \I__2898\ : InMux
    port map (
            O => \N__16229\,
            I => \scaler_2.un2_source_data_0_cry_9\
        );

    \I__2897\ : InMux
    port map (
            O => \N__16226\,
            I => \N__16223\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__16223\,
            I => \N__16220\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__16217\,
            I => \N__16214\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__16214\,
            I => scaler_4_data_5
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__16211\,
            I => \N__16208\
        );

    \I__2891\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16205\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__16205\,
            I => \scaler_2.un2_source_data_0_cry_1_c_RNO_0\
        );

    \I__2889\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16197\
        );

    \I__2888\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16194\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__16200\,
            I => \N__16191\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__16197\,
            I => \N__16187\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16184\
        );

    \I__2884\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16179\
        );

    \I__2883\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16179\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__16187\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__16184\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__16179\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__2879\ : InMux
    port map (
            O => \N__16172\,
            I => \scaler_2.un2_source_data_0_cry_1\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__2877\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16160\
        );

    \I__2876\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16160\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__16160\,
            I => \scaler_2.un3_source_data_0_cry_1_c_RNILSPH\
        );

    \I__2874\ : InMux
    port map (
            O => \N__16157\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_17\
        );

    \I__2873\ : InMux
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__16151\,
            I => \ppm_encoder_1.un1_init_pulses_10_18\
        );

    \I__2871\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16143\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__16147\,
            I => \N__16140\
        );

    \I__2869\ : InMux
    port map (
            O => \N__16146\,
            I => \N__16136\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__16143\,
            I => \N__16133\
        );

    \I__2867\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16128\
        );

    \I__2866\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16128\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__16136\,
            I => \N__16120\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__16133\,
            I => \N__16115\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__16128\,
            I => \N__16115\
        );

    \I__2862\ : InMux
    port map (
            O => \N__16127\,
            I => \N__16108\
        );

    \I__2861\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16108\
        );

    \I__2860\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16108\
        );

    \I__2859\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16103\
        );

    \I__2858\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16103\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__16120\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__16115\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__16108\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__16103\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2853\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16091\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__16091\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_18\
        );

    \I__2851\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16085\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__2849\ : Span4Mux_v
    port map (
            O => \N__16082\,
            I => \N__16079\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__16079\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__16076\,
            I => \N__16073\
        );

    \I__2846\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16068\
        );

    \I__2845\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16065\
        );

    \I__2844\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16062\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__16068\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__16065\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__16062\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__2840\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16052\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__16052\,
            I => \N__16047\
        );

    \I__2838\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16042\
        );

    \I__2837\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16042\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__16047\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__16042\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__16037\,
            I => \N__16034\
        );

    \I__2833\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16030\
        );

    \I__2832\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16027\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16024\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__16027\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__16024\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__16019\,
            I => \N__16013\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__16018\,
            I => \N__16010\
        );

    \I__2826\ : InMux
    port map (
            O => \N__16017\,
            I => \N__16001\
        );

    \I__2825\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16001\
        );

    \I__2824\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16001\
        );

    \I__2823\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16001\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__2821\ : Span12Mux_s8_v
    port map (
            O => \N__15998\,
            I => \N__15994\
        );

    \I__2820\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15991\
        );

    \I__2819\ : Odrv12
    port map (
            O => \N__15994\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_162_d\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__15991\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_162_d\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__15986\,
            I => \N__15982\
        );

    \I__2816\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15979\
        );

    \I__2815\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15975\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__15979\,
            I => \N__15972\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__15978\,
            I => \N__15969\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__15975\,
            I => \N__15964\
        );

    \I__2811\ : Span4Mux_h
    port map (
            O => \N__15972\,
            I => \N__15964\
        );

    \I__2810\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15961\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__15964\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__15961\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__2807\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15951\
        );

    \I__2806\ : InMux
    port map (
            O => \N__15955\,
            I => \N__15946\
        );

    \I__2805\ : InMux
    port map (
            O => \N__15954\,
            I => \N__15946\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__15951\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__15946\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__2802\ : InMux
    port map (
            O => \N__15941\,
            I => \N__15938\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__15938\,
            I => \N__15935\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__15935\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_16\
        );

    \I__2799\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__15929\,
            I => \ppm_encoder_1.un1_init_pulses_10_10\
        );

    \I__2797\ : InMux
    port map (
            O => \N__15926\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_9\
        );

    \I__2796\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__15920\,
            I => \N__15916\
        );

    \I__2794\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15913\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__15916\,
            I => \N__15910\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__15913\,
            I => \N__15907\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__15910\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__15907\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__2788\ : InMux
    port map (
            O => \N__15899\,
            I => \N__15896\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__15896\,
            I => \N__15893\
        );

    \I__2786\ : Odrv12
    port map (
            O => \N__15893\,
            I => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\
        );

    \I__2785\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15887\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__15887\,
            I => \ppm_encoder_1.un1_init_pulses_10_11\
        );

    \I__2783\ : InMux
    port map (
            O => \N__15884\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_10\
        );

    \I__2782\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15878\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__15878\,
            I => \ppm_encoder_1.un1_init_pulses_10_12\
        );

    \I__2780\ : InMux
    port map (
            O => \N__15875\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_11\
        );

    \I__2779\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15869\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__15869\,
            I => \N__15866\
        );

    \I__2777\ : Span4Mux_h
    port map (
            O => \N__15866\,
            I => \N__15863\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__15863\,
            I => \ppm_encoder_1.un1_init_pulses_10_13\
        );

    \I__2775\ : InMux
    port map (
            O => \N__15860\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_12\
        );

    \I__2774\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15854\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__15854\,
            I => \ppm_encoder_1.un1_init_pulses_10_14\
        );

    \I__2772\ : InMux
    port map (
            O => \N__15851\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_13\
        );

    \I__2771\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15845\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__15845\,
            I => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__15842\,
            I => \N__15839\
        );

    \I__2768\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15836\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__15836\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\
        );

    \I__2766\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15830\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__15830\,
            I => \ppm_encoder_1.un1_init_pulses_10_15\
        );

    \I__2764\ : InMux
    port map (
            O => \N__15827\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_14\
        );

    \I__2763\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15821\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__15821\,
            I => \ppm_encoder_1.un1_init_pulses_10_16\
        );

    \I__2761\ : InMux
    port map (
            O => \N__15818\,
            I => \bfn_9_26_0_\
        );

    \I__2760\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__15812\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_17\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__15809\,
            I => \N__15806\
        );

    \I__2757\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15803\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__15803\,
            I => \ppm_encoder_1.un1_init_pulses_10_17\
        );

    \I__2755\ : InMux
    port map (
            O => \N__15800\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_16\
        );

    \I__2754\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15794\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__15794\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__15791\,
            I => \N__15788\
        );

    \I__2751\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15785\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__15785\,
            I => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__2748\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__15773\,
            I => \ppm_encoder_1.un1_init_pulses_10_2\
        );

    \I__2745\ : InMux
    port map (
            O => \N__15770\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_1\
        );

    \I__2744\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__15764\,
            I => \N__15760\
        );

    \I__2742\ : InMux
    port map (
            O => \N__15763\,
            I => \N__15757\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__15760\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__15757\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__15752\,
            I => \N__15749\
        );

    \I__2738\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__15743\,
            I => \ppm_encoder_1.init_pulses_RNI60223Z0Z_3\
        );

    \I__2735\ : InMux
    port map (
            O => \N__15740\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_2\
        );

    \I__2734\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15733\
        );

    \I__2733\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15730\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__15733\,
            I => \N__15727\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15724\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__15727\,
            I => \N__15721\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__15724\,
            I => \N__15718\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__15721\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__15718\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__15713\,
            I => \N__15710\
        );

    \I__2725\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15707\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__15707\,
            I => \N__15704\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__15704\,
            I => \ppm_encoder_1.aileron_esr_RNI8CGI5Z0Z_4\
        );

    \I__2722\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15698\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__15692\,
            I => \ppm_encoder_1.un1_init_pulses_10_4\
        );

    \I__2718\ : InMux
    port map (
            O => \N__15689\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_3\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__2716\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__15680\,
            I => \ppm_encoder_1.aileron_esr_RNIDHGI5Z0Z_5\
        );

    \I__2714\ : InMux
    port map (
            O => \N__15677\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_4\
        );

    \I__2713\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__15671\,
            I => \N__15668\
        );

    \I__2711\ : Span4Mux_h
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__15665\,
            I => \ppm_encoder_1.un1_init_pulses_10_6\
        );

    \I__2709\ : InMux
    port map (
            O => \N__15662\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_5\
        );

    \I__2708\ : InMux
    port map (
            O => \N__15659\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_6\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__2706\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15650\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__15650\,
            I => \N__15647\
        );

    \I__2704\ : Odrv12
    port map (
            O => \N__15647\,
            I => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\
        );

    \I__2703\ : InMux
    port map (
            O => \N__15644\,
            I => \bfn_9_25_0_\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__2701\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__2699\ : Odrv12
    port map (
            O => \N__15632\,
            I => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\
        );

    \I__2698\ : InMux
    port map (
            O => \N__15629\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_8\
        );

    \I__2697\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15621\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__15625\,
            I => \N__15618\
        );

    \I__2695\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15612\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__15621\,
            I => \N__15609\
        );

    \I__2693\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15604\
        );

    \I__2692\ : InMux
    port map (
            O => \N__15617\,
            I => \N__15604\
        );

    \I__2691\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15599\
        );

    \I__2690\ : InMux
    port map (
            O => \N__15615\,
            I => \N__15599\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__15612\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__2688\ : Odrv12
    port map (
            O => \N__15609\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__15604\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__15599\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__15590\,
            I => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\
        );

    \I__2684\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15584\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__15584\,
            I => \ppm_encoder_1.un2_throttle_iv_1_5\
        );

    \I__2682\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15575\
        );

    \I__2681\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15575\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__15575\,
            I => \N__15572\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__15572\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__2678\ : InMux
    port map (
            O => \N__15569\,
            I => \N__15563\
        );

    \I__2677\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15563\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__15560\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__15557\,
            I => \ppm_encoder_1.N_300_cascade_\
        );

    \I__2673\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15551\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__2671\ : Odrv12
    port map (
            O => \N__15548\,
            I => scaler_2_data_5
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__15545\,
            I => \N__15541\
        );

    \I__2669\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15538\
        );

    \I__2668\ : InMux
    port map (
            O => \N__15541\,
            I => \N__15535\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__15538\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__15535\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__2665\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15526\
        );

    \I__2664\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15523\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__15526\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__15523\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__2661\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__15515\,
            I => \N__15511\
        );

    \I__2659\ : InMux
    port map (
            O => \N__15514\,
            I => \N__15508\
        );

    \I__2658\ : Odrv12
    port map (
            O => \N__15511\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__15508\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__15503\,
            I => \N__15500\
        );

    \I__2655\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15497\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__15494\,
            I => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\
        );

    \I__2652\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15488\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__15488\,
            I => \ppm_encoder_1.un1_init_pulses_10_1\
        );

    \I__2650\ : InMux
    port map (
            O => \N__15485\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_0\
        );

    \I__2649\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__15479\,
            I => \ppm_encoder_1.un2_throttle_iv_1_9\
        );

    \I__2647\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15471\
        );

    \I__2646\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15468\
        );

    \I__2645\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15465\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__15471\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__15468\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__15465\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__15458\,
            I => \N__15453\
        );

    \I__2640\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15450\
        );

    \I__2639\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15447\
        );

    \I__2638\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15444\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__15450\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__15447\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__15444\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__2634\ : InMux
    port map (
            O => \N__15437\,
            I => \N__15433\
        );

    \I__2633\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15430\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__15433\,
            I => \N__15425\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__15430\,
            I => \N__15425\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__15425\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__2629\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15418\
        );

    \I__2628\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15415\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__15418\,
            I => \N__15412\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__15415\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__15412\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__15407\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\
        );

    \I__2623\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15400\
        );

    \I__2622\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15397\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__15400\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__15397\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\
        );

    \I__2619\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15388\
        );

    \I__2618\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15385\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__15388\,
            I => \N__15380\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15380\
        );

    \I__2615\ : Span4Mux_v
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__15377\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__15371\,
            I => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\
        );

    \I__2611\ : InMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__15365\,
            I => \ppm_encoder_1.un2_throttle_iv_1_4\
        );

    \I__2609\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__15359\,
            I => \ppm_encoder_1.un2_throttle_iv_1_11\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__15356\,
            I => \ppm_encoder_1.N_306_cascade_\
        );

    \I__2606\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15344\
        );

    \I__2605\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15344\
        );

    \I__2604\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15344\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__15344\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\
        );

    \I__2601\ : InMux
    port map (
            O => \N__15338\,
            I => \N__15335\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__15335\,
            I => \ppm_encoder_1.un2_throttle_iv_1_8\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__15332\,
            I => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\
        );

    \I__2598\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15322\
        );

    \I__2597\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15322\
        );

    \I__2596\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15319\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__15322\,
            I => \N__15310\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__15319\,
            I => \N__15310\
        );

    \I__2593\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15306\
        );

    \I__2592\ : InMux
    port map (
            O => \N__15317\,
            I => \N__15301\
        );

    \I__2591\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15301\
        );

    \I__2590\ : InMux
    port map (
            O => \N__15315\,
            I => \N__15298\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__15310\,
            I => \N__15295\
        );

    \I__2588\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15292\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__15306\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__15301\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__15298\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__15295\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__15292\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2582\ : InMux
    port map (
            O => \N__15281\,
            I => \N__15275\
        );

    \I__2581\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15275\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__15275\,
            I => \uart_frame_decoder.count8_THRU_CO\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \N__15263\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__15271\,
            I => \N__15260\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__15270\,
            I => \N__15257\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__15269\,
            I => \N__15254\
        );

    \I__2575\ : InMux
    port map (
            O => \N__15268\,
            I => \N__15248\
        );

    \I__2574\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15243\
        );

    \I__2573\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15240\
        );

    \I__2572\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15225\
        );

    \I__2571\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15225\
        );

    \I__2570\ : InMux
    port map (
            O => \N__15257\,
            I => \N__15225\
        );

    \I__2569\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15225\
        );

    \I__2568\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15225\
        );

    \I__2567\ : InMux
    port map (
            O => \N__15252\,
            I => \N__15225\
        );

    \I__2566\ : InMux
    port map (
            O => \N__15251\,
            I => \N__15225\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__15248\,
            I => \N__15222\
        );

    \I__2564\ : InMux
    port map (
            O => \N__15247\,
            I => \N__15218\
        );

    \I__2563\ : InMux
    port map (
            O => \N__15246\,
            I => \N__15215\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__15243\,
            I => \N__15212\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__15240\,
            I => \N__15209\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__15225\,
            I => \N__15206\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__15222\,
            I => \N__15203\
        );

    \I__2558\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15200\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__15218\,
            I => \N__15193\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__15215\,
            I => \N__15193\
        );

    \I__2555\ : Sp12to4
    port map (
            O => \N__15212\,
            I => \N__15193\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__15209\,
            I => \N__15190\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__15206\,
            I => \N__15187\
        );

    \I__2552\ : Span4Mux_v
    port map (
            O => \N__15203\,
            I => \N__15184\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__15200\,
            I => \N__15181\
        );

    \I__2550\ : Span12Mux_v
    port map (
            O => \N__15193\,
            I => \N__15178\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__15190\,
            I => uart_input_pc_sync
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__15187\,
            I => uart_input_pc_sync
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__15184\,
            I => uart_input_pc_sync
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__15181\,
            I => uart_input_pc_sync
        );

    \I__2545\ : Odrv12
    port map (
            O => \N__15178\,
            I => uart_input_pc_sync
        );

    \I__2544\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15160\
        );

    \I__2543\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15160\
        );

    \I__2542\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15157\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__15160\,
            I => \N__15154\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__15157\,
            I => \N__15151\
        );

    \I__2539\ : Span4Mux_h
    port map (
            O => \N__15154\,
            I => \N__15148\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__15151\,
            I => \N__15145\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__15148\,
            I => \N__15142\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__15145\,
            I => \uart_pc.state_1_sqmuxa\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__15142\,
            I => \uart_pc.state_1_sqmuxa\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__15137\,
            I => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\
        );

    \I__2533\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15131\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__15131\,
            I => \scaler_2.N_520_i_l_ofxZ0\
        );

    \I__2531\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15125\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__15125\,
            I => \N__15122\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__15122\,
            I => \N__15119\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__15119\,
            I => scaler_1_data_5
        );

    \I__2527\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15113\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__15110\,
            I => \N__15107\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__15107\,
            I => scaler_3_data_5
        );

    \I__2523\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__15101\,
            I => \N__15098\
        );

    \I__2521\ : Span4Mux_v
    port map (
            O => \N__15098\,
            I => \N__15094\
        );

    \I__2520\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15091\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__15094\,
            I => scaler_1_data_4
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__15091\,
            I => scaler_1_data_4
        );

    \I__2517\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15082\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__15085\,
            I => \N__15077\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__15082\,
            I => \N__15074\
        );

    \I__2514\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15071\
        );

    \I__2513\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15068\
        );

    \I__2512\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15065\
        );

    \I__2511\ : Span4Mux_v
    port map (
            O => \N__15074\,
            I => \N__15060\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__15071\,
            I => \N__15060\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__15068\,
            I => \N__15057\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__15065\,
            I => \N__15054\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__15060\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__15057\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__15054\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__2504\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15043\
        );

    \I__2503\ : InMux
    port map (
            O => \N__15046\,
            I => \N__15040\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__15043\,
            I => \N__15033\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__15040\,
            I => \N__15033\
        );

    \I__2500\ : InMux
    port map (
            O => \N__15039\,
            I => \N__15030\
        );

    \I__2499\ : InMux
    port map (
            O => \N__15038\,
            I => \N__15027\
        );

    \I__2498\ : Odrv12
    port map (
            O => \N__15033\,
            I => \frame_decoder_CH2data_0\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__15030\,
            I => \frame_decoder_CH2data_0\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__15027\,
            I => \frame_decoder_CH2data_0\
        );

    \I__2495\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15017\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__15017\,
            I => \N__15013\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__15016\,
            I => \N__15010\
        );

    \I__2492\ : Span4Mux_h
    port map (
            O => \N__15013\,
            I => \N__15007\
        );

    \I__2491\ : InMux
    port map (
            O => \N__15010\,
            I => \N__15004\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__15007\,
            I => scaler_2_data_4
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__15004\,
            I => scaler_2_data_4
        );

    \I__2488\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14995\
        );

    \I__2487\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14992\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__14995\,
            I => \N__14989\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__14992\,
            I => \N__14986\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__14989\,
            I => scaler_3_data_4
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__14986\,
            I => scaler_3_data_4
        );

    \I__2482\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14978\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__14978\,
            I => \N__14974\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__14977\,
            I => \N__14971\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__14974\,
            I => \N__14968\
        );

    \I__2478\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14965\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__14968\,
            I => scaler_4_data_4
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__14965\,
            I => scaler_4_data_4
        );

    \I__2475\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14957\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__14957\,
            I => \frame_decoder_CH2data_4\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__14954\,
            I => \N__14951\
        );

    \I__2472\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14948\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__14948\,
            I => \frame_decoder_OFF2data_4\
        );

    \I__2470\ : InMux
    port map (
            O => \N__14945\,
            I => \scaler_2.un3_source_data_0_cry_3\
        );

    \I__2469\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14939\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__14939\,
            I => \frame_decoder_CH2data_5\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__14936\,
            I => \N__14933\
        );

    \I__2466\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14930\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__14930\,
            I => \frame_decoder_OFF2data_5\
        );

    \I__2464\ : InMux
    port map (
            O => \N__14927\,
            I => \scaler_2.un3_source_data_0_cry_4\
        );

    \I__2463\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__14921\,
            I => \frame_decoder_CH2data_6\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__2460\ : InMux
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__14912\,
            I => \frame_decoder_OFF2data_6\
        );

    \I__2458\ : InMux
    port map (
            O => \N__14909\,
            I => \scaler_2.un3_source_data_0_cry_5\
        );

    \I__2457\ : InMux
    port map (
            O => \N__14906\,
            I => \scaler_2.un3_source_data_0_cry_6\
        );

    \I__2456\ : InMux
    port map (
            O => \N__14903\,
            I => \bfn_9_15_0_\
        );

    \I__2455\ : InMux
    port map (
            O => \N__14900\,
            I => \scaler_2.un3_source_data_0_cry_8\
        );

    \I__2454\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14894\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__14894\,
            I => \N__14890\
        );

    \I__2452\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14887\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__14890\,
            I => \N__14884\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__14887\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__14884\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__2448\ : InMux
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__2446\ : Sp12to4
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__2445\ : Odrv12
    port map (
            O => \N__14870\,
            I => \uart_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__14867\,
            I => \uart_frame_decoder.source_CH2data_1_sqmuxa_cascade_\
        );

    \I__2443\ : InMux
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__14861\,
            I => \frame_decoder_CH2data_1\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__14858\,
            I => \N__14855\
        );

    \I__2440\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__14852\,
            I => \frame_decoder_OFF2data_1\
        );

    \I__2438\ : InMux
    port map (
            O => \N__14849\,
            I => \scaler_2.un3_source_data_0_cry_0\
        );

    \I__2437\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__14843\,
            I => \frame_decoder_CH2data_2\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__14840\,
            I => \N__14837\
        );

    \I__2434\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14834\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__14834\,
            I => \frame_decoder_OFF2data_2\
        );

    \I__2432\ : InMux
    port map (
            O => \N__14831\,
            I => \scaler_2.un3_source_data_0_cry_1\
        );

    \I__2431\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__14825\,
            I => \frame_decoder_CH2data_3\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__2428\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14816\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__14816\,
            I => \frame_decoder_OFF2data_3\
        );

    \I__2426\ : InMux
    port map (
            O => \N__14813\,
            I => \scaler_2.un3_source_data_0_cry_2\
        );

    \I__2425\ : SRMux
    port map (
            O => \N__14810\,
            I => \N__14805\
        );

    \I__2424\ : SRMux
    port map (
            O => \N__14809\,
            I => \N__14802\
        );

    \I__2423\ : SRMux
    port map (
            O => \N__14808\,
            I => \N__14799\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__14805\,
            I => \N__14796\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__14802\,
            I => \N__14791\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__14799\,
            I => \N__14791\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__14796\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__14791\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__2417\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__14783\,
            I => \uart_frame_decoder.state_1_ns_i_i_0_0\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__14780\,
            I => \N__14777\
        );

    \I__2414\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14774\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__14774\,
            I => \uart_frame_decoder.N_39_i_1\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__14771\,
            I => \N__14766\
        );

    \I__2411\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14763\
        );

    \I__2410\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14758\
        );

    \I__2409\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14758\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__14763\,
            I => \uart_frame_decoder.state_1Z0Z_0\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__14758\,
            I => \uart_frame_decoder.state_1Z0Z_0\
        );

    \I__2406\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14749\
        );

    \I__2405\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14746\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__14749\,
            I => \uart_frame_decoder.state_1Z0Z_9\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__14746\,
            I => \uart_frame_decoder.state_1Z0Z_9\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__2401\ : InMux
    port map (
            O => \N__14738\,
            I => \N__14735\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__14735\,
            I => \uart_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__14732\,
            I => \uart_frame_decoder.source_offset4data_1_sqmuxa_cascade_\
        );

    \I__2398\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14722\
        );

    \I__2396\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14718\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__14722\,
            I => \N__14715\
        );

    \I__2394\ : InMux
    port map (
            O => \N__14721\,
            I => \N__14712\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__14718\,
            I => \uart_frame_decoder.countZ0Z_2\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__14715\,
            I => \uart_frame_decoder.countZ0Z_2\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__14712\,
            I => \uart_frame_decoder.countZ0Z_2\
        );

    \I__2390\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14701\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__14704\,
            I => \N__14698\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__14701\,
            I => \N__14694\
        );

    \I__2387\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14688\
        );

    \I__2386\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14688\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__14694\,
            I => \N__14685\
        );

    \I__2384\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14682\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__14688\,
            I => \uart_frame_decoder.countZ0Z_1\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__14685\,
            I => \uart_frame_decoder.countZ0Z_1\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__14682\,
            I => \uart_frame_decoder.countZ0Z_1\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \uart_frame_decoder.state_1_RNINMHJZ0Z_10_cascade_\
        );

    \I__2379\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14666\
        );

    \I__2378\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14666\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__14666\,
            I => \uart_frame_decoder.state_1_ns_0_i_o2_0_10\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__2375\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14657\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__14657\,
            I => \ppm_encoder_1.un1_init_pulses_11_10\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__2372\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__14648\,
            I => \ppm_encoder_1.un1_init_pulses_11_16\
        );

    \I__2370\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__14642\,
            I => \ppm_encoder_1.un1_init_pulses_11_17\
        );

    \I__2368\ : InMux
    port map (
            O => \N__14639\,
            I => \N__14636\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__14636\,
            I => \ppm_encoder_1.un1_init_pulses_11_4\
        );

    \I__2366\ : InMux
    port map (
            O => \N__14633\,
            I => \N__14630\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__14630\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_4\
        );

    \I__2364\ : InMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__14624\,
            I => \N__14620\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__14623\,
            I => \N__14617\
        );

    \I__2361\ : Span4Mux_h
    port map (
            O => \N__14620\,
            I => \N__14614\
        );

    \I__2360\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14611\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__14614\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__14611\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__2357\ : CEMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__14603\,
            I => \N__14598\
        );

    \I__2355\ : CEMux
    port map (
            O => \N__14602\,
            I => \N__14595\
        );

    \I__2354\ : CEMux
    port map (
            O => \N__14601\,
            I => \N__14592\
        );

    \I__2353\ : Span4Mux_h
    port map (
            O => \N__14598\,
            I => \N__14589\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__14595\,
            I => \N__14586\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__14592\,
            I => \N__14583\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__14589\,
            I => \uart_pc.state_1_sqmuxa_0\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__14586\,
            I => \uart_pc.state_1_sqmuxa_0\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__14583\,
            I => \uart_pc.state_1_sqmuxa_0\
        );

    \I__2347\ : InMux
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__14573\,
            I => \N__14570\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__14570\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_12\
        );

    \I__2344\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14564\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__14564\,
            I => \N__14561\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__14561\,
            I => \ppm_encoder_1.un1_init_pulses_11_14\
        );

    \I__2341\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14555\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__14555\,
            I => \ppm_encoder_1.un1_init_pulses_11_15\
        );

    \I__2339\ : InMux
    port map (
            O => \N__14552\,
            I => \N__14549\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__14549\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_15\
        );

    \I__2337\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14543\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__14543\,
            I => \N__14540\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__14540\,
            I => \ppm_encoder_1.un1_init_pulses_11_18\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__14537\,
            I => \N__14534\
        );

    \I__2333\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14531\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__14531\,
            I => \N__14528\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__14528\,
            I => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__14525\,
            I => \N__14521\
        );

    \I__2329\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14516\
        );

    \I__2328\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14516\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N__14506\
        );

    \I__2326\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14499\
        );

    \I__2325\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14499\
        );

    \I__2324\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14499\
        );

    \I__2323\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14490\
        );

    \I__2322\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14490\
        );

    \I__2321\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14490\
        );

    \I__2320\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14490\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__14506\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__14499\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__14490\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__2316\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14480\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__14480\,
            I => \N__14477\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__14477\,
            I => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\
        );

    \I__2313\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14471\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__14471\,
            I => \N__14468\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__14468\,
            I => \ppm_encoder_1.un1_init_pulses_11_2\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \ppm_encoder_1.un1_init_pulses_0_2_cascade_\
        );

    \I__2309\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14459\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__14459\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_2\
        );

    \I__2307\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__14450\,
            I => \ppm_encoder_1.un1_init_pulses_11_11\
        );

    \I__2304\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14444\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__14444\,
            I => \N__14441\
        );

    \I__2302\ : Span4Mux_v
    port map (
            O => \N__14441\,
            I => \N__14438\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__14438\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_11\
        );

    \I__2300\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14432\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__14432\,
            I => \N__14429\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__14429\,
            I => \ppm_encoder_1.un1_init_pulses_11_12\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__14426\,
            I => \N__14423\
        );

    \I__2296\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14420\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__14420\,
            I => \N__14417\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__14417\,
            I => \ppm_encoder_1.un1_init_pulses_11_1\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__14414\,
            I => \ppm_encoder_1.PPM_STATE_62_d_cascade_\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__14411\,
            I => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\
        );

    \I__2291\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14405\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__14405\,
            I => \N__14402\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__14402\,
            I => \N__14399\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__14399\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_10\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__14396\,
            I => \N__14392\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__14395\,
            I => \N__14389\
        );

    \I__2285\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14386\
        );

    \I__2284\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__14386\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__14383\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__2281\ : InMux
    port map (
            O => \N__14378\,
            I => \N__14375\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__14375\,
            I => \N__14372\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__14372\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__14369\,
            I => \N__14364\
        );

    \I__2277\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14361\
        );

    \I__2276\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14356\
        );

    \I__2275\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14356\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__14361\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__14356\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__2272\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14345\
        );

    \I__2271\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14338\
        );

    \I__2270\ : InMux
    port map (
            O => \N__14349\,
            I => \N__14338\
        );

    \I__2269\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14338\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__14345\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__14338\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__14333\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__14330\,
            I => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\
        );

    \I__2264\ : InMux
    port map (
            O => \N__14327\,
            I => \N__14324\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__14324\,
            I => \N__14321\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__14321\,
            I => \N__14318\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__14318\,
            I => \ppm_encoder_1.N_299\
        );

    \I__2260\ : InMux
    port map (
            O => \N__14315\,
            I => \uart_frame_decoder.count8\
        );

    \I__2259\ : CEMux
    port map (
            O => \N__14312\,
            I => \N__14309\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__14309\,
            I => \N__14305\
        );

    \I__2257\ : CEMux
    port map (
            O => \N__14308\,
            I => \N__14302\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__14305\,
            I => \N__14297\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__14302\,
            I => \N__14297\
        );

    \I__2254\ : Span4Mux_h
    port map (
            O => \N__14297\,
            I => \N__14294\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__14294\,
            I => \uart_frame_decoder.source_CH1data_1_sqmuxa_0\
        );

    \I__2252\ : InMux
    port map (
            O => \N__14291\,
            I => \scaler_1.un3_source_data_0_cry_8\
        );

    \I__2251\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14285\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__14285\,
            I => \scaler_1.un3_source_data_0_axb_7\
        );

    \I__2249\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14276\
        );

    \I__2248\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14276\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__14276\,
            I => \frame_decoder_CH1data_7\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__14273\,
            I => \N__14270\
        );

    \I__2245\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14264\
        );

    \I__2244\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14264\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__14264\,
            I => \frame_decoder_OFF1data_7\
        );

    \I__2242\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14258\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__14258\,
            I => \scaler_1.N_508_i_l_ofxZ0\
        );

    \I__2240\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14249\
        );

    \I__2239\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14249\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__14249\,
            I => \N__14246\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__14246\,
            I => \uart_frame_decoder.count_RNIHJ501Z0Z_0\
        );

    \I__2236\ : InMux
    port map (
            O => \N__14243\,
            I => \N__14240\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__14240\,
            I => \uart_frame_decoder.count8_axb_1\
        );

    \I__2234\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14234\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__14234\,
            I => \uart_frame_decoder.count_i_2\
        );

    \I__2232\ : InMux
    port map (
            O => \N__14231\,
            I => \N__14228\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__14228\,
            I => \frame_decoder_CH1data_1\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__2229\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14219\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__14219\,
            I => \frame_decoder_OFF1data_1\
        );

    \I__2227\ : InMux
    port map (
            O => \N__14216\,
            I => \scaler_1.un3_source_data_0_cry_0\
        );

    \I__2226\ : InMux
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__14210\,
            I => \frame_decoder_CH1data_2\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__2223\ : InMux
    port map (
            O => \N__14204\,
            I => \N__14201\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__14201\,
            I => \frame_decoder_OFF1data_2\
        );

    \I__2221\ : InMux
    port map (
            O => \N__14198\,
            I => \scaler_1.un3_source_data_0_cry_1\
        );

    \I__2220\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__14192\,
            I => \frame_decoder_CH1data_3\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__14189\,
            I => \N__14186\
        );

    \I__2217\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14183\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__14183\,
            I => \frame_decoder_OFF1data_3\
        );

    \I__2215\ : InMux
    port map (
            O => \N__14180\,
            I => \scaler_1.un3_source_data_0_cry_2\
        );

    \I__2214\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14174\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__14174\,
            I => \frame_decoder_CH1data_4\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__14171\,
            I => \N__14168\
        );

    \I__2211\ : InMux
    port map (
            O => \N__14168\,
            I => \N__14165\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__14165\,
            I => \frame_decoder_OFF1data_4\
        );

    \I__2209\ : InMux
    port map (
            O => \N__14162\,
            I => \scaler_1.un3_source_data_0_cry_3\
        );

    \I__2208\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14156\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__14156\,
            I => \frame_decoder_CH1data_5\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__14153\,
            I => \N__14150\
        );

    \I__2205\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14147\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__14147\,
            I => \frame_decoder_OFF1data_5\
        );

    \I__2203\ : InMux
    port map (
            O => \N__14144\,
            I => \scaler_1.un3_source_data_0_cry_4\
        );

    \I__2202\ : InMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__14138\,
            I => \frame_decoder_CH1data_6\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__14135\,
            I => \N__14132\
        );

    \I__2199\ : InMux
    port map (
            O => \N__14132\,
            I => \N__14129\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__14129\,
            I => \frame_decoder_OFF1data_6\
        );

    \I__2197\ : InMux
    port map (
            O => \N__14126\,
            I => \scaler_1.un3_source_data_0_cry_5\
        );

    \I__2196\ : InMux
    port map (
            O => \N__14123\,
            I => \scaler_1.un3_source_data_0_cry_6\
        );

    \I__2195\ : InMux
    port map (
            O => \N__14120\,
            I => \bfn_8_18_0_\
        );

    \I__2194\ : CEMux
    port map (
            O => \N__14117\,
            I => \N__14114\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__14114\,
            I => \uart_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__2192\ : InMux
    port map (
            O => \N__14111\,
            I => \N__14107\
        );

    \I__2191\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14104\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__14107\,
            I => \uart_frame_decoder.WDTZ0Z_6\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__14104\,
            I => \uart_frame_decoder.WDTZ0Z_6\
        );

    \I__2188\ : InMux
    port map (
            O => \N__14099\,
            I => \N__14094\
        );

    \I__2187\ : InMux
    port map (
            O => \N__14098\,
            I => \N__14089\
        );

    \I__2186\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14089\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__14094\,
            I => \uart_frame_decoder.WDTZ0Z_11\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__14089\,
            I => \uart_frame_decoder.WDTZ0Z_11\
        );

    \I__2183\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14080\
        );

    \I__2182\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14077\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__14080\,
            I => \uart_frame_decoder.WDTZ0Z_10\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__14077\,
            I => \uart_frame_decoder.WDTZ0Z_10\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__14072\,
            I => \N__14068\
        );

    \I__2178\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__2177\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14062\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__14065\,
            I => \uart_frame_decoder.WDTZ0Z_13\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__14062\,
            I => \uart_frame_decoder.WDTZ0Z_13\
        );

    \I__2174\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14052\
        );

    \I__2173\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14047\
        );

    \I__2172\ : InMux
    port map (
            O => \N__14055\,
            I => \N__14047\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__14052\,
            I => \uart_frame_decoder.WDTZ0Z_12\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__14047\,
            I => \uart_frame_decoder.WDTZ0Z_12\
        );

    \I__2169\ : InMux
    port map (
            O => \N__14042\,
            I => \N__14038\
        );

    \I__2168\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__14038\,
            I => \uart_frame_decoder.WDTZ0Z_7\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__14035\,
            I => \uart_frame_decoder.WDTZ0Z_7\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__14030\,
            I => \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_\
        );

    \I__2164\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14024\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__14024\,
            I => \uart_frame_decoder.WDT8lto13_1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__14021\,
            I => \N__14018\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__14015\,
            I => \uart_frame_decoder.WDT8lt14_0\
        );

    \I__2159\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__14009\,
            I => \N__14005\
        );

    \I__2157\ : InMux
    port map (
            O => \N__14008\,
            I => \N__14001\
        );

    \I__2156\ : Span4Mux_h
    port map (
            O => \N__14005\,
            I => \N__13998\
        );

    \I__2155\ : InMux
    port map (
            O => \N__14004\,
            I => \N__13995\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__14001\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__13998\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__13995\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \uart_frame_decoder.WDT8lt14_0_cascade_\
        );

    \I__2150\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__13982\,
            I => \N__13978\
        );

    \I__2148\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13974\
        );

    \I__2147\ : Span4Mux_h
    port map (
            O => \N__13978\,
            I => \N__13971\
        );

    \I__2146\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13968\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__13974\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__13971\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__13968\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__13961\,
            I => \N__13957\
        );

    \I__2141\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13954\
        );

    \I__2140\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__13954\,
            I => \uart_frame_decoder.WDT8_0_i\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__13951\,
            I => \uart_frame_decoder.WDT8_0_i\
        );

    \I__2137\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13942\
        );

    \I__2136\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13939\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__13942\,
            I => \uart_frame_decoder.WDTZ0Z_8\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__13939\,
            I => \uart_frame_decoder.WDTZ0Z_8\
        );

    \I__2133\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13930\
        );

    \I__2132\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13927\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__13930\,
            I => \uart_frame_decoder.WDTZ0Z_5\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__13927\,
            I => \uart_frame_decoder.WDTZ0Z_5\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__13922\,
            I => \N__13918\
        );

    \I__2128\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13915\
        );

    \I__2127\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13912\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__13915\,
            I => \uart_frame_decoder.WDTZ0Z_9\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__13912\,
            I => \uart_frame_decoder.WDTZ0Z_9\
        );

    \I__2124\ : InMux
    port map (
            O => \N__13907\,
            I => \N__13903\
        );

    \I__2123\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13900\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__13903\,
            I => \uart_frame_decoder.WDTZ0Z_4\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__13900\,
            I => \uart_frame_decoder.WDTZ0Z_4\
        );

    \I__2120\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__13892\,
            I => \uart_frame_decoder.WDT_RNIQAB11Z0Z_4\
        );

    \I__2118\ : SRMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__13886\,
            I => \N__13882\
        );

    \I__2116\ : SRMux
    port map (
            O => \N__13885\,
            I => \N__13879\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__13882\,
            I => \N__13876\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__13879\,
            I => \N__13873\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__13876\,
            I => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__13873\,
            I => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__2111\ : CEMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__2109\ : Span4Mux_h
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__2108\ : Span4Mux_h
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__13856\,
            I => \uart_frame_decoder.source_offset2data_1_sqmuxa_0\
        );

    \I__2106\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13849\
        );

    \I__2105\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13846\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__13849\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__13846\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__2102\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13837\
        );

    \I__2101\ : InMux
    port map (
            O => \N__13840\,
            I => \N__13834\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__13837\,
            I => \uart_frame_decoder.source_offset1data_1_sqmuxa\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__13834\,
            I => \uart_frame_decoder.source_offset1data_1_sqmuxa\
        );

    \I__2098\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13825\
        );

    \I__2097\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__13825\,
            I => \uart_frame_decoder.state_1Z0Z_7\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__13822\,
            I => \uart_frame_decoder.state_1Z0Z_7\
        );

    \I__2094\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13814\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__13811\,
            I => \uart_frame_decoder.source_offset2data_1_sqmuxa\
        );

    \I__2091\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13804\
        );

    \I__2090\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13801\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__13804\,
            I => \uart_frame_decoder.state_1Z0Z_8\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__13801\,
            I => \uart_frame_decoder.state_1Z0Z_8\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__13796\,
            I => \N__13793\
        );

    \I__2086\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13789\
        );

    \I__2085\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13786\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__13789\,
            I => \uart_frame_decoder.source_offset3data_1_sqmuxa\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__13786\,
            I => \uart_frame_decoder.source_offset3data_1_sqmuxa\
        );

    \I__2082\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13778\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__13778\,
            I => \uart_frame_decoder.N_138_4\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__13775\,
            I => \uart_frame_decoder.N_138_4_cascade_\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__13772\,
            I => \N__13769\
        );

    \I__2078\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13766\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__13766\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\
        );

    \I__2076\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13756\
        );

    \I__2075\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13749\
        );

    \I__2074\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13749\
        );

    \I__2073\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13749\
        );

    \I__2072\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13746\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__13756\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__13749\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__13746\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__2068\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__13736\,
            I => \uart_frame_decoder.state_1_RNO_2Z0Z_0\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__13733\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__13730\,
            I => \uart_frame_decoder.N_85_cascade_\
        );

    \I__2064\ : InMux
    port map (
            O => \N__13727\,
            I => \N__13724\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__13724\,
            I => \uart_pc_sync.aux_0__0_Z0Z_0\
        );

    \I__2062\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13718\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__13718\,
            I => \uart_pc_sync.aux_1__0_Z0Z_0\
        );

    \I__2060\ : InMux
    port map (
            O => \N__13715\,
            I => \N__13712\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__13712\,
            I => \uart_pc_sync.aux_2__0_Z0Z_0\
        );

    \I__2058\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__13706\,
            I => \N__13703\
        );

    \I__2056\ : Odrv12
    port map (
            O => \N__13703\,
            I => \uart_pc_sync.aux_3__0_Z0Z_0\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__13700\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__13697\,
            I => \uart_frame_decoder.state_1_RNO_3Z0Z_0_cascade_\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__13694\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\
        );

    \I__2052\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13688\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__13688\,
            I => \N__13685\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__13685\,
            I => \N__13682\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__13682\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__2048\ : InMux
    port map (
            O => \N__13679\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13\
        );

    \I__2047\ : InMux
    port map (
            O => \N__13676\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_14\
        );

    \I__2046\ : InMux
    port map (
            O => \N__13673\,
            I => \bfn_7_28_0_\
        );

    \I__2045\ : InMux
    port map (
            O => \N__13670\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_16\
        );

    \I__2044\ : InMux
    port map (
            O => \N__13667\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_17\
        );

    \I__2043\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__13661\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_17\
        );

    \I__2041\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__13655\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_16\
        );

    \I__2039\ : InMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__13649\,
            I => \N__13646\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__13646\,
            I => uart_input_pc_c
        );

    \I__2036\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__2034\ : Odrv12
    port map (
            O => \N__13637\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__13634\,
            I => \N__13631\
        );

    \I__2032\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13628\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__13628\,
            I => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__13625\,
            I => \N__13622\
        );

    \I__2029\ : InMux
    port map (
            O => \N__13622\,
            I => \N__13619\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__13619\,
            I => \ppm_encoder_1.un1_init_pulses_11_6\
        );

    \I__2027\ : InMux
    port map (
            O => \N__13616\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_5\
        );

    \I__2026\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13610\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__13610\,
            I => \N__13607\
        );

    \I__2024\ : Odrv12
    port map (
            O => \N__13607\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_7\
        );

    \I__2023\ : InMux
    port map (
            O => \N__13604\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_6\
        );

    \I__2022\ : InMux
    port map (
            O => \N__13601\,
            I => \bfn_7_27_0_\
        );

    \I__2021\ : InMux
    port map (
            O => \N__13598\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_8\
        );

    \I__2020\ : InMux
    port map (
            O => \N__13595\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_9\
        );

    \I__2019\ : InMux
    port map (
            O => \N__13592\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_10\
        );

    \I__2018\ : InMux
    port map (
            O => \N__13589\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_11\
        );

    \I__2017\ : InMux
    port map (
            O => \N__13586\,
            I => \N__13583\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__2015\ : Odrv12
    port map (
            O => \N__13580\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__13577\,
            I => \N__13574\
        );

    \I__2013\ : InMux
    port map (
            O => \N__13574\,
            I => \N__13571\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__13571\,
            I => \N__13568\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__13568\,
            I => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\
        );

    \I__2010\ : InMux
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__13559\,
            I => \ppm_encoder_1.un1_init_pulses_11_13\
        );

    \I__2007\ : InMux
    port map (
            O => \N__13556\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_12\
        );

    \I__2006\ : InMux
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__13550\,
            I => \N__13547\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__13547\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\
        );

    \I__2003\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__13541\,
            I => \N__13538\
        );

    \I__2001\ : Odrv12
    port map (
            O => \N__13538\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_1\
        );

    \I__2000\ : InMux
    port map (
            O => \N__13535\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_0\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__13532\,
            I => \N__13529\
        );

    \I__1998\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13526\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__13526\,
            I => \N__13523\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__13523\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\
        );

    \I__1995\ : InMux
    port map (
            O => \N__13520\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_1\
        );

    \I__1994\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13514\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__13514\,
            I => \N__13511\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__13511\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_3\
        );

    \I__1991\ : InMux
    port map (
            O => \N__13508\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_2\
        );

    \I__1990\ : InMux
    port map (
            O => \N__13505\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_3\
        );

    \I__1989\ : InMux
    port map (
            O => \N__13502\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_4\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__13499\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\
        );

    \I__1987\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13487\
        );

    \I__1986\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13487\
        );

    \I__1985\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13487\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__13487\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__13484\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__13481\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__13478\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\
        );

    \I__1980\ : CEMux
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__13466\,
            I => \uart_frame_decoder.source_offset1data_1_sqmuxa_0\
        );

    \I__1976\ : InMux
    port map (
            O => \N__13463\,
            I => \uart_frame_decoder.un1_WDT_cry_10\
        );

    \I__1975\ : InMux
    port map (
            O => \N__13460\,
            I => \uart_frame_decoder.un1_WDT_cry_11\
        );

    \I__1974\ : InMux
    port map (
            O => \N__13457\,
            I => \uart_frame_decoder.un1_WDT_cry_12\
        );

    \I__1973\ : InMux
    port map (
            O => \N__13454\,
            I => \uart_frame_decoder.un1_WDT_cry_13\
        );

    \I__1972\ : InMux
    port map (
            O => \N__13451\,
            I => \uart_frame_decoder.un1_WDT_cry_14\
        );

    \I__1971\ : InMux
    port map (
            O => \N__13448\,
            I => \uart_frame_decoder.un1_WDT_cry_1\
        );

    \I__1970\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__13442\,
            I => \uart_frame_decoder.WDTZ0Z_3\
        );

    \I__1968\ : InMux
    port map (
            O => \N__13439\,
            I => \uart_frame_decoder.un1_WDT_cry_2\
        );

    \I__1967\ : InMux
    port map (
            O => \N__13436\,
            I => \uart_frame_decoder.un1_WDT_cry_3\
        );

    \I__1966\ : InMux
    port map (
            O => \N__13433\,
            I => \uart_frame_decoder.un1_WDT_cry_4\
        );

    \I__1965\ : InMux
    port map (
            O => \N__13430\,
            I => \uart_frame_decoder.un1_WDT_cry_5\
        );

    \I__1964\ : InMux
    port map (
            O => \N__13427\,
            I => \uart_frame_decoder.un1_WDT_cry_6\
        );

    \I__1963\ : InMux
    port map (
            O => \N__13424\,
            I => \bfn_7_16_0_\
        );

    \I__1962\ : InMux
    port map (
            O => \N__13421\,
            I => \uart_frame_decoder.un1_WDT_cry_8\
        );

    \I__1961\ : InMux
    port map (
            O => \N__13418\,
            I => \uart_frame_decoder.un1_WDT_cry_9\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__13415\,
            I => \uart_frame_decoder.source_offset2data_1_sqmuxa_cascade_\
        );

    \I__1959\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13409\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__13409\,
            I => \uart_frame_decoder.WDTZ0Z_0\
        );

    \I__1957\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13403\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__13403\,
            I => \uart_frame_decoder.WDTZ0Z_1\
        );

    \I__1955\ : InMux
    port map (
            O => \N__13400\,
            I => \uart_frame_decoder.un1_WDT_cry_0\
        );

    \I__1954\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13394\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__13394\,
            I => \uart_frame_decoder.WDTZ0Z_2\
        );

    \I__1952\ : InMux
    port map (
            O => \N__13391\,
            I => \N__13388\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__13388\,
            I => uart_input_drone_c
        );

    \I__1950\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13382\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__13382\,
            I => \uart_drone_sync.aux_0__0__0_0\
        );

    \I__1948\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13376\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__1946\ : Odrv4
    port map (
            O => \N__13373\,
            I => \uart_drone_sync.aux_1__0__0_0\
        );

    \I__1945\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13367\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__13367\,
            I => \N__13364\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__13364\,
            I => \N__13360\
        );

    \I__1942\ : InMux
    port map (
            O => \N__13363\,
            I => \N__13357\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__13360\,
            I => \uart_pc.data_AuxZ0Z_1\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__13357\,
            I => \uart_pc.data_AuxZ0Z_1\
        );

    \I__1939\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13349\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__13349\,
            I => \N__13345\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__13348\,
            I => \N__13342\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__13345\,
            I => \N__13339\
        );

    \I__1935\ : InMux
    port map (
            O => \N__13342\,
            I => \N__13336\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__13339\,
            I => \uart_pc.data_AuxZ0Z_0\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__13336\,
            I => \uart_pc.data_AuxZ0Z_0\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__1931\ : InMux
    port map (
            O => \N__13328\,
            I => \N__13324\
        );

    \I__1930\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13321\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__13324\,
            I => \N__13318\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13315\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__13318\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__13315\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__1925\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13306\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__13309\,
            I => \N__13303\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__13306\,
            I => \N__13300\
        );

    \I__1922\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13297\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__13300\,
            I => \uart_pc.data_AuxZ0Z_2\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__13297\,
            I => \uart_pc.data_AuxZ0Z_2\
        );

    \I__1919\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13289\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__13289\,
            I => \N__13285\
        );

    \I__1917\ : InMux
    port map (
            O => \N__13288\,
            I => \N__13282\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__13285\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__13282\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__1914\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__13274\,
            I => \N__13270\
        );

    \I__1912\ : InMux
    port map (
            O => \N__13273\,
            I => \N__13267\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__13270\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__13267\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__1909\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13258\
        );

    \I__1908\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13255\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__13258\,
            I => \N__13250\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__13255\,
            I => \N__13250\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__13250\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__13247\,
            I => \uart_pc.N_143_cascade_\
        );

    \I__1903\ : InMux
    port map (
            O => \N__13244\,
            I => \N__13241\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__13241\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_1\
        );

    \I__1901\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13234\
        );

    \I__1900\ : InMux
    port map (
            O => \N__13237\,
            I => \N__13231\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__13234\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__13231\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__13226\,
            I => \N__13220\
        );

    \I__1896\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13215\
        );

    \I__1895\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13215\
        );

    \I__1894\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13210\
        );

    \I__1893\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13210\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__13215\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__13210\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__13205\,
            I => \N__13202\
        );

    \I__1889\ : InMux
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__13199\,
            I => \uart_pc.un1_state_2_0_a3_0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__13196\,
            I => \uart_pc.un4_timer_Count_1_cry_1\
        );

    \I__1886\ : InMux
    port map (
            O => \N__13193\,
            I => \uart_pc.un4_timer_Count_1_cry_2\
        );

    \I__1885\ : InMux
    port map (
            O => \N__13190\,
            I => \uart_pc.un4_timer_Count_1_cry_3\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_4_cascade_\
        );

    \I__1883\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13178\
        );

    \I__1882\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13175\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__13182\,
            I => \N__13170\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__13181\,
            I => \N__13166\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__13178\,
            I => \N__13160\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13160\
        );

    \I__1877\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13156\
        );

    \I__1876\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13147\
        );

    \I__1875\ : InMux
    port map (
            O => \N__13170\,
            I => \N__13147\
        );

    \I__1874\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13147\
        );

    \I__1873\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13147\
        );

    \I__1872\ : InMux
    port map (
            O => \N__13165\,
            I => \N__13144\
        );

    \I__1871\ : Span4Mux_v
    port map (
            O => \N__13160\,
            I => \N__13141\
        );

    \I__1870\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13138\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__13156\,
            I => \N__13133\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__13147\,
            I => \N__13133\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__13144\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__13141\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__13138\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__1864\ : Odrv12
    port map (
            O => \N__13133\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__1863\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__13121\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_2\
        );

    \I__1861\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13113\
        );

    \I__1860\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13110\
        );

    \I__1859\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13107\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__13113\,
            I => \N__13104\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__13110\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__13107\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__13104\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__1854\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13094\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__13094\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_3\
        );

    \I__1852\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13084\
        );

    \I__1851\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13081\
        );

    \I__1850\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13076\
        );

    \I__1849\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13076\
        );

    \I__1848\ : InMux
    port map (
            O => \N__13087\,
            I => \N__13073\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__13084\,
            I => \uart_pc.N_143\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__13081\,
            I => \uart_pc.N_143\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__13076\,
            I => \uart_pc.N_143\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__13073\,
            I => \uart_pc.N_143\
        );

    \I__1843\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13055\
        );

    \I__1842\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13055\
        );

    \I__1841\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13055\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__13055\,
            I => \N__13050\
        );

    \I__1839\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13045\
        );

    \I__1838\ : InMux
    port map (
            O => \N__13053\,
            I => \N__13045\
        );

    \I__1837\ : Odrv12
    port map (
            O => \N__13050\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__13045\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__1835\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13036\
        );

    \I__1834\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13027\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__13036\,
            I => \N__13024\
        );

    \I__1832\ : InMux
    port map (
            O => \N__13035\,
            I => \N__13015\
        );

    \I__1831\ : InMux
    port map (
            O => \N__13034\,
            I => \N__13015\
        );

    \I__1830\ : InMux
    port map (
            O => \N__13033\,
            I => \N__13015\
        );

    \I__1829\ : InMux
    port map (
            O => \N__13032\,
            I => \N__13015\
        );

    \I__1828\ : InMux
    port map (
            O => \N__13031\,
            I => \N__13012\
        );

    \I__1827\ : InMux
    port map (
            O => \N__13030\,
            I => \N__13009\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__13027\,
            I => \N__13006\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__13024\,
            I => \N__13001\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__13015\,
            I => \N__13001\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__13012\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__13009\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__1821\ : Odrv12
    port map (
            O => \N__13006\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__13001\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__12992\,
            I => \uart_pc.N_145_cascade_\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__12989\,
            I => \N__12984\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__12988\,
            I => \N__12981\
        );

    \I__1816\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12977\
        );

    \I__1815\ : InMux
    port map (
            O => \N__12984\,
            I => \N__12972\
        );

    \I__1814\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12972\
        );

    \I__1813\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12969\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__12977\,
            I => \N__12964\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__12972\,
            I => \N__12964\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__12969\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__12964\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__1808\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12954\
        );

    \I__1807\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12951\
        );

    \I__1806\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12947\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__12954\,
            I => \N__12944\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__12951\,
            I => \N__12941\
        );

    \I__1803\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12938\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__12947\,
            I => \uart_pc.N_152\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__12944\,
            I => \uart_pc.N_152\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__12941\,
            I => \uart_pc.N_152\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__12938\,
            I => \uart_pc.N_152\
        );

    \I__1798\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12923\
        );

    \I__1797\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12923\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__12923\,
            I => \uart_pc.N_144_1\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__12920\,
            I => \N__12913\
        );

    \I__1794\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12910\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__12918\,
            I => \N__12906\
        );

    \I__1792\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12901\
        );

    \I__1791\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12896\
        );

    \I__1790\ : InMux
    port map (
            O => \N__12913\,
            I => \N__12896\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__12910\,
            I => \N__12893\
        );

    \I__1788\ : InMux
    port map (
            O => \N__12909\,
            I => \N__12890\
        );

    \I__1787\ : InMux
    port map (
            O => \N__12906\,
            I => \N__12883\
        );

    \I__1786\ : InMux
    port map (
            O => \N__12905\,
            I => \N__12883\
        );

    \I__1785\ : InMux
    port map (
            O => \N__12904\,
            I => \N__12883\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__12901\,
            I => \N__12878\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__12896\,
            I => \N__12878\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__12893\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__12890\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__12883\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__12878\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__1778\ : InMux
    port map (
            O => \N__12869\,
            I => \N__12859\
        );

    \I__1777\ : InMux
    port map (
            O => \N__12868\,
            I => \N__12844\
        );

    \I__1776\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12844\
        );

    \I__1775\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12844\
        );

    \I__1774\ : InMux
    port map (
            O => \N__12865\,
            I => \N__12844\
        );

    \I__1773\ : InMux
    port map (
            O => \N__12864\,
            I => \N__12844\
        );

    \I__1772\ : InMux
    port map (
            O => \N__12863\,
            I => \N__12844\
        );

    \I__1771\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12844\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__12859\,
            I => \N__12839\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__12844\,
            I => \N__12839\
        );

    \I__1768\ : Odrv12
    port map (
            O => \N__12839\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__1766\ : InMux
    port map (
            O => \N__12833\,
            I => \N__12830\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__12830\,
            I => \N__12826\
        );

    \I__1764\ : InMux
    port map (
            O => \N__12829\,
            I => \N__12823\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__12826\,
            I => \uart_pc.N_126_li\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__12823\,
            I => \uart_pc.N_126_li\
        );

    \I__1761\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12813\
        );

    \I__1760\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12808\
        );

    \I__1759\ : InMux
    port map (
            O => \N__12816\,
            I => \N__12804\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12801\
        );

    \I__1757\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12796\
        );

    \I__1756\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12796\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__12808\,
            I => \N__12793\
        );

    \I__1754\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12790\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__12804\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__1752\ : Odrv12
    port map (
            O => \N__12801\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__12796\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__12793\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__12790\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__12779\,
            I => \uart_pc.N_126_li_cascade_\
        );

    \I__1747\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__12773\,
            I => \uart_pc.data_Auxce_0_0_0\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__12770\,
            I => \N__12765\
        );

    \I__1744\ : InMux
    port map (
            O => \N__12769\,
            I => \N__12760\
        );

    \I__1743\ : InMux
    port map (
            O => \N__12768\,
            I => \N__12760\
        );

    \I__1742\ : InMux
    port map (
            O => \N__12765\,
            I => \N__12751\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__12760\,
            I => \N__12748\
        );

    \I__1740\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12737\
        );

    \I__1739\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12737\
        );

    \I__1738\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12737\
        );

    \I__1737\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12737\
        );

    \I__1736\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12737\
        );

    \I__1735\ : InMux
    port map (
            O => \N__12754\,
            I => \N__12734\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__12751\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__12748\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__12737\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__12734\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__12725\,
            I => \uart_pc.un1_state_4_0_cascade_\
        );

    \I__1729\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__12719\,
            I => \uart_pc.CO0\
        );

    \I__1727\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12712\
        );

    \I__1726\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12709\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__12712\,
            I => \uart_pc.un1_state_7_0\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__12709\,
            I => \uart_pc.un1_state_7_0\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__12704\,
            I => \N__12696\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__12703\,
            I => \N__12693\
        );

    \I__1721\ : InMux
    port map (
            O => \N__12702\,
            I => \N__12685\
        );

    \I__1720\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12685\
        );

    \I__1719\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12682\
        );

    \I__1718\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12671\
        );

    \I__1717\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12671\
        );

    \I__1716\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12671\
        );

    \I__1715\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12671\
        );

    \I__1714\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12671\
        );

    \I__1713\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12667\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__12685\,
            I => \N__12664\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__12682\,
            I => \N__12659\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__12671\,
            I => \N__12659\
        );

    \I__1709\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12656\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__12667\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__1707\ : Odrv12
    port map (
            O => \N__12664\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__12659\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__12656\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__12647\,
            I => \N__12643\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__12646\,
            I => \N__12640\
        );

    \I__1702\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12635\
        );

    \I__1701\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12635\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__12635\,
            I => \N__12631\
        );

    \I__1699\ : InMux
    port map (
            O => \N__12634\,
            I => \N__12628\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__12631\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__12628\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__1696\ : InMux
    port map (
            O => \N__12623\,
            I => \N__12610\
        );

    \I__1695\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12610\
        );

    \I__1694\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12599\
        );

    \I__1693\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12599\
        );

    \I__1692\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12599\
        );

    \I__1691\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12599\
        );

    \I__1690\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12599\
        );

    \I__1689\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12592\
        );

    \I__1688\ : InMux
    port map (
            O => \N__12615\,
            I => \N__12592\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__12610\,
            I => \N__12587\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__12599\,
            I => \N__12587\
        );

    \I__1685\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12582\
        );

    \I__1684\ : InMux
    port map (
            O => \N__12597\,
            I => \N__12582\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__12592\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__12587\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__12582\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__1680\ : SRMux
    port map (
            O => \N__12575\,
            I => \N__12571\
        );

    \I__1679\ : SRMux
    port map (
            O => \N__12574\,
            I => \N__12568\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__12571\,
            I => \N__12565\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__12568\,
            I => \N__12562\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__12565\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__12562\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__1674\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12554\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__12554\,
            I => \uart_pc.data_Auxce_0_0_2\
        );

    \I__1672\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12548\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__12548\,
            I => \uart_pc.data_Auxce_0_3\
        );

    \I__1670\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12542\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__12542\,
            I => \uart_pc.data_Auxce_0_5\
        );

    \I__1668\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__12536\,
            I => \N__12533\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__12533\,
            I => \uart_pc.data_Auxce_0_0_4\
        );

    \I__1665\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12524\
        );

    \I__1664\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12519\
        );

    \I__1663\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12514\
        );

    \I__1662\ : InMux
    port map (
            O => \N__12527\,
            I => \N__12514\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__12524\,
            I => \N__12511\
        );

    \I__1660\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12508\
        );

    \I__1659\ : InMux
    port map (
            O => \N__12522\,
            I => \N__12505\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__12519\,
            I => \N__12500\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__12514\,
            I => \N__12500\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__12511\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__12508\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__12505\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__12500\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__12491\,
            I => \N__12488\
        );

    \I__1651\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12485\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__12485\,
            I => \N__12481\
        );

    \I__1649\ : InMux
    port map (
            O => \N__12484\,
            I => \N__12478\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__12481\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__12478\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__1645\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12464\
        );

    \I__1644\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12461\
        );

    \I__1643\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12456\
        );

    \I__1642\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12456\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__12464\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__12461\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__12456\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__1638\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12436\
        );

    \I__1637\ : InMux
    port map (
            O => \N__12448\,
            I => \N__12436\
        );

    \I__1636\ : InMux
    port map (
            O => \N__12447\,
            I => \N__12431\
        );

    \I__1635\ : InMux
    port map (
            O => \N__12446\,
            I => \N__12431\
        );

    \I__1634\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12424\
        );

    \I__1633\ : InMux
    port map (
            O => \N__12444\,
            I => \N__12424\
        );

    \I__1632\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12424\
        );

    \I__1631\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12417\
        );

    \I__1630\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12417\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__12436\,
            I => \N__12414\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__12431\,
            I => \N__12411\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__12424\,
            I => \N__12408\
        );

    \I__1626\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12403\
        );

    \I__1625\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12403\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__12417\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__12414\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__1622\ : Odrv12
    port map (
            O => \N__12411\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__12408\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__12403\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__1619\ : InMux
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__12389\,
            I => \uart_drone.CO0\
        );

    \I__1617\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12382\
        );

    \I__1616\ : InMux
    port map (
            O => \N__12385\,
            I => \N__12379\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__12382\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__12379\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__12374\,
            I => \N__12367\
        );

    \I__1612\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12358\
        );

    \I__1611\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12358\
        );

    \I__1610\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12353\
        );

    \I__1609\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12353\
        );

    \I__1608\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12346\
        );

    \I__1607\ : InMux
    port map (
            O => \N__12366\,
            I => \N__12346\
        );

    \I__1606\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12346\
        );

    \I__1605\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12342\
        );

    \I__1604\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12339\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__12358\,
            I => \N__12336\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__12353\,
            I => \N__12333\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__12346\,
            I => \N__12330\
        );

    \I__1600\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12327\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__12342\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__12339\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__12336\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__12333\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__12330\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__12327\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__1593\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12304\
        );

    \I__1592\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12304\
        );

    \I__1591\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12297\
        );

    \I__1590\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12297\
        );

    \I__1589\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12297\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__12309\,
            I => \N__12292\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__12304\,
            I => \N__12287\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__12297\,
            I => \N__12287\
        );

    \I__1585\ : InMux
    port map (
            O => \N__12296\,
            I => \N__12282\
        );

    \I__1584\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12282\
        );

    \I__1583\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12278\
        );

    \I__1582\ : Sp12to4
    port map (
            O => \N__12287\,
            I => \N__12273\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__12282\,
            I => \N__12273\
        );

    \I__1580\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12270\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__12278\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__12273\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__12270\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__1576\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12260\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__12260\,
            I => \uart_drone_sync.aux_2__0__0_0\
        );

    \I__1574\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12254\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__12254\,
            I => \uart_pc.data_Auxce_0_6\
        );

    \I__1572\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12248\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__12248\,
            I => \uart_pc.data_Auxce_0_1\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__12245\,
            I => \N__12242\
        );

    \I__1569\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12233\
        );

    \I__1568\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12233\
        );

    \I__1567\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12230\
        );

    \I__1566\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12225\
        );

    \I__1565\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12225\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__12233\,
            I => \uart_drone.N_143\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__12230\,
            I => \uart_drone.N_143\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__12225\,
            I => \uart_drone.N_143\
        );

    \I__1561\ : InMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__12215\,
            I => \uart_drone.N_144_1\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__12212\,
            I => \uart_drone.N_144_1_cascade_\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__12209\,
            I => \N__12204\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__12208\,
            I => \N__12201\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__12207\,
            I => \N__12197\
        );

    \I__1555\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12192\
        );

    \I__1554\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12192\
        );

    \I__1553\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12187\
        );

    \I__1552\ : InMux
    port map (
            O => \N__12197\,
            I => \N__12187\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__12192\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__12187\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__1549\ : InMux
    port map (
            O => \N__12182\,
            I => \N__12179\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__12179\,
            I => \uart_drone.N_145\
        );

    \I__1547\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12166\
        );

    \I__1546\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12163\
        );

    \I__1545\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12160\
        );

    \I__1544\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12153\
        );

    \I__1543\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12153\
        );

    \I__1542\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12153\
        );

    \I__1541\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12148\
        );

    \I__1540\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12148\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__12166\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__12163\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__12160\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__12153\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__12148\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__12137\,
            I => \N__12130\
        );

    \I__1533\ : InMux
    port map (
            O => \N__12136\,
            I => \N__12126\
        );

    \I__1532\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12123\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__12134\,
            I => \N__12119\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__12133\,
            I => \N__12115\
        );

    \I__1529\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12112\
        );

    \I__1528\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12109\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__12126\,
            I => \N__12104\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__12123\,
            I => \N__12104\
        );

    \I__1525\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12101\
        );

    \I__1524\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12094\
        );

    \I__1523\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12094\
        );

    \I__1522\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12094\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__12112\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__12109\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__12104\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__12101\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__12094\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__1516\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12079\
        );

    \I__1515\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12074\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__12079\,
            I => \N__12071\
        );

    \I__1513\ : InMux
    port map (
            O => \N__12078\,
            I => \N__12068\
        );

    \I__1512\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12065\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__12074\,
            I => \uart_drone.N_152\
        );

    \I__1510\ : Odrv12
    port map (
            O => \N__12071\,
            I => \uart_drone.N_152\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__12068\,
            I => \uart_drone.N_152\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__12065\,
            I => \uart_drone.N_152\
        );

    \I__1507\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12052\
        );

    \I__1506\ : IoInMux
    port map (
            O => \N__12055\,
            I => \N__12047\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__12052\,
            I => \N__12044\
        );

    \I__1504\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12036\
        );

    \I__1503\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12033\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__12047\,
            I => \N__12030\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__12044\,
            I => \N__12027\
        );

    \I__1500\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12018\
        );

    \I__1499\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12018\
        );

    \I__1498\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12018\
        );

    \I__1497\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12018\
        );

    \I__1496\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12010\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__12036\,
            I => \N__12007\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__12033\,
            I => \N__12004\
        );

    \I__1493\ : IoSpan4Mux
    port map (
            O => \N__12030\,
            I => \N__12001\
        );

    \I__1492\ : Sp12to4
    port map (
            O => \N__12027\,
            I => \N__11998\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__12018\,
            I => \N__11995\
        );

    \I__1490\ : InMux
    port map (
            O => \N__12017\,
            I => \N__11990\
        );

    \I__1489\ : InMux
    port map (
            O => \N__12016\,
            I => \N__11990\
        );

    \I__1488\ : InMux
    port map (
            O => \N__12015\,
            I => \N__11987\
        );

    \I__1487\ : InMux
    port map (
            O => \N__12014\,
            I => \N__11984\
        );

    \I__1486\ : InMux
    port map (
            O => \N__12013\,
            I => \N__11981\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__12010\,
            I => \N__11974\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__12007\,
            I => \N__11974\
        );

    \I__1483\ : Span4Mux_h
    port map (
            O => \N__12004\,
            I => \N__11974\
        );

    \I__1482\ : Span4Mux_s1_v
    port map (
            O => \N__12001\,
            I => \N__11971\
        );

    \I__1481\ : Span12Mux_h
    port map (
            O => \N__11998\,
            I => \N__11958\
        );

    \I__1480\ : Sp12to4
    port map (
            O => \N__11995\,
            I => \N__11958\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__11990\,
            I => \N__11958\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__11987\,
            I => \N__11958\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__11984\,
            I => \N__11958\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__11981\,
            I => \N__11958\
        );

    \I__1475\ : Span4Mux_v
    port map (
            O => \N__11974\,
            I => \N__11955\
        );

    \I__1474\ : Span4Mux_h
    port map (
            O => \N__11971\,
            I => \N__11952\
        );

    \I__1473\ : Span12Mux_v
    port map (
            O => \N__11958\,
            I => \N__11947\
        );

    \I__1472\ : Sp12to4
    port map (
            O => \N__11955\,
            I => \N__11947\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__11952\,
            I => uart_input_debug_c
        );

    \I__1470\ : Odrv12
    port map (
            O => \N__11947\,
            I => uart_input_debug_c
        );

    \I__1469\ : InMux
    port map (
            O => \N__11942\,
            I => \N__11934\
        );

    \I__1468\ : InMux
    port map (
            O => \N__11941\,
            I => \N__11929\
        );

    \I__1467\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11929\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__11939\,
            I => \N__11923\
        );

    \I__1465\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11920\
        );

    \I__1464\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11917\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__11934\,
            I => \N__11912\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__11929\,
            I => \N__11912\
        );

    \I__1461\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11905\
        );

    \I__1460\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11905\
        );

    \I__1459\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11905\
        );

    \I__1458\ : InMux
    port map (
            O => \N__11923\,
            I => \N__11902\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__11920\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__11917\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__11912\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__11905\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__11902\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__1452\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11888\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__11888\,
            I => \N__11884\
        );

    \I__1450\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11881\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__11884\,
            I => \uart_drone.N_126_li\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__11881\,
            I => \uart_drone.N_126_li\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__11876\,
            I => \uart_drone.state_srsts_0_0_0_cascade_\
        );

    \I__1446\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__11870\,
            I => \uart_drone.data_Auxce_0_5\
        );

    \I__1444\ : InMux
    port map (
            O => \N__11867\,
            I => \N__11861\
        );

    \I__1443\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11861\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__11861\,
            I => \N__11852\
        );

    \I__1441\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11847\
        );

    \I__1440\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11847\
        );

    \I__1439\ : InMux
    port map (
            O => \N__11858\,
            I => \N__11838\
        );

    \I__1438\ : InMux
    port map (
            O => \N__11857\,
            I => \N__11838\
        );

    \I__1437\ : InMux
    port map (
            O => \N__11856\,
            I => \N__11838\
        );

    \I__1436\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11838\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__11852\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__11847\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__11838\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__11831\,
            I => \N__11827\
        );

    \I__1431\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11824\
        );

    \I__1430\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11821\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__11824\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__11821\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__1427\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11813\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__11813\,
            I => \uart_drone.data_Auxce_0_6\
        );

    \I__1425\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11807\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__11807\,
            I => \N__11804\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__11804\,
            I => \uart_drone.data_Auxce_0_0_2\
        );

    \I__1422\ : SRMux
    port map (
            O => \N__11801\,
            I => \N__11797\
        );

    \I__1421\ : SRMux
    port map (
            O => \N__11800\,
            I => \N__11794\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__11797\,
            I => \N__11790\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__11794\,
            I => \N__11787\
        );

    \I__1418\ : SRMux
    port map (
            O => \N__11793\,
            I => \N__11784\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__11790\,
            I => \N__11777\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__11787\,
            I => \N__11777\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__11784\,
            I => \N__11777\
        );

    \I__1414\ : Span4Mux_h
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__11774\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__1412\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__11768\,
            I => \uart_drone.timer_Count_RNO_0_0_4\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__11765\,
            I => \uart_drone.N_143_cascade_\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__11762\,
            I => \N__11756\
        );

    \I__1408\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11751\
        );

    \I__1407\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11751\
        );

    \I__1406\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11746\
        );

    \I__1405\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11746\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__11751\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__11746\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__11741\,
            I => \N__11736\
        );

    \I__1401\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11731\
        );

    \I__1400\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11726\
        );

    \I__1399\ : InMux
    port map (
            O => \N__11736\,
            I => \N__11726\
        );

    \I__1398\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11721\
        );

    \I__1397\ : InMux
    port map (
            O => \N__11734\,
            I => \N__11721\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__11731\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__11726\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__11721\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__11714\,
            I => \uart_drone.timer_Count_RNO_0_0_1_cascade_\
        );

    \I__1392\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11707\
        );

    \I__1391\ : InMux
    port map (
            O => \N__11710\,
            I => \N__11704\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__11707\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__11704\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__1388\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11696\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__11696\,
            I => \uart_drone_sync.aux_3__0__0_0\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__11693\,
            I => \N__11689\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__11692\,
            I => \N__11685\
        );

    \I__1384\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11682\
        );

    \I__1383\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11679\
        );

    \I__1382\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11676\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__11682\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__11679\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__11676\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__11669\,
            I => \uart_pc.state_srsts_i_0_2_cascade_\
        );

    \I__1377\ : InMux
    port map (
            O => \N__11666\,
            I => \N__11663\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__11663\,
            I => \uart_pc.state_srsts_0_0_0\
        );

    \I__1375\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__11657\,
            I => \N__11653\
        );

    \I__1373\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11650\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__11653\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__11650\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__11645\,
            I => \N__11641\
        );

    \I__1369\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11638\
        );

    \I__1368\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11635\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__11638\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__11635\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__1365\ : InMux
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__11627\,
            I => \N__11623\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__11626\,
            I => \N__11620\
        );

    \I__1362\ : Span12Mux_v
    port map (
            O => \N__11623\,
            I => \N__11617\
        );

    \I__1361\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11614\
        );

    \I__1360\ : Odrv12
    port map (
            O => \N__11617\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__11614\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__11609\,
            I => \N__11605\
        );

    \I__1357\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11602\
        );

    \I__1356\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11599\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__11602\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__11599\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__1353\ : InMux
    port map (
            O => \N__11594\,
            I => \N__11591\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__11591\,
            I => \uart_drone.timer_Count_RNO_0_0_3\
        );

    \I__1351\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11585\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__11585\,
            I => \uart_drone.timer_Count_RNO_0_0_2\
        );

    \I__1349\ : InMux
    port map (
            O => \N__11582\,
            I => \N__11577\
        );

    \I__1348\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11572\
        );

    \I__1347\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11572\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__11577\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__11572\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__11567\,
            I => \uart_drone.state_srsts_i_0_2_cascade_\
        );

    \I__1343\ : InMux
    port map (
            O => \N__11564\,
            I => \N__11559\
        );

    \I__1342\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11556\
        );

    \I__1341\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11553\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__11559\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__11556\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__11553\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__1337\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11540\
        );

    \I__1336\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11537\
        );

    \I__1335\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11532\
        );

    \I__1334\ : InMux
    port map (
            O => \N__11543\,
            I => \N__11532\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__11540\,
            I => \N__11529\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__11537\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__11532\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__11529\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__1329\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11517\
        );

    \I__1328\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11512\
        );

    \I__1327\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11512\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__11517\,
            I => \reset_module_System.reset6_15\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__11512\,
            I => \reset_module_System.reset6_15\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__11507\,
            I => \N__11503\
        );

    \I__1323\ : InMux
    port map (
            O => \N__11506\,
            I => \N__11496\
        );

    \I__1322\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11496\
        );

    \I__1321\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11491\
        );

    \I__1320\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11491\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__11496\,
            I => \reset_module_System.reset6_14\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__11491\,
            I => \reset_module_System.reset6_14\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__11486\,
            I => \reset_module_System.count_1_1_cascade_\
        );

    \I__1316\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11475\
        );

    \I__1315\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11475\
        );

    \I__1314\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11470\
        );

    \I__1313\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11470\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__11475\,
            I => \reset_module_System.reset6_19\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__11470\,
            I => \reset_module_System.reset6_19\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__11465\,
            I => \N__11462\
        );

    \I__1309\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11458\
        );

    \I__1308\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11454\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__11458\,
            I => \N__11451\
        );

    \I__1306\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11448\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__11454\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__11451\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__11448\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__1302\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11436\
        );

    \I__1301\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11431\
        );

    \I__1300\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11431\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__11436\,
            I => \N__11428\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__11431\,
            I => \N__11425\
        );

    \I__1297\ : Odrv12
    port map (
            O => \N__11428\,
            I => \uart_drone.state_1_sqmuxa\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__11425\,
            I => \uart_drone.state_1_sqmuxa\
        );

    \I__1295\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11417\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__11417\,
            I => \uart_drone.data_Auxce_0_1\
        );

    \I__1293\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11411\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__11411\,
            I => \uart_drone.data_Auxce_0_3\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__11408\,
            I => \uart_drone.N_126_li_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11402\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__11402\,
            I => \uart_drone.un1_state_2_0_a3_0\
        );

    \I__1288\ : InMux
    port map (
            O => \N__11399\,
            I => \uart_drone.un4_timer_Count_1_cry_1\
        );

    \I__1287\ : InMux
    port map (
            O => \N__11396\,
            I => \uart_drone.un4_timer_Count_1_cry_2\
        );

    \I__1286\ : InMux
    port map (
            O => \N__11393\,
            I => \uart_drone.un4_timer_Count_1_cry_3\
        );

    \I__1285\ : InMux
    port map (
            O => \N__11390\,
            I => \N__11383\
        );

    \I__1284\ : InMux
    port map (
            O => \N__11389\,
            I => \N__11383\
        );

    \I__1283\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11380\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__11383\,
            I => \N__11376\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__11380\,
            I => \N__11373\
        );

    \I__1280\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11370\
        );

    \I__1279\ : Span4Mux_s3_h
    port map (
            O => \N__11376\,
            I => \N__11367\
        );

    \I__1278\ : Span4Mux_s3_h
    port map (
            O => \N__11373\,
            I => \N__11364\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__11370\,
            I => uart_drone_data_6
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__11367\,
            I => uart_drone_data_6
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__11364\,
            I => uart_drone_data_6
        );

    \I__1274\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11354\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__11354\,
            I => uart_drone_data_7
        );

    \I__1272\ : CEMux
    port map (
            O => \N__11351\,
            I => \N__11348\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__11348\,
            I => \N__11344\
        );

    \I__1270\ : CEMux
    port map (
            O => \N__11347\,
            I => \N__11341\
        );

    \I__1269\ : Span4Mux_v
    port map (
            O => \N__11344\,
            I => \N__11338\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__11341\,
            I => \N__11335\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__11338\,
            I => \uart_drone.state_1_sqmuxa_0\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__11335\,
            I => \uart_drone.state_1_sqmuxa_0\
        );

    \I__1265\ : SRMux
    port map (
            O => \N__11330\,
            I => \N__11327\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__11327\,
            I => \N__11323\
        );

    \I__1263\ : SRMux
    port map (
            O => \N__11326\,
            I => \N__11320\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__11323\,
            I => \N__11315\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__11320\,
            I => \N__11315\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__11315\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__11312\,
            I => \N__11308\
        );

    \I__1258\ : InMux
    port map (
            O => \N__11311\,
            I => \N__11305\
        );

    \I__1257\ : InMux
    port map (
            O => \N__11308\,
            I => \N__11302\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__11305\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__11302\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__11297\,
            I => \N__11293\
        );

    \I__1253\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__1252\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__11290\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__11287\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \N__11278\
        );

    \I__1248\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11275\
        );

    \I__1247\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11272\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__11275\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__11272\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__11267\,
            I => \uart_drone.data_Auxce_0_0_4_cascade_\
        );

    \I__1243\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11261\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__1241\ : Span4Mux_v
    port map (
            O => \N__11258\,
            I => \N__11254\
        );

    \I__1240\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11251\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__11254\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__11251\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__1237\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11243\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__11243\,
            I => \uart_drone.data_Auxce_0_0_0\
        );

    \I__1235\ : InMux
    port map (
            O => \N__11240\,
            I => \N__11237\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__11237\,
            I => \N__11234\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__11234\,
            I => \N__11229\
        );

    \I__1232\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11226\
        );

    \I__1231\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11223\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__11229\,
            I => \frame_dron_decoder_1.stateZ0Z_6\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__11226\,
            I => \frame_dron_decoder_1.stateZ0Z_6\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__11223\,
            I => \frame_dron_decoder_1.stateZ0Z_6\
        );

    \I__1227\ : IoInMux
    port map (
            O => \N__11216\,
            I => \N__11213\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__11213\,
            I => \N__11210\
        );

    \I__1225\ : Span12Mux_s1_v
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1224\ : Span12Mux_v
    port map (
            O => \N__11207\,
            I => \N__11203\
        );

    \I__1223\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11200\
        );

    \I__1222\ : Odrv12
    port map (
            O => \N__11203\,
            I => drone_frame_decoder_data_rdy_debug_c
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__11200\,
            I => drone_frame_decoder_data_rdy_debug_c
        );

    \I__1220\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11192\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__11192\,
            I => \N__11189\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__11189\,
            I => uart_drone_data_2
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__11186\,
            I => \frame_dron_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_\
        );

    \I__1216\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11179\
        );

    \I__1215\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11175\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__11179\,
            I => \N__11172\
        );

    \I__1213\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11169\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__11175\,
            I => \N__11164\
        );

    \I__1211\ : Span4Mux_s3_h
    port map (
            O => \N__11172\,
            I => \N__11164\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__11169\,
            I => \N__11161\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__11164\,
            I => \frame_dron_decoder_1.N_255\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__11161\,
            I => \frame_dron_decoder_1.N_255\
        );

    \I__1207\ : IoInMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__1205\ : Span4Mux_s1_v
    port map (
            O => \N__11150\,
            I => \N__11145\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__11149\,
            I => \N__11142\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__11148\,
            I => \N__11138\
        );

    \I__1202\ : Sp12to4
    port map (
            O => \N__11145\,
            I => \N__11131\
        );

    \I__1201\ : InMux
    port map (
            O => \N__11142\,
            I => \N__11122\
        );

    \I__1200\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11122\
        );

    \I__1199\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11122\
        );

    \I__1198\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11122\
        );

    \I__1197\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11118\
        );

    \I__1196\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11115\
        );

    \I__1195\ : InMux
    port map (
            O => \N__11134\,
            I => \N__11112\
        );

    \I__1194\ : Span12Mux_h
    port map (
            O => \N__11131\,
            I => \N__11109\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__11122\,
            I => \N__11106\
        );

    \I__1192\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11103\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__11118\,
            I => \N__11100\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__11115\,
            I => \N__11095\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__11112\,
            I => \N__11095\
        );

    \I__1188\ : Span12Mux_v
    port map (
            O => \N__11109\,
            I => \N__11090\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__11106\,
            I => \N__11081\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__11103\,
            I => \N__11081\
        );

    \I__1185\ : Span4Mux_s2_h
    port map (
            O => \N__11100\,
            I => \N__11081\
        );

    \I__1184\ : Span4Mux_v
    port map (
            O => \N__11095\,
            I => \N__11081\
        );

    \I__1183\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11076\
        );

    \I__1182\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11076\
        );

    \I__1181\ : Odrv12
    port map (
            O => \N__11090\,
            I => uart_data_rdy_debug_c
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__11081\,
            I => uart_data_rdy_debug_c
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__11076\,
            I => uart_data_rdy_debug_c
        );

    \I__1178\ : SRMux
    port map (
            O => \N__11069\,
            I => \N__11065\
        );

    \I__1177\ : SRMux
    port map (
            O => \N__11068\,
            I => \N__11062\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__11065\,
            I => \frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__11062\,
            I => \frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__1174\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__11054\,
            I => \N__11051\
        );

    \I__1172\ : Span4Mux_s3_h
    port map (
            O => \N__11051\,
            I => \N__11046\
        );

    \I__1171\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11041\
        );

    \I__1170\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11041\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__11046\,
            I => uart_drone_data_1
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__11041\,
            I => uart_drone_data_1
        );

    \I__1167\ : InMux
    port map (
            O => \N__11036\,
            I => \N__11033\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__11033\,
            I => \N__11030\
        );

    \I__1165\ : Span4Mux_s3_h
    port map (
            O => \N__11030\,
            I => \N__11025\
        );

    \I__1164\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11020\
        );

    \I__1163\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11020\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__11025\,
            I => uart_drone_data_3
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__11020\,
            I => uart_drone_data_3
        );

    \I__1160\ : InMux
    port map (
            O => \N__11015\,
            I => \N__11012\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__11012\,
            I => uart_drone_data_0
        );

    \I__1158\ : InMux
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__11006\,
            I => uart_drone_data_5
        );

    \I__1156\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10999\
        );

    \I__1155\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10996\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__10999\,
            I => \N__10993\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__10996\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__10993\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__1151\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10984\
        );

    \I__1150\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10981\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__10984\,
            I => \N__10978\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__10981\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__10978\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__1146\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10969\
        );

    \I__1145\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10966\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__10969\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__10966\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__1142\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10957\
        );

    \I__1141\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10954\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__10957\,
            I => \N__10951\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__10954\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__10951\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__10946\,
            I => \reset_module_System.reset6_3_cascade_\
        );

    \I__1136\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10940\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__10940\,
            I => \reset_module_System.reset6_13\
        );

    \I__1134\ : InMux
    port map (
            O => \N__10937\,
            I => \N__10934\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10930\
        );

    \I__1132\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10927\
        );

    \I__1131\ : Odrv12
    port map (
            O => \N__10930\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__10927\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__10922\,
            I => \reset_module_System.reset6_17_cascade_\
        );

    \I__1128\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10916\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__10916\,
            I => \reset_module_System.reset6_11\
        );

    \I__1126\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10910\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__10910\,
            I => \N__10906\
        );

    \I__1124\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10903\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__10906\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__10903\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__1121\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__10895\,
            I => \N__10891\
        );

    \I__1119\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10888\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__10891\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__10888\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__1116\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10879\
        );

    \I__1115\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10876\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__10879\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__10876\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__10871\,
            I => \reset_module_System.reset6_15_cascade_\
        );

    \I__1111\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__10862\,
            I => \reset_module_System.count_1_2\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__10859\,
            I => \N__10855\
        );

    \I__1107\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10852\
        );

    \I__1106\ : InMux
    port map (
            O => \N__10855\,
            I => \N__10849\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__10852\,
            I => \N__10846\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__10849\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__1103\ : Odrv12
    port map (
            O => \N__10846\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__1102\ : InMux
    port map (
            O => \N__10841\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__1101\ : InMux
    port map (
            O => \N__10838\,
            I => \bfn_2_19_0_\
        );

    \I__1100\ : InMux
    port map (
            O => \N__10835\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__1099\ : InMux
    port map (
            O => \N__10832\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__1098\ : InMux
    port map (
            O => \N__10829\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__1097\ : InMux
    port map (
            O => \N__10826\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__1096\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10819\
        );

    \I__1095\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10816\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__10819\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__10816\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__1091\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10802\
        );

    \I__1090\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10802\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__10802\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__10799\,
            I => \N__10795\
        );

    \I__1087\ : InMux
    port map (
            O => \N__10798\,
            I => \N__10790\
        );

    \I__1086\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10790\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__10790\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__1084\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10783\
        );

    \I__1083\ : InMux
    port map (
            O => \N__10786\,
            I => \N__10780\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__10783\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__10780\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__1080\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10771\
        );

    \I__1079\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10768\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__10771\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__10768\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__1076\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10759\
        );

    \I__1075\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10756\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__10759\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__10756\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__1071\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10744\
        );

    \I__1070\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10741\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__10744\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__10741\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__1067\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10730\
        );

    \I__1066\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10730\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__10730\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__1064\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10723\
        );

    \I__1063\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10720\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__10723\,
            I => \N__10717\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__10720\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__10717\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__1059\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10708\
        );

    \I__1058\ : InMux
    port map (
            O => \N__10711\,
            I => \N__10705\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__10708\,
            I => \N__10702\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__10705\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__10702\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__10697\,
            I => \N__10693\
        );

    \I__1053\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10690\
        );

    \I__1052\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10687\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__10690\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__10687\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__1049\ : InMux
    port map (
            O => \N__10682\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__1048\ : InMux
    port map (
            O => \N__10679\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__1047\ : InMux
    port map (
            O => \N__10676\,
            I => \bfn_2_18_0_\
        );

    \I__1046\ : InMux
    port map (
            O => \N__10673\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__1045\ : InMux
    port map (
            O => \N__10670\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__1044\ : InMux
    port map (
            O => \N__10667\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__1043\ : InMux
    port map (
            O => \N__10664\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__1042\ : InMux
    port map (
            O => \N__10661\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__1041\ : InMux
    port map (
            O => \N__10658\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__1040\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10651\
        );

    \I__1039\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10646\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__10651\,
            I => \N__10643\
        );

    \I__1037\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10640\
        );

    \I__1036\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10637\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__10646\,
            I => \frame_dron_decoder_1.stateZ0Z_0\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__10643\,
            I => \frame_dron_decoder_1.stateZ0Z_0\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__10640\,
            I => \frame_dron_decoder_1.stateZ0Z_0\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__10637\,
            I => \frame_dron_decoder_1.stateZ0Z_0\
        );

    \I__1031\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__10625\,
            I => \frame_dron_decoder_1.state_ns_i_a2_1_2_0\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__10622\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\
        );

    \I__1028\ : InMux
    port map (
            O => \N__10619\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__1027\ : InMux
    port map (
            O => \N__10616\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__1026\ : InMux
    port map (
            O => \N__10613\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__1025\ : InMux
    port map (
            O => \N__10610\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__1024\ : InMux
    port map (
            O => \N__10607\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__1023\ : InMux
    port map (
            O => \N__10604\,
            I => \frame_dron_decoder_1.un1_WDT_cry_8\
        );

    \I__1022\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10597\
        );

    \I__1021\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10594\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__10597\,
            I => \frame_dron_decoder_1.WDTZ0Z_10\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__10594\,
            I => \frame_dron_decoder_1.WDTZ0Z_10\
        );

    \I__1018\ : InMux
    port map (
            O => \N__10589\,
            I => \frame_dron_decoder_1.un1_WDT_cry_9\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__10586\,
            I => \N__10582\
        );

    \I__1016\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10578\
        );

    \I__1015\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10573\
        );

    \I__1014\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10573\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__10578\,
            I => \frame_dron_decoder_1.WDTZ0Z_11\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__10573\,
            I => \frame_dron_decoder_1.WDTZ0Z_11\
        );

    \I__1011\ : InMux
    port map (
            O => \N__10568\,
            I => \frame_dron_decoder_1.un1_WDT_cry_10\
        );

    \I__1010\ : InMux
    port map (
            O => \N__10565\,
            I => \N__10560\
        );

    \I__1009\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10555\
        );

    \I__1008\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10555\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__10560\,
            I => \frame_dron_decoder_1.WDTZ0Z_12\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__10555\,
            I => \frame_dron_decoder_1.WDTZ0Z_12\
        );

    \I__1005\ : InMux
    port map (
            O => \N__10550\,
            I => \frame_dron_decoder_1.un1_WDT_cry_11\
        );

    \I__1004\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10543\
        );

    \I__1003\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__10543\,
            I => \frame_dron_decoder_1.WDTZ0Z_13\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__10540\,
            I => \frame_dron_decoder_1.WDTZ0Z_13\
        );

    \I__1000\ : InMux
    port map (
            O => \N__10535\,
            I => \frame_dron_decoder_1.un1_WDT_cry_12\
        );

    \I__999\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10525\
        );

    \I__998\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10525\
        );

    \I__997\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10522\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__10525\,
            I => \N__10519\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__10522\,
            I => \frame_dron_decoder_1.WDTZ0Z_14\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__10519\,
            I => \frame_dron_decoder_1.WDTZ0Z_14\
        );

    \I__993\ : InMux
    port map (
            O => \N__10514\,
            I => \frame_dron_decoder_1.un1_WDT_cry_13\
        );

    \I__992\ : InMux
    port map (
            O => \N__10511\,
            I => \frame_dron_decoder_1.un1_WDT_cry_14\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__10508\,
            I => \N__10505\
        );

    \I__990\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10498\
        );

    \I__989\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10498\
        );

    \I__988\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10495\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__10498\,
            I => \N__10492\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__10495\,
            I => \frame_dron_decoder_1.WDTZ0Z_15\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__10492\,
            I => \frame_dron_decoder_1.WDTZ0Z_15\
        );

    \I__984\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__10484\,
            I => \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__981\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10473\
        );

    \I__980\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10470\
        );

    \I__979\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10467\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__10473\,
            I => \frame_dron_decoder_1.stateZ0Z_1\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__10470\,
            I => \frame_dron_decoder_1.stateZ0Z_1\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__10467\,
            I => \frame_dron_decoder_1.stateZ0Z_1\
        );

    \I__975\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10456\
        );

    \I__974\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10449\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10446\
        );

    \I__971\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10443\
        );

    \I__970\ : Span4Mux_v
    port map (
            O => \N__10449\,
            I => \N__10436\
        );

    \I__969\ : Span4Mux_h
    port map (
            O => \N__10446\,
            I => \N__10436\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10436\
        );

    \I__967\ : Span4Mux_v
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__10433\,
            I => uart_drone_data_4
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__10430\,
            I => \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3_cascade_\
        );

    \I__964\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__10421\,
            I => \frame_dron_decoder_1.state_ns_0_a3_0_3_3\
        );

    \I__961\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__10415\,
            I => \frame_dron_decoder_1.WDTZ0Z_1\
        );

    \I__959\ : InMux
    port map (
            O => \N__10412\,
            I => \frame_dron_decoder_1.un1_WDT_cry_0\
        );

    \I__958\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__10406\,
            I => \frame_dron_decoder_1.WDTZ0Z_2\
        );

    \I__956\ : InMux
    port map (
            O => \N__10403\,
            I => \frame_dron_decoder_1.un1_WDT_cry_1\
        );

    \I__955\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__10397\,
            I => \frame_dron_decoder_1.WDTZ0Z_3\
        );

    \I__953\ : InMux
    port map (
            O => \N__10394\,
            I => \frame_dron_decoder_1.un1_WDT_cry_2\
        );

    \I__952\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10387\
        );

    \I__951\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10384\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__10387\,
            I => \frame_dron_decoder_1.WDTZ0Z_4\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__10384\,
            I => \frame_dron_decoder_1.WDTZ0Z_4\
        );

    \I__948\ : InMux
    port map (
            O => \N__10379\,
            I => \frame_dron_decoder_1.un1_WDT_cry_3\
        );

    \I__947\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10372\
        );

    \I__946\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10369\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__10372\,
            I => \frame_dron_decoder_1.WDTZ0Z_5\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__10369\,
            I => \frame_dron_decoder_1.WDTZ0Z_5\
        );

    \I__943\ : InMux
    port map (
            O => \N__10364\,
            I => \frame_dron_decoder_1.un1_WDT_cry_4\
        );

    \I__942\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10357\
        );

    \I__941\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10354\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__10357\,
            I => \frame_dron_decoder_1.WDTZ0Z_6\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__10354\,
            I => \frame_dron_decoder_1.WDTZ0Z_6\
        );

    \I__938\ : InMux
    port map (
            O => \N__10349\,
            I => \frame_dron_decoder_1.un1_WDT_cry_5\
        );

    \I__937\ : InMux
    port map (
            O => \N__10346\,
            I => \N__10342\
        );

    \I__936\ : InMux
    port map (
            O => \N__10345\,
            I => \N__10339\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__10342\,
            I => \frame_dron_decoder_1.WDTZ0Z_7\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__10339\,
            I => \frame_dron_decoder_1.WDTZ0Z_7\
        );

    \I__933\ : InMux
    port map (
            O => \N__10334\,
            I => \frame_dron_decoder_1.un1_WDT_cry_6\
        );

    \I__932\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10327\
        );

    \I__931\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10324\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__10327\,
            I => \frame_dron_decoder_1.WDTZ0Z_8\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__10324\,
            I => \frame_dron_decoder_1.WDTZ0Z_8\
        );

    \I__928\ : InMux
    port map (
            O => \N__10319\,
            I => \bfn_2_15_0_\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__10316\,
            I => \N__10312\
        );

    \I__926\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10309\
        );

    \I__925\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10306\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__10309\,
            I => \frame_dron_decoder_1.WDTZ0Z_9\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__10306\,
            I => \frame_dron_decoder_1.WDTZ0Z_9\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__10301\,
            I => \frame_dron_decoder_1.N_229_cascade_\
        );

    \I__921\ : InMux
    port map (
            O => \N__10298\,
            I => \N__10295\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__10295\,
            I => \frame_dron_decoder_1.state_ns_i_a2_0_2_0\
        );

    \I__919\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__10289\,
            I => \frame_dron_decoder_1.N_231\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \frame_dron_decoder_1.state_ns_0_a3_0_0_1_cascade_\
        );

    \I__916\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__10280\,
            I => \frame_dron_decoder_1.state_ns_0_a3_0_3_1\
        );

    \I__914\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10273\
        );

    \I__913\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10264\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__10273\,
            I => \N__10261\
        );

    \I__911\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10256\
        );

    \I__910\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10256\
        );

    \I__909\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10247\
        );

    \I__908\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10247\
        );

    \I__907\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10247\
        );

    \I__906\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10247\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__10264\,
            I => \frame_dron_decoder_1.N_249\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__10261\,
            I => \frame_dron_decoder_1.N_249\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__10256\,
            I => \frame_dron_decoder_1.N_249\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__10247\,
            I => \frame_dron_decoder_1.N_249\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__10238\,
            I => \N__10234\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__10237\,
            I => \N__10231\
        );

    \I__899\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10228\
        );

    \I__898\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__10228\,
            I => \frame_dron_decoder_1.stateZ0Z_3\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__10225\,
            I => \frame_dron_decoder_1.stateZ0Z_3\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__10220\,
            I => \N__10216\
        );

    \I__894\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10213\
        );

    \I__893\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10210\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__10213\,
            I => \frame_dron_decoder_1.WDT10_0_i\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__10210\,
            I => \frame_dron_decoder_1.WDT10_0_i\
        );

    \I__890\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10202\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__10202\,
            I => \frame_dron_decoder_1.WDTZ0Z_0\
        );

    \I__888\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__10196\,
            I => \frame_dron_decoder_1.WDT_RNIMRG3Z0Z_4\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__10193\,
            I => \frame_dron_decoder_1.WDT_RNI6TFJ1Z0Z_10_cascade_\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__10190\,
            I => \frame_dron_decoder_1.WDT10lt14_0_cascade_\
        );

    \I__884\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__10184\,
            I => \frame_dron_decoder_1.WDT10lt14_0\
        );

    \I__882\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__10178\,
            I => \frame_dron_decoder_1.WDT10lto13_1\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__879\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__10169\,
            I => \N__10165\
        );

    \I__877\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__10165\,
            I => \frame_dron_decoder_1.stateZ0Z_7\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__10162\,
            I => \frame_dron_decoder_1.stateZ0Z_7\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__10157\,
            I => \frame_dron_decoder_1.state_ns_i_a2_0_2_0_cascade_\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__10154\,
            I => \frame_dron_decoder_1.state_ns_i_a3_1_0_cascade_\
        );

    \I__872\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10145\
        );

    \I__871\ : InMux
    port map (
            O => \N__10150\,
            I => \N__10145\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__10145\,
            I => \frame_dron_decoder_1.stateZ0Z_2\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__868\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10133\
        );

    \I__867\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10133\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__10133\,
            I => \frame_dron_decoder_1.stateZ0Z_5\
        );

    \I__865\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10124\
        );

    \I__864\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10124\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__10124\,
            I => \frame_dron_decoder_1.stateZ0Z_4\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un3_source_data_0_cry_7\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un2_source_data_0_cry_8\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un3_source_data_0_cry_7\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un2_source_data_0_cry_8\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un3_source_data_0_cry_7\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un2_source_data_0_cry_8\,
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_1.un3_source_data_0_cry_7\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_1.un2_source_data_0_cry_8\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_throttle_cry_13\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_rudder_cry_13\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_elevator_cry_13\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_11_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_aileron_cry_13\,
            carryinitout => \bfn_11_25_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_7_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            carryinitout => \bfn_7_27_0_\
        );

    \IN_MUX_bfv_7_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            carryinitout => \bfn_7_28_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_10_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_27_0_\
        );

    \IN_MUX_bfv_10_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.counter24_0_data_tmp_7\,
            carryinitout => \bfn_10_28_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_11_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_28_0_\
        );

    \IN_MUX_bfv_11_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_7\,
            carryinitout => \bfn_11_29_0_\
        );

    \IN_MUX_bfv_11_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_15\,
            carryinitout => \bfn_11_30_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \frame_dron_decoder_1.un1_WDT_cry_7\,
            carryinitout => \bfn_2_15_0_\
        );

    \reset_module_System.reset_RNITC69\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24213\,
            GLOBALBUFFEROUTPUT => reset_system_g
        );

    \pc_frame_decoder_dv_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20138\,
            GLOBALBUFFEROUTPUT => pc_frame_decoder_dv_0_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23969\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_228_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_2_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__10150\,
            in1 => \N__11137\,
            in2 => \N__10238\,
            in3 => \N__10267\,
            lcout => \frame_dron_decoder_1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25295\,
            ce => 'H',
            sr => \N__24755\
        );

    \frame_dron_decoder_1.state_5_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__10151\,
            in1 => \N__11141\,
            in2 => \N__10142\,
            in3 => \N__10269\,
            lcout => \frame_dron_decoder_1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25295\,
            ce => 'H',
            sr => \N__24755\
        );

    \frame_dron_decoder_1.state_4_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__10268\,
            in1 => \N__10138\,
            in2 => \N__11148\,
            in3 => \N__10129\,
            lcout => \frame_dron_decoder_1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25295\,
            ce => 'H',
            sr => \N__24755\
        );

    \frame_dron_decoder_1.state_7_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__10270\,
            in1 => \N__10168\,
            in2 => \N__11149\,
            in3 => \N__10130\,
            lcout => \frame_dron_decoder_1.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25295\,
            ce => 'H',
            sr => \N__24755\
        );

    \frame_dron_decoder_1.WDT_RNIMRG3_4_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10330\,
            in1 => \N__10375\,
            in2 => \N__10316\,
            in3 => \N__10390\,
            lcout => \frame_dron_decoder_1.WDT_RNIMRG3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.WDT_RNI6TFJ1_10_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__10600\,
            in1 => \N__10546\,
            in2 => \N__10586\,
            in3 => \N__10564\,
            lcout => OPEN,
            ltout => \frame_dron_decoder_1.WDT_RNI6TFJ1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.WDT_RNIA5HI2_7_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__10345\,
            in1 => \N__10199\,
            in2 => \N__10193\,
            in3 => \N__10181\,
            lcout => \frame_dron_decoder_1.WDT10lt14_0\,
            ltout => \frame_dron_decoder_1.WDT10lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.WDT_RNI3A9C3_15_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10504\,
            in2 => \N__10190\,
            in3 => \N__10531\,
            lcout => \frame_dron_decoder_1.WDT10_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.WDT_RNICPRL3_15_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010011"
        )
    port map (
            in0 => \N__10532\,
            in1 => \N__11136\,
            in2 => \N__10508\,
            in3 => \N__10187\,
            lcout => \frame_dron_decoder_1.N_249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.WDT_RNI05KQ_6_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10581\,
            in1 => \N__10563\,
            in2 => \_gnd_net_\,
            in3 => \N__10360\,
            lcout => \frame_dron_decoder_1.WDT10lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_6_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__11233\,
            in1 => \N__11135\,
            in2 => \N__10175\,
            in3 => \N__10271\,
            lcout => \frame_dron_decoder_1.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25290\,
            ce => 'H',
            sr => \N__24764\
        );

    \frame_dron_decoder_1.state_RNIOTUU_6_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11232\,
            in2 => \_gnd_net_\,
            in3 => \N__10649\,
            lcout => \frame_dron_decoder_1.state_ns_i_a2_0_2_0\,
            ltout => \frame_dron_decoder_1.state_ns_i_a2_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_RNO_3_0_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__10452\,
            in1 => \N__11389\,
            in2 => \N__10157\,
            in3 => \N__10487\,
            lcout => OPEN,
            ltout => \frame_dron_decoder_1.state_ns_i_a3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_RNO_0_0_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100000000000"
        )
    port map (
            in0 => \N__11390\,
            in1 => \N__10628\,
            in2 => \N__10154\,
            in3 => \N__11178\,
            lcout => OPEN,
            ltout => \frame_dron_decoder_1.N_229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_0_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__10272\,
            in1 => \N__10292\,
            in2 => \N__10301\,
            in3 => \N__10654\,
            lcout => \frame_dron_decoder_1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25290\,
            ce => 'H',
            sr => \N__24764\
        );

    \frame_dron_decoder_1.state_1_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__10283\,
            in1 => \N__11183\,
            in2 => \N__10481\,
            in3 => \N__10277\,
            lcout => \frame_dron_decoder_1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25285\,
            ce => 'H',
            sr => \N__24770\
        );

    \frame_dron_decoder_1.state_RNO_1_0_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10476\,
            in1 => \N__10298\,
            in2 => \_gnd_net_\,
            in3 => \N__11134\,
            lcout => \frame_dron_decoder_1.N_231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_RNO_1_1_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11388\,
            in2 => \_gnd_net_\,
            in3 => \N__11057\,
            lcout => OPEN,
            ltout => \frame_dron_decoder_1.state_ns_0_a3_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_RNO_0_1_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10460\,
            in1 => \N__10655\,
            in2 => \N__10286\,
            in3 => \N__11036\,
            lcout => \frame_dron_decoder_1.state_ns_0_a3_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_esr_4_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11264\,
            lcout => uart_drone_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25296\,
            ce => \N__11351\,
            sr => \N__11330\
        );

    \uart_drone.data_esr_2_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11630\,
            lcout => uart_drone_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25296\,
            ce => \N__11351\,
            sr => \N__11330\
        );

    \frame_dron_decoder_1.state_3_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__11182\,
            in1 => \N__10427\,
            in2 => \N__10237\,
            in3 => \N__10276\,
            lcout => \frame_dron_decoder_1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25294\,
            ce => 'H',
            sr => \N__24750\
        );

    \frame_dron_decoder_1.WDT_0_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10205\,
            in2 => \N__10220\,
            in3 => \N__10219\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_0\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_1_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__10412\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_0\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_1\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_2_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10409\,
            in2 => \_gnd_net_\,
            in3 => \N__10403\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_1\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_2\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_3_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10400\,
            in2 => \_gnd_net_\,
            in3 => \N__10394\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_2\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_3\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_4_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10391\,
            in2 => \_gnd_net_\,
            in3 => \N__10379\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_3\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_4\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_5_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10376\,
            in2 => \_gnd_net_\,
            in3 => \N__10364\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_4\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_5\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_6_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10361\,
            in2 => \_gnd_net_\,
            in3 => \N__10349\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_5\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_6\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_7_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10346\,
            in2 => \_gnd_net_\,
            in3 => \N__10334\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_6\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_7\,
            clk => \N__25291\,
            ce => 'H',
            sr => \N__11069\
        );

    \frame_dron_decoder_1.WDT_8_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10331\,
            in2 => \_gnd_net_\,
            in3 => \N__10319\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_8\,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.WDT_9_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10315\,
            in2 => \_gnd_net_\,
            in3 => \N__10604\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_8\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_9\,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.WDT_10_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10601\,
            in2 => \_gnd_net_\,
            in3 => \N__10589\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_9\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_10\,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.WDT_11_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10585\,
            in2 => \_gnd_net_\,
            in3 => \N__10568\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_10\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_11\,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.WDT_12_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10565\,
            in2 => \_gnd_net_\,
            in3 => \N__10550\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_11\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_12\,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.WDT_13_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10547\,
            in2 => \_gnd_net_\,
            in3 => \N__10535\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_12\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_13\,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.WDT_14_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10530\,
            in2 => \_gnd_net_\,
            in3 => \N__10514\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \frame_dron_decoder_1.un1_WDT_cry_13\,
            carryout => \frame_dron_decoder_1.un1_WDT_cry_14\,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.WDT_15_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10503\,
            in2 => \_gnd_net_\,
            in3 => \N__10511\,
            lcout => \frame_dron_decoder_1.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25286\,
            ce => 'H',
            sr => \N__11068\
        );

    \frame_dron_decoder_1.state_ns_0_a3_0_1_3_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11049\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11028\,
            lcout => \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3\,
            ltout => \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_RNO_0_3_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10477\,
            in1 => \N__10459\,
            in2 => \N__10430\,
            in3 => \N__11379\,
            lcout => \frame_dron_decoder_1.state_ns_0_a3_0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_RNO_2_0_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11029\,
            in1 => \N__10650\,
            in2 => \_gnd_net_\,
            in3 => \N__11050\,
            lcout => \frame_dron_decoder_1.state_ns_i_a2_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIES9Q1_2_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__12050\,
            in1 => \N__11439\,
            in2 => \_gnd_net_\,
            in3 => \N__24191\,
            lcout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\,
            ltout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIRC5U2_2_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11440\,
            in1 => \_gnd_net_\,
            in2 => \N__10622\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.state_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11546\,
            in2 => \N__11465\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10858\,
            in2 => \_gnd_net_\,
            in3 => \N__10619\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10894\,
            in2 => \_gnd_net_\,
            in3 => \N__10616\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__25277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10987\,
            in2 => \_gnd_net_\,
            in3 => \N__10613\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__25277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11002\,
            in2 => \_gnd_net_\,
            in3 => \N__10610\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__25277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10909\,
            in2 => \_gnd_net_\,
            in3 => \N__10607\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__25277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10711\,
            in2 => \_gnd_net_\,
            in3 => \N__10682\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__25277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10726\,
            in2 => \_gnd_net_\,
            in3 => \N__10679\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__25277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10696\,
            in2 => \_gnd_net_\,
            in3 => \N__10676\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10762\,
            in2 => \_gnd_net_\,
            in3 => \N__10673\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10747\,
            in2 => \_gnd_net_\,
            in3 => \N__10670\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10933\,
            in2 => \_gnd_net_\,
            in3 => \N__10667\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10823\,
            in2 => \_gnd_net_\,
            in3 => \N__10664\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10774\,
            in2 => \_gnd_net_\,
            in3 => \N__10661\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10787\,
            in2 => \_gnd_net_\,
            in3 => \N__10658\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10960\,
            in2 => \_gnd_net_\,
            in3 => \N__10841\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__25272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10735\,
            in2 => \_gnd_net_\,
            in3 => \N__10838\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__25268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10973\,
            in2 => \_gnd_net_\,
            in3 => \N__10835\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__25268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10811\,
            in3 => \N__10832\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__25268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10883\,
            in2 => \_gnd_net_\,
            in3 => \N__10829\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__25268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10798\,
            in2 => \_gnd_net_\,
            in3 => \N__10826\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10822\,
            in1 => \N__10807\,
            in2 => \N__10799\,
            in3 => \N__10786\,
            lcout => \reset_module_System.reset6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNISRMR1_10_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10775\,
            in1 => \N__10763\,
            in2 => \N__10751\,
            in3 => \N__10736\,
            lcout => \reset_module_System.reset6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10727\,
            in1 => \N__10712\,
            in2 => \N__10697\,
            in3 => \N__11003\,
            lcout => \reset_module_System.reset6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__11544\,
            in1 => \N__11522\,
            in2 => \N__11507\,
            in3 => \N__11482\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIR9N6_1_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10988\,
            in2 => \_gnd_net_\,
            in3 => \N__11457\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIA72I1_16_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10972\,
            in1 => \N__10961\,
            in2 => \N__10946\,
            in3 => \N__10943\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIMJ304_12_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10937\,
            in1 => \N__11543\,
            in2 => \N__10922\,
            in3 => \N__10919\,
            lcout => \reset_module_System.reset6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10913\,
            in1 => \N__10898\,
            in2 => \N__10859\,
            in3 => \N__10882\,
            lcout => \reset_module_System.reset6_15\,
            ltout => \reset_module_System.reset6_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11483\,
            in1 => \N__11506\,
            in2 => \N__10871\,
            in3 => \N__10868\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_1_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__12056\,
            in1 => \N__11564\,
            in2 => \N__12491\,
            in3 => \N__24919\,
            lcout => \uart_drone.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_rdy_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12039\,
            in2 => \_gnd_net_\,
            in3 => \N__11441\,
            lcout => uart_data_rdy_debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25287\,
            ce => 'H',
            sr => \N__24751\
        );

    \frame_dron_decoder_1.source_data_valid_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__11206\,
            in1 => \N__11240\,
            in2 => \_gnd_net_\,
            in3 => \N__11121\,
            lcout => drone_frame_decoder_data_rdy_debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25287\,
            ce => 'H',
            sr => \N__24751\
        );

    \frame_dron_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11357\,
            in2 => \_gnd_net_\,
            in3 => \N__11093\,
            lcout => OPEN,
            ltout => \frame_dron_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.state_ns_i_a2_2_0_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11009\,
            in1 => \N__11195\,
            in2 => \N__11186\,
            in3 => \N__11015\,
            lcout => \frame_dron_decoder_1.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \frame_dron_decoder_1.source_data_valid_2_sqmuxa_i_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24897\,
            lcout => \frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_0_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__11656\,
            in1 => \N__15267\,
            in2 => \_gnd_net_\,
            in3 => \N__24896\,
            lcout => \uart_pc.state_srsts_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_esr_1_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11296\,
            lcout => uart_drone_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25278\,
            ce => \N__11347\,
            sr => \N__11326\
        );

    \uart_drone.data_esr_3_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11281\,
            lcout => uart_drone_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25278\,
            ce => \N__11347\,
            sr => \N__11326\
        );

    \uart_drone.data_esr_0_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11311\,
            lcout => uart_drone_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25278\,
            ce => \N__11347\,
            sr => \N__11326\
        );

    \uart_drone.data_esr_5_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11830\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_drone_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25278\,
            ce => \N__11347\,
            sr => \N__11326\
        );

    \uart_drone.data_esr_6_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11608\,
            lcout => uart_drone_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25278\,
            ce => \N__11347\,
            sr => \N__11326\
        );

    \uart_drone.data_esr_7_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11644\,
            lcout => uart_drone_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25278\,
            ce => \N__11347\,
            sr => \N__11326\
        );

    \uart_drone.data_Aux_0_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__12040\,
            in1 => \N__11246\,
            in2 => \N__11312\,
            in3 => \N__11855\,
            lcout => \uart_drone.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25273\,
            ce => 'H',
            sr => \N__11801\
        );

    \uart_drone.data_Aux_1_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__11856\,
            in1 => \N__11420\,
            in2 => \N__11297\,
            in3 => \N__12041\,
            lcout => \uart_drone.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25273\,
            ce => 'H',
            sr => \N__11801\
        );

    \uart_drone.data_Aux_3_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__11857\,
            in1 => \N__11414\,
            in2 => \N__11282\,
            in3 => \N__12042\,
            lcout => \uart_drone.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25273\,
            ce => 'H',
            sr => \N__11801\
        );

    \uart_drone.data_Aux_RNO_0_4_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12314\,
            in1 => \N__12371\,
            in2 => \_gnd_net_\,
            in3 => \N__12447\,
            lcout => OPEN,
            ltout => \uart_drone.data_Auxce_0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_4_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__12043\,
            in1 => \N__11257\,
            in2 => \N__11267\,
            in3 => \N__11858\,
            lcout => \uart_drone.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25273\,
            ce => 'H',
            sr => \N__11801\
        );

    \uart_drone.data_Aux_RNO_0_5_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12313\,
            in1 => \N__12370\,
            in2 => \_gnd_net_\,
            in3 => \N__12446\,
            lcout => \uart_drone.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_0_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12310\,
            in1 => \N__12365\,
            in2 => \_gnd_net_\,
            in3 => \N__12443\,
            lcout => \uart_drone.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIDGR31_2_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__12169\,
            in1 => \N__12527\,
            in2 => \N__11939\,
            in3 => \N__11580\,
            lcout => \uart_drone.state_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_1_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__12311\,
            in1 => \N__12366\,
            in2 => \_gnd_net_\,
            in3 => \N__12444\,
            lcout => \uart_drone.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_3_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__12445\,
            in1 => \_gnd_net_\,
            in2 => \N__12374\,
            in3 => \N__12312\,
            lcout => \uart_drone.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI9E9J_2_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12170\,
            lcout => \uart_drone.N_126_li\,
            ltout => \uart_drone.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI9ADK1_4_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__11405\,
            in1 => \N__12528\,
            in2 => \N__11408\,
            in3 => \N__12135\,
            lcout => \uart_drone.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI5A9J_1_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__11759\,
            in1 => \N__11710\,
            in2 => \N__11762\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \uart_drone.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_2_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11582\,
            in2 => \_gnd_net_\,
            in3 => \N__11399\,
            lcout => \uart_drone.timer_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_1\,
            carryout => \uart_drone.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_3_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12174\,
            in2 => \_gnd_net_\,
            in3 => \N__11396\,
            lcout => \uart_drone.timer_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_2\,
            carryout => \uart_drone.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_4_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11938\,
            in2 => \_gnd_net_\,
            in3 => \N__11393\,
            lcout => \uart_drone.timer_Count_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_3_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__11735\,
            in1 => \N__24120\,
            in2 => \N__12245\,
            in3 => \N__11594\,
            lcout => \uart_drone.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_2_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__11588\,
            in1 => \N__12241\,
            in2 => \N__24169\,
            in3 => \N__11734\,
            lcout => \uart_drone.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_2_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110100"
        )
    port map (
            in0 => \N__12051\,
            in1 => \N__11562\,
            in2 => \N__12209\,
            in3 => \N__24899\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_2_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__11941\,
            in1 => \N__12176\,
            in2 => \N__11567\,
            in3 => \N__11563\,
            lcout => \uart_drone.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__11520\,
            in1 => \N__11501\,
            in2 => \_gnd_net_\,
            in3 => \N__11480\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11545\,
            in2 => \_gnd_net_\,
            in3 => \N__11461\,
            lcout => OPEN,
            ltout => \reset_module_System.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__11521\,
            in1 => \N__11502\,
            in2 => \N__11486\,
            in3 => \N__11481\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI40411_2_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__12129\,
            in1 => \N__11940\,
            in2 => \N__12208\,
            in3 => \N__12175\,
            lcout => \uart_drone.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_1_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__12442\,
            in1 => \N__12363\,
            in2 => \N__12473\,
            in3 => \N__12385\,
            lcout => \uart_drone.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25250\,
            ce => 'H',
            sr => \N__24781\
        );

    \uart_drone.bit_Count_0_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001100100"
        )
    port map (
            in0 => \N__12469\,
            in1 => \N__12441\,
            in2 => \N__12137\,
            in3 => \N__12082\,
            lcout => \uart_drone.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25250\,
            ce => 'H',
            sr => \N__24781\
        );

    \uart_drone_sync.Q_0__0_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11699\,
            lcout => uart_input_debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_3__0__0_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12263\,
            lcout => \uart_drone_sync.aux_3__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_1_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__11660\,
            in1 => \N__15247\,
            in2 => \N__11693\,
            in3 => \N__24918\,
            lcout => \uart_pc.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_2_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__12980\,
            in1 => \N__15246\,
            in2 => \N__11692\,
            in3 => \N__24898\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_2_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__11688\,
            in1 => \N__13183\,
            in2 => \N__11669\,
            in3 => \N__13040\,
            lcout => \uart_pc.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_0_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110101010101"
        )
    port map (
            in0 => \N__11666\,
            in1 => \N__13184\,
            in2 => \N__12836\,
            in3 => \N__12816\,
            lcout => \uart_pc.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_7_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__12015\,
            in1 => \N__11867\,
            in2 => \N__11645\,
            in3 => \N__12083\,
            lcout => \uart_drone.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25274\,
            ce => 'H',
            sr => \N__11800\
        );

    \uart_drone.data_Aux_2_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__11810\,
            in1 => \N__12014\,
            in2 => \N__11626\,
            in3 => \N__11866\,
            lcout => \uart_drone.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25274\,
            ce => 'H',
            sr => \N__11800\
        );

    \uart_drone.data_Aux_6_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__11816\,
            in1 => \N__12017\,
            in2 => \N__11609\,
            in3 => \N__11860\,
            lcout => \uart_drone.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25269\,
            ce => 'H',
            sr => \N__11793\
        );

    \uart_drone.data_Aux_5_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__11873\,
            in1 => \N__12016\,
            in2 => \N__11831\,
            in3 => \N__11859\,
            lcout => \uart_drone.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25269\,
            ce => 'H',
            sr => \N__11793\
        );

    \uart_drone.data_Aux_RNO_0_6_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12296\,
            in1 => \N__12373\,
            in2 => \_gnd_net_\,
            in3 => \N__12449\,
            lcout => \uart_drone.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_2_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__12295\,
            in1 => \N__12372\,
            in2 => \_gnd_net_\,
            in3 => \N__12448\,
            lcout => \uart_drone.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIOU0N_4_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__12136\,
            in1 => \N__12529\,
            in2 => \_gnd_net_\,
            in3 => \N__24903\,
            lcout => \uart_drone.state_RNIOU0NZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_0_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__24118\,
            in1 => \N__11761\,
            in2 => \N__11741\,
            in3 => \N__12238\,
            lcout => \uart_drone.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIAT1D1_4_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__11937\,
            in1 => \N__12523\,
            in2 => \N__24199\,
            in3 => \N__11887\,
            lcout => \uart_drone.N_143\,
            ltout => \uart_drone.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_4_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__11771\,
            in1 => \N__24168\,
            in2 => \N__11765\,
            in3 => \N__11740\,
            lcout => \uart_drone.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_1_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11760\,
            in2 => \_gnd_net_\,
            in3 => \N__11711\,
            lcout => OPEN,
            ltout => \uart_drone.timer_Count_RNO_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_1_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__12239\,
            in1 => \N__11739\,
            in2 => \N__11714\,
            in3 => \N__24119\,
            lcout => \uart_drone.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_4_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__24116\,
            in1 => \N__12218\,
            in2 => \N__12134\,
            in3 => \N__12240\,
            lcout => \uart_drone.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIU8TV1_3_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11927\,
            in1 => \N__12078\,
            in2 => \_gnd_net_\,
            in3 => \N__12173\,
            lcout => \uart_drone.N_144_1\,
            ltout => \uart_drone.N_144_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_3_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__12200\,
            in1 => \N__12182\,
            in2 => \N__12212\,
            in3 => \N__24117\,
            lcout => \uart_drone.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_3_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__12172\,
            in1 => \N__12118\,
            in2 => \N__12207\,
            in3 => \N__11928\,
            lcout => \uart_drone.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI62411_4_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__11926\,
            in1 => \N__12171\,
            in2 => \N__12133\,
            in3 => \N__12522\,
            lcout => \uart_drone.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI63LK2_3_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__12122\,
            in1 => \N__12468\,
            in2 => \_gnd_net_\,
            in3 => \N__12077\,
            lcout => \uart_drone.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNIJOJC1_2_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12281\,
            in1 => \N__12345\,
            in2 => \_gnd_net_\,
            in3 => \N__12422\,
            lcout => \uart_drone.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_0_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__12484\,
            in1 => \N__12013\,
            in2 => \_gnd_net_\,
            in3 => \N__24900\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_0_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__11942\,
            in1 => \N__11891\,
            in2 => \N__11876\,
            in3 => \N__12530\,
            lcout => \uart_drone.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNO_0_2_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12467\,
            in2 => \_gnd_net_\,
            in3 => \N__12423\,
            lcout => \uart_drone.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_2_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__12392\,
            in1 => \N__12386\,
            in2 => \N__12309\,
            in3 => \N__12364\,
            lcout => \uart_drone.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25238\,
            ce => 'H',
            sr => \N__24782\
        );

    \uart_drone_sync.aux_2__0__0_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13379\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone_sync.aux_2__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_6_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__12257\,
            in1 => \N__15266\,
            in2 => \N__14623\,
            in3 => \N__12869\,
            lcout => \uart_pc.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25297\,
            ce => 'H',
            sr => \N__12575\
        );

    \uart_pc.data_Aux_RNO_0_6_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12702\,
            in1 => \N__12769\,
            in2 => \_gnd_net_\,
            in3 => \N__12623\,
            lcout => \uart_pc.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_1_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__12701\,
            in1 => \N__12768\,
            in2 => \_gnd_net_\,
            in3 => \N__12622\,
            lcout => \uart_pc.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__12776\,
            in1 => \N__15251\,
            in2 => \N__13348\,
            in3 => \N__12862\,
            lcout => \uart_pc.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25292\,
            ce => 'H',
            sr => \N__12574\
        );

    \uart_pc.data_Aux_1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__12863\,
            in1 => \N__13363\,
            in2 => \N__15269\,
            in3 => \N__12251\,
            lcout => \uart_pc.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25292\,
            ce => 'H',
            sr => \N__12574\
        );

    \uart_pc.data_Aux_2_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__12557\,
            in1 => \N__15252\,
            in2 => \N__13309\,
            in3 => \N__12864\,
            lcout => \uart_pc.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25292\,
            ce => 'H',
            sr => \N__12574\
        );

    \uart_pc.data_Aux_3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__12865\,
            in1 => \N__13288\,
            in2 => \N__15270\,
            in3 => \N__12551\,
            lcout => \uart_pc.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25292\,
            ce => 'H',
            sr => \N__12574\
        );

    \uart_pc.data_Aux_4_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__12539\,
            in1 => \N__15253\,
            in2 => \N__13331\,
            in3 => \N__12866\,
            lcout => \uart_pc.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25292\,
            ce => 'H',
            sr => \N__12574\
        );

    \uart_pc.data_Aux_5_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__12867\,
            in1 => \N__13273\,
            in2 => \N__15271\,
            in3 => \N__12545\,
            lcout => \uart_pc.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25292\,
            ce => 'H',
            sr => \N__12574\
        );

    \uart_pc.data_Aux_7_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__12868\,
            in1 => \N__13261\,
            in2 => \N__15272\,
            in3 => \N__12959\,
            lcout => \uart_pc.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25292\,
            ce => 'H',
            sr => \N__12574\
        );

    \uart_pc.state_RNIEAGS_4_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__12919\,
            in1 => \N__12818\,
            in2 => \_gnd_net_\,
            in3 => \N__24901\,
            lcout => \uart_pc.state_RNIEAGSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_2_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__12756\,
            in1 => \N__12692\,
            in2 => \_gnd_net_\,
            in3 => \N__12618\,
            lcout => \uart_pc.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_3_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__12619\,
            in1 => \_gnd_net_\,
            in2 => \N__12703\,
            in3 => \N__12757\,
            lcout => \uart_pc.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12759\,
            in1 => \N__12699\,
            in2 => \_gnd_net_\,
            in3 => \N__12621\,
            lcout => \uart_pc.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_4_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__12620\,
            in1 => \_gnd_net_\,
            in2 => \N__12704\,
            in3 => \N__12758\,
            lcout => \uart_pc.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12755\,
            in1 => \N__12691\,
            in2 => \_gnd_net_\,
            in3 => \N__12617\,
            lcout => \uart_pc.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_2_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__12722\,
            in1 => \N__12700\,
            in2 => \N__12770\,
            in3 => \N__12716\,
            lcout => \uart_pc.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25283\,
            ce => 'H',
            sr => \N__24741\
        );

    \uart_pc.bit_Count_RNI4U6E1_2_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12754\,
            in1 => \N__12670\,
            in2 => \_gnd_net_\,
            in3 => \N__12597\,
            lcout => \uart_pc.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIITIF1_4_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__13174\,
            in1 => \N__13039\,
            in2 => \N__12920\,
            in3 => \N__12817\,
            lcout => \uart_pc.un1_state_4_0\,
            ltout => \uart_pc.un1_state_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIUPE73_3_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12916\,
            in2 => \N__12725\,
            in3 => \N__12950\,
            lcout => \uart_pc.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNO_0_2_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12634\,
            in2 => \_gnd_net_\,
            in3 => \N__12598\,
            lcout => \uart_pc.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_1_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__12690\,
            in1 => \N__12715\,
            in2 => \N__12647\,
            in3 => \N__12616\,
            lcout => \uart_pc.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25275\,
            ce => 'H',
            sr => \N__24746\
        );

    \uart_pc.bit_Count_0_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100100000"
        )
    port map (
            in0 => \N__12917\,
            in1 => \N__12957\,
            in2 => \N__12646\,
            in3 => \N__12615\,
            lcout => \uart_pc.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25275\,
            ce => 'H',
            sr => \N__24746\
        );

    \uart_pc.timer_Count_RNIPD2K1_2_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__13032\,
            in1 => \N__13118\,
            in2 => \N__13181\,
            in3 => \N__12807\,
            lcout => \uart_pc.state_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_3_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__12905\,
            in1 => \N__13173\,
            in2 => \N__12989\,
            in3 => \N__13035\,
            lcout => OPEN,
            ltout => \uart_pc.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_3_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__12987\,
            in1 => \N__12928\,
            in2 => \N__12992\,
            in3 => \N__24193\,
            lcout => \uart_pc.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIGRIF1_2_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__12904\,
            in1 => \N__13169\,
            in2 => \N__12988\,
            in3 => \N__13034\,
            lcout => \uart_pc.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_4_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__12929\,
            in1 => \N__24192\,
            in2 => \N__12918\,
            in3 => \N__13091\,
            lcout => \uart_pc.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNI5UFA2_3_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__13033\,
            in1 => \_gnd_net_\,
            in2 => \N__13182\,
            in3 => \N__12958\,
            lcout => \uart_pc.N_144_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_0_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__13225\,
            in1 => \N__13087\,
            in2 => \N__24212\,
            in3 => \N__13053\,
            lcout => \uart_pc.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIBLRB2_4_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__12812\,
            in1 => \N__12829\,
            in2 => \N__13205\,
            in3 => \N__12909\,
            lcout => \uart_pc.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_1_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13224\,
            in2 => \_gnd_net_\,
            in3 => \N__13238\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIVT8S_2_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13030\,
            in2 => \_gnd_net_\,
            in3 => \N__13116\,
            lcout => \uart_pc.N_126_li\,
            ltout => \uart_pc.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIMQ8T1_4_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__13159\,
            in1 => \N__12811\,
            in2 => \N__12779\,
            in3 => \N__24194\,
            lcout => \uart_pc.N_143\,
            ltout => \uart_pc.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_1_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__13054\,
            in1 => \N__24195\,
            in2 => \N__13247\,
            in3 => \N__13244\,
            lcout => \uart_pc.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIRP8S_1_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__13223\,
            in1 => \N__13237\,
            in2 => \N__13226\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => \uart_pc.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_2_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13117\,
            in2 => \_gnd_net_\,
            in3 => \N__13196\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_1\,
            carryout => \uart_pc.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_3_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13031\,
            in2 => \_gnd_net_\,
            in3 => \N__13193\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_2\,
            carryout => \uart_pc.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_4_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13165\,
            in2 => \_gnd_net_\,
            in3 => \N__13190\,
            lcout => OPEN,
            ltout => \uart_pc.timer_Count_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_4_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__13064\,
            in1 => \N__13090\,
            in2 => \N__13187\,
            in3 => \N__24184\,
            lcout => \uart_pc.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_2_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__13124\,
            in1 => \N__13088\,
            in2 => \N__24210\,
            in3 => \N__13062\,
            lcout => \uart_pc.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_3_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__13097\,
            in1 => \N__13089\,
            in2 => \N__24211\,
            in3 => \N__13063\,
            lcout => \uart_pc.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_0__0__0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13391\,
            lcout => \uart_drone_sync.aux_0__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_1__0__0_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13385\,
            lcout => \uart_drone_sync.aux_1__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_esr_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13370\,
            lcout => uart_pc_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25289\,
            ce => \N__14601\,
            sr => \N__14808\
        );

    \uart_pc.data_esr_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13352\,
            lcout => uart_pc_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25289\,
            ce => \N__14601\,
            sr => \N__14808\
        );

    \uart_pc.data_esr_4_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13327\,
            lcout => uart_pc_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25284\,
            ce => \N__14606\,
            sr => \N__14810\
        );

    \uart_pc.data_esr_2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13310\,
            lcout => uart_pc_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25284\,
            ce => \N__14606\,
            sr => \N__14810\
        );

    \uart_pc.data_esr_3_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13292\,
            lcout => uart_pc_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25284\,
            ce => \N__14606\,
            sr => \N__14810\
        );

    \uart_pc.data_esr_5_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_pc_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25284\,
            ce => \N__14606\,
            sr => \N__14810\
        );

    \uart_pc.data_esr_7_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_pc_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25284\,
            ce => \N__14606\,
            sr => \N__14810\
        );

    \uart_frame_decoder.state_1_1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__13763\,
            in1 => \N__23932\,
            in2 => \N__13772\,
            in3 => \N__23904\,
            lcout => \uart_frame_decoder.state_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25280\,
            ce => 'H',
            sr => \N__24740\
        );

    \uart_frame_decoder.state_1_RNIC4PK_6_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13852\,
            in2 => \_gnd_net_\,
            in3 => \N__23823\,
            lcout => \uart_frame_decoder.source_offset1data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIE6PK_8_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13807\,
            lcout => \uart_frame_decoder.source_offset3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNID5PK_7_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23825\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13828\,
            lcout => \uart_frame_decoder.source_offset2data_1_sqmuxa\,
            ltout => \uart_frame_decoder.source_offset2data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIAIVT_7_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13415\,
            in3 => \N__24904\,
            lcout => \uart_frame_decoder.source_offset2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI9HVT_6_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13840\,
            in2 => \_gnd_net_\,
            in3 => \N__24905\,
            lcout => \uart_frame_decoder.source_offset1data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIBJVT_8_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13792\,
            in2 => \_gnd_net_\,
            in3 => \N__24906\,
            lcout => \uart_frame_decoder.source_offset3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13412\,
            in2 => \N__13961\,
            in3 => \N__13960\,
            lcout => \uart_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \uart_frame_decoder.un1_WDT_cry_0\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13406\,
            in2 => \_gnd_net_\,
            in3 => \N__13400\,
            lcout => \uart_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_0\,
            carryout => \uart_frame_decoder.un1_WDT_cry_1\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_2_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13397\,
            in2 => \_gnd_net_\,
            in3 => \N__13448\,
            lcout => \uart_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_1\,
            carryout => \uart_frame_decoder.un1_WDT_cry_2\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_3_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13445\,
            in2 => \_gnd_net_\,
            in3 => \N__13439\,
            lcout => \uart_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_2\,
            carryout => \uart_frame_decoder.un1_WDT_cry_3\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_4_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13907\,
            in2 => \_gnd_net_\,
            in3 => \N__13436\,
            lcout => \uart_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_3\,
            carryout => \uart_frame_decoder.un1_WDT_cry_4\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_5_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13934\,
            in2 => \_gnd_net_\,
            in3 => \N__13433\,
            lcout => \uart_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_4\,
            carryout => \uart_frame_decoder.un1_WDT_cry_5\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_6_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14111\,
            in2 => \_gnd_net_\,
            in3 => \N__13430\,
            lcout => \uart_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_5\,
            carryout => \uart_frame_decoder.un1_WDT_cry_6\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_7_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14042\,
            in2 => \_gnd_net_\,
            in3 => \N__13427\,
            lcout => \uart_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_6\,
            carryout => \uart_frame_decoder.un1_WDT_cry_7\,
            clk => \N__25265\,
            ce => 'H',
            sr => \N__13889\
        );

    \uart_frame_decoder.WDT_8_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13946\,
            in2 => \_gnd_net_\,
            in3 => \N__13424\,
            lcout => \uart_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \uart_frame_decoder.un1_WDT_cry_8\,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.WDT_9_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13921\,
            in2 => \_gnd_net_\,
            in3 => \N__13421\,
            lcout => \uart_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_8\,
            carryout => \uart_frame_decoder.un1_WDT_cry_9\,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.WDT_10_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14084\,
            in2 => \_gnd_net_\,
            in3 => \N__13418\,
            lcout => \uart_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_9\,
            carryout => \uart_frame_decoder.un1_WDT_cry_10\,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.WDT_11_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14099\,
            in2 => \_gnd_net_\,
            in3 => \N__13463\,
            lcout => \uart_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_10\,
            carryout => \uart_frame_decoder.un1_WDT_cry_11\,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.WDT_12_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14057\,
            in2 => \_gnd_net_\,
            in3 => \N__13460\,
            lcout => \uart_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_11\,
            carryout => \uart_frame_decoder.un1_WDT_cry_12\,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.WDT_13_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14071\,
            in2 => \_gnd_net_\,
            in3 => \N__13457\,
            lcout => \uart_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_12\,
            carryout => \uart_frame_decoder.un1_WDT_cry_13\,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.WDT_14_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14008\,
            in2 => \_gnd_net_\,
            in3 => \N__13454\,
            lcout => \uart_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_13\,
            carryout => \uart_frame_decoder.un1_WDT_cry_14\,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.WDT_15_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13981\,
            in2 => \_gnd_net_\,
            in3 => \N__13451\,
            lcout => \uart_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25258\,
            ce => 'H',
            sr => \N__13885\
        );

    \uart_frame_decoder.source_offset1data_esr_0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21103\,
            lcout => \frame_decoder_OFF1data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_offset1data_esr_1_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20974\,
            lcout => \frame_decoder_OFF1data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_offset1data_esr_2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20898\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF1data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_offset1data_esr_3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF1data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_offset1data_esr_4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20727\,
            lcout => \frame_decoder_OFF1data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_offset1data_esr_5_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF1data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_offset1data_esr_6_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20632\,
            lcout => \frame_decoder_OFF1data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_offset1data_esr_7_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20527\,
            lcout => \frame_decoder_OFF1data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25252\,
            ce => \N__13475\,
            sr => \N__24756\
        );

    \uart_frame_decoder.source_CH1data_esr_0_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21110\,
            lcout => \frame_decoder_CH1data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25245\,
            ce => \N__14312\,
            sr => \N__24759\
        );

    \uart_frame_decoder.source_CH1data_esr_1_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20975\,
            lcout => \frame_decoder_CH1data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25245\,
            ce => \N__14312\,
            sr => \N__24759\
        );

    \uart_frame_decoder.source_CH1data_esr_2_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20899\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH1data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25245\,
            ce => \N__14312\,
            sr => \N__24759\
        );

    \uart_frame_decoder.source_CH1data_esr_3_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20813\,
            lcout => \frame_decoder_CH1data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25245\,
            ce => \N__14312\,
            sr => \N__24759\
        );

    \uart_frame_decoder.source_CH1data_esr_4_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20716\,
            lcout => \frame_decoder_CH1data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25245\,
            ce => \N__14312\,
            sr => \N__24759\
        );

    \uart_frame_decoder.source_CH1data_esr_5_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH1data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25245\,
            ce => \N__14312\,
            sr => \N__24759\
        );

    \uart_frame_decoder.source_CH1data_esr_6_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20633\,
            lcout => \frame_decoder_CH1data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25245\,
            ce => \N__14312\,
            sr => \N__24759\
        );

    \uart_frame_decoder.source_CH1data_esr_7_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20536\,
            lcout => \frame_decoder_CH1data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25239\,
            ce => \N__14308\,
            sr => \N__24765\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26102\,
            in1 => \N__14327\,
            in2 => \_gnd_net_\,
            in3 => \N__15421\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_4_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14981\,
            lcout => \ppm_encoder_1.rudderZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25228\,
            ce => \N__21739\,
            sr => \N__24774\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23594\,
            in1 => \_gnd_net_\,
            in2 => \N__22771\,
            in3 => \N__22330\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19418\,
            in1 => \N__22705\,
            in2 => \_gnd_net_\,
            in3 => \N__23592\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23593\,
            in1 => \_gnd_net_\,
            in2 => \N__22770\,
            in3 => \N__19417\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__23086\,
            in1 => \N__22704\,
            in2 => \_gnd_net_\,
            in3 => \N__23591\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000001010"
        )
    port map (
            in0 => \N__22188\,
            in1 => \N__26071\,
            in2 => \N__23192\,
            in3 => \N__25800\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__24920\,
            in1 => \N__22189\,
            in2 => \N__13478\,
            in3 => \N__23589\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__23160\,
            in1 => \N__26072\,
            in2 => \N__25807\,
            in3 => \N__22693\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIE3D21_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15626\,
            in1 => \N__22239\,
            in2 => \N__22195\,
            in3 => \N__23156\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_162_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14510\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIGD613_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14512\,
            in1 => \N__15997\,
            in2 => \_gnd_net_\,
            in3 => \N__23510\,
            lcout => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15404\,
            in2 => \N__22695\,
            in3 => \N__25931\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13484\,
            in3 => \N__23506\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22190\,
            in3 => \N__14351\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13481\,
            in3 => \N__23505\,
            lcout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14509\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23509\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIR7352_3_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001000101101"
        )
    port map (
            in0 => \N__18637\,
            in1 => \N__19988\,
            in2 => \N__22511\,
            in3 => \N__16124\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI60223_3_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13499\,
            in3 => \N__15763\,
            lcout => \ppm_encoder_1.init_pulses_RNI60223Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__22649\,
            in1 => \N__22503\,
            in2 => \_gnd_net_\,
            in3 => \N__23511\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__23512\,
            in1 => \_gnd_net_\,
            in2 => \N__22510\,
            in3 => \N__22650\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_1_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19989\,
            in2 => \_gnd_net_\,
            in3 => \N__25542\,
            lcout => \ppm_encoder_1.throttleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25214\,
            ce => 'H',
            sr => \N__24787\
        );

    \ppm_encoder_1.throttle_2_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13496\,
            lcout => \ppm_encoder_1.throttleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25214\,
            ce => 'H',
            sr => \N__24787\
        );

    \ppm_encoder_1.throttle_RNIR7352_2_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__13494\,
            in1 => \N__22136\,
            in2 => \N__18665\,
            in3 => \N__16123\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__26063\,
            in1 => \N__25808\,
            in2 => \_gnd_net_\,
            in3 => \N__13495\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22345\,
            in1 => \N__23655\,
            in2 => \N__14525\,
            in3 => \N__16139\,
            lcout => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_6_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19515\,
            in1 => \N__19700\,
            in2 => \N__13625\,
            in3 => \N__15674\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25208\,
            ce => 'H',
            sr => \N__24793\
        );

    \ppm_encoder_1.init_pulses_RNIERUS_6_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22344\,
            in1 => \N__22779\,
            in2 => \_gnd_net_\,
            in3 => \N__23653\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__23656\,
            in1 => \N__22414\,
            in2 => \N__16147\,
            in3 => \N__14524\,
            lcout => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_13_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19699\,
            in1 => \N__13565\,
            in2 => \N__19549\,
            in3 => \N__15872\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25208\,
            ce => 'H',
            sr => \N__24793\
        );

    \ppm_encoder_1.init_pulses_RNISFRP_13_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23654\,
            in1 => \_gnd_net_\,
            in2 => \N__22822\,
            in3 => \N__22413\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13553\,
            in2 => \N__14537\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_1_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13544\,
            in2 => \_gnd_net_\,
            in3 => \N__13535\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_2_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14483\,
            in2 => \N__13532\,
            in3 => \N__13520\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_3_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13517\,
            in2 => \_gnd_net_\,
            in3 => \N__13508\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_4_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14633\,
            in2 => \_gnd_net_\,
            in3 => \N__13505\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_5_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19721\,
            in2 => \_gnd_net_\,
            in3 => \N__13502\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_6_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13643\,
            in2 => \N__13634\,
            in3 => \N__13616\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_7_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13613\,
            in2 => \_gnd_net_\,
            in3 => \N__13604\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_8_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17402\,
            in2 => \_gnd_net_\,
            in3 => \N__13601\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_8\,
            ltout => OPEN,
            carryin => \bfn_7_27_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_9_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17354\,
            in2 => \_gnd_net_\,
            in3 => \N__13598\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_10_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14408\,
            in2 => \_gnd_net_\,
            in3 => \N__13595\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_11_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14447\,
            in2 => \_gnd_net_\,
            in3 => \N__13592\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_12_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14576\,
            in2 => \_gnd_net_\,
            in3 => \N__13589\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_13_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13586\,
            in2 => \N__13577\,
            in3 => \N__13556\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13691\,
            in2 => \_gnd_net_\,
            in3 => \N__13679\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_15_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14552\,
            in2 => \_gnd_net_\,
            in3 => \N__13676\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_16_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13658\,
            in2 => \_gnd_net_\,
            in3 => \N__13673\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_16\,
            ltout => OPEN,
            carryin => \bfn_7_28_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_17_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13664\,
            in2 => \_gnd_net_\,
            in3 => \N__13670\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_18_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__23707\,
            in1 => \N__15985\,
            in2 => \N__22840\,
            in3 => \N__13667\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23706\,
            in1 => \_gnd_net_\,
            in2 => \N__22839\,
            in3 => \N__16072\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__15956\,
            in1 => \N__22827\,
            in2 => \_gnd_net_\,
            in3 => \N__23705\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_0__0__0_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_2__0__0_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13721\,
            lcout => \uart_pc_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_1__0__0_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13727\,
            lcout => \uart_pc_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_3__0__0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13715\,
            lcout => \uart_pc_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.Q_0__0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13709\,
            lcout => uart_input_pc_sync,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNILR1B2_2_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__15221\,
            in1 => \N__15166\,
            in2 => \_gnd_net_\,
            in3 => \N__24173\,
            lcout => \uart_pc.timer_Count_RNILR1B2Z0Z_2\,
            ltout => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIE94V3_2_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__15167\,
            in1 => \_gnd_net_\,
            in2 => \N__13700\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.state_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13762\,
            in1 => \N__15317\,
            in2 => \_gnd_net_\,
            in3 => \N__14770\,
            lcout => \uart_frame_decoder.N_39_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_3_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13761\,
            in1 => \N__15316\,
            in2 => \_gnd_net_\,
            in3 => \N__13781\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_RNO_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_1_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__13739\,
            in1 => \N__23953\,
            in2 => \N__13697\,
            in3 => \N__23931\,
            lcout => \uart_frame_decoder.state_1_ns_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26310\,
            in2 => \_gnd_net_\,
            in3 => \N__21065\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIDPNH_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20483\,
            in1 => \N__13760\,
            in2 => \N__13694\,
            in3 => \N__20851\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26309\,
            in1 => \N__20850\,
            in2 => \N__20505\,
            in3 => \N__21069\,
            lcout => \uart_frame_decoder.N_138_4\,
            ltout => \uart_frame_decoder.N_138_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14769\,
            in2 => \N__13775\,
            in3 => \_gnd_net_\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_2_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__15309\,
            in1 => \N__13759\,
            in2 => \N__14771\,
            in3 => \N__23826\,
            lcout => \uart_frame_decoder.state_1_RNO_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__20599\,
            in1 => \N__20955\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23827\,
            in1 => \N__20673\,
            in2 => \N__13733\,
            in3 => \N__20766\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNI5CUL2_15_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__14012\,
            in1 => \N__13985\,
            in2 => \N__23831\,
            in3 => \N__14021\,
            lcout => \uart_frame_decoder.N_85\,
            ltout => \uart_frame_decoder.N_85_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_3_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14893\,
            in2 => \N__13730\,
            in3 => \N__21362\,
            lcout => \uart_frame_decoder.state_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25271\,
            ce => 'H',
            sr => \N__24743\
        );

    \uart_frame_decoder.state_1_4_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__14879\,
            in1 => \N__23845\,
            in2 => \_gnd_net_\,
            in3 => \N__23898\,
            lcout => \uart_frame_decoder.state_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25271\,
            ce => 'H',
            sr => \N__24743\
        );

    \uart_frame_decoder.state_1_5_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__23899\,
            in1 => \N__17794\,
            in2 => \_gnd_net_\,
            in3 => \N__26381\,
            lcout => \uart_frame_decoder.state_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25271\,
            ce => 'H',
            sr => \N__24743\
        );

    \uart_frame_decoder.state_1_6_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__13853\,
            in1 => \N__17780\,
            in2 => \_gnd_net_\,
            in3 => \N__23900\,
            lcout => \uart_frame_decoder.state_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25271\,
            ce => 'H',
            sr => \N__24743\
        );

    \uart_frame_decoder.state_1_7_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__23901\,
            in1 => \N__13841\,
            in2 => \_gnd_net_\,
            in3 => \N__13829\,
            lcout => \uart_frame_decoder.state_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25271\,
            ce => 'H',
            sr => \N__24743\
        );

    \uart_frame_decoder.state_1_8_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__13817\,
            in1 => \N__13808\,
            in2 => \_gnd_net_\,
            in3 => \N__23902\,
            lcout => \uart_frame_decoder.state_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25271\,
            ce => 'H',
            sr => \N__24743\
        );

    \uart_frame_decoder.state_1_9_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__23903\,
            in1 => \_gnd_net_\,
            in2 => \N__13796\,
            in3 => \N__14753\,
            lcout => \uart_frame_decoder.state_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25271\,
            ce => 'H',
            sr => \N__24743\
        );

    \uart_frame_decoder.source_offset2data_esr_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21101\,
            lcout => \frame_decoder_OFF2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset2data_esr_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20988\,
            lcout => \frame_decoder_OFF2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset2data_esr_2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20882\,
            lcout => \frame_decoder_OFF2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset2data_esr_7_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20507\,
            lcout => \frame_decoder_OFF2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset2data_esr_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20725\,
            lcout => \frame_decoder_OFF2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset2data_esr_5_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26342\,
            lcout => \frame_decoder_OFF2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset2data_esr_6_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20619\,
            lcout => \frame_decoder_OFF2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset2data_esr_3_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25266\,
            ce => \N__13868\,
            sr => \N__24747\
        );

    \uart_frame_decoder.source_offset3data_esr_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21102\,
            lcout => \frame_decoder_OFF3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.source_offset3data_esr_1_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20989\,
            lcout => \frame_decoder_OFF3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.source_offset3data_esr_2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20897\,
            lcout => \frame_decoder_OFF3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.source_offset3data_esr_3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20811\,
            lcout => \frame_decoder_OFF3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.source_offset3data_esr_4_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20726\,
            lcout => \frame_decoder_OFF3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.source_offset3data_esr_5_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26359\,
            lcout => \frame_decoder_OFF3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.source_offset3data_esr_6_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.source_offset3data_esr_7_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20526\,
            lcout => \frame_decoder_OFF3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25259\,
            ce => \N__14117\,
            sr => \N__24752\
        );

    \uart_frame_decoder.WDT_RNIBI7E_6_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14055\,
            in1 => \N__14097\,
            in2 => \_gnd_net_\,
            in3 => \N__14110\,
            lcout => \uart_frame_decoder.WDT8lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIAGPB_10_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__14098\,
            in1 => \N__14083\,
            in2 => \N__14072\,
            in3 => \N__14056\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIM8N32_7_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__14041\,
            in1 => \N__13895\,
            in2 => \N__14030\,
            in3 => \N__14027\,
            lcout => \uart_frame_decoder.WDT8lt14_0\,
            ltout => \uart_frame_decoder.WDT8lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNI17K92_15_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14004\,
            in2 => \N__13988\,
            in3 => \N__13977\,
            lcout => \uart_frame_decoder.WDT8_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIQAB11_4_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13945\,
            in1 => \N__13933\,
            in2 => \N__13922\,
            in3 => \N__13906\,
            lcout => \uart_frame_decoder.WDT_RNIQAB11Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_RNIHJ501_0_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__16618\,
            in1 => \N__23816\,
            in2 => \_gnd_net_\,
            in3 => \N__15327\,
            lcout => \uart_frame_decoder.count_RNIHJ501Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__23817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24902\,
            lcout => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16536\,
            in2 => \N__16583\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \scaler_1.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14231\,
            in2 => \N__14225\,
            in3 => \N__14216\,
            lcout => \scaler_1.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_0\,
            carryout => \scaler_1.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14213\,
            in2 => \N__14207\,
            in3 => \N__14198\,
            lcout => \scaler_1.un3_source_data_0_cry_1_c_RNIISC11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_1\,
            carryout => \scaler_1.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14195\,
            in2 => \N__14189\,
            in3 => \N__14180\,
            lcout => \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_2\,
            carryout => \scaler_1.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14177\,
            in2 => \N__14171\,
            in3 => \N__14162\,
            lcout => \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_3\,
            carryout => \scaler_1.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14159\,
            in2 => \N__14153\,
            in3 => \N__14144\,
            lcout => \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_4\,
            carryout => \scaler_1.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14141\,
            in2 => \N__14135\,
            in3 => \N__14126\,
            lcout => \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_5\,
            carryout => \scaler_1.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14288\,
            in2 => \_gnd_net_\,
            in3 => \N__14123\,
            lcout => \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_6\,
            carryout => \scaler_1.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14261\,
            in2 => \N__21850\,
            in3 => \N__14120\,
            lcout => \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \scaler_1.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14291\,
            lcout => \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_1_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__14254\,
            in1 => \N__14697\,
            in2 => \_gnd_net_\,
            in3 => \N__16635\,
            lcout => \uart_frame_decoder.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14269\,
            in2 => \_gnd_net_\,
            in3 => \N__14281\,
            lcout => \scaler_1.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.N_508_i_l_ofx_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__14282\,
            in1 => \_gnd_net_\,
            in2 => \N__14273\,
            in3 => \_gnd_net_\,
            lcout => \scaler_1.N_508_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_2_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__16636\,
            in1 => \N__14255\,
            in2 => \N__14704\,
            in3 => \N__14725\,
            lcout => \uart_frame_decoder.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_0_c_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16694\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \uart_frame_decoder.count8_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_1_c_inv_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14243\,
            in2 => \_gnd_net_\,
            in3 => \N__14693\,
            lcout => \uart_frame_decoder.count8_axb_1\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.count8_cry_0\,
            carryout => \uart_frame_decoder.count8_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_2_c_inv_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14237\,
            in2 => \N__21848\,
            in3 => \N__14721\,
            lcout => \uart_frame_decoder.count_i_2\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.count8_cry_1\,
            carryout => \uart_frame_decoder.count8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_THRU_LUT4_0_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14315\,
            lcout => \uart_frame_decoder.count8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_4_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15020\,
            lcout => \ppm_encoder_1.aileronZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25229\,
            ce => \N__21707\,
            sr => \N__24775\
        );

    \ppm_encoder_1.elevator_esr_4_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14999\,
            lcout => \ppm_encoder_1.elevatorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25229\,
            ce => \N__21707\,
            sr => \N__24775\
        );

    \ppm_encoder_1.rudder_esr_5_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16226\,
            lcout => \ppm_encoder_1.rudderZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25229\,
            ce => \N__21707\,
            sr => \N__24775\
        );

    \ppm_encoder_1.throttle_esr_4_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15104\,
            lcout => \ppm_encoder_1.throttleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25229\,
            ce => \N__21707\,
            sr => \N__24775\
        );

    \ppm_encoder_1.elevator_esr_5_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15116\,
            lcout => \ppm_encoder_1.elevatorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25229\,
            ce => \N__21707\,
            sr => \N__24775\
        );

    \ppm_encoder_1.throttle_esr_5_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15128\,
            lcout => \ppm_encoder_1.throttleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25229\,
            ce => \N__21707\,
            sr => \N__24775\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__23628\,
            in1 => \N__23166\,
            in2 => \N__14396\,
            in3 => \N__24215\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25225\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111111010"
        )
    port map (
            in0 => \N__22240\,
            in1 => \N__22751\,
            in2 => \N__24930\,
            in3 => \N__23630\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25225\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI5DVT_2_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21361\,
            in2 => \_gnd_net_\,
            in3 => \N__24912\,
            lcout => \uart_frame_decoder.source_CH1data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__23629\,
            in1 => \N__24916\,
            in2 => \N__26090\,
            in3 => \N__15476\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25225\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22024\,
            in1 => \N__22750\,
            in2 => \_gnd_net_\,
            in3 => \N__23627\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14369\,
            in3 => \N__14348\,
            lcout => \ppm_encoder_1.N_230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111111010"
        )
    port map (
            in0 => \N__15457\,
            in1 => \N__22694\,
            in2 => \N__24931\,
            in3 => \N__23556\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23554\,
            in1 => \N__24214\,
            in2 => \N__14395\,
            in3 => \N__14350\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__14368\,
            in1 => \N__14378\,
            in2 => \N__24932\,
            in3 => \N__23555\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__14367\,
            in1 => \N__14349\,
            in2 => \N__15458\,
            in3 => \N__15474\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__18517\,
            in1 => \N__23553\,
            in2 => \N__14333\,
            in3 => \N__18440\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIALN65_1_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001111"
        )
    port map (
            in0 => \N__19995\,
            in1 => \N__15518\,
            in2 => \N__14330\,
            in3 => \N__18644\,
            lcout => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15437\,
            in1 => \N__15392\,
            in2 => \_gnd_net_\,
            in3 => \N__15624\,
            lcout => \ppm_encoder_1.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22242\,
            in1 => \N__25932\,
            in2 => \N__15625\,
            in3 => \N__23995\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_1_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19473\,
            in1 => \N__19701\,
            in2 => \N__14426\,
            in3 => \N__15491\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25215\,
            ce => 'H',
            sr => \N__24788\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__22687\,
            in1 => \N__23079\,
            in2 => \_gnd_net_\,
            in3 => \N__23572\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21468\,
            in3 => \N__23994\,
            lcout => \ppm_encoder_1.PPM_STATE_62_d\,
            ltout => \ppm_encoder_1.PPM_STATE_62_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22241\,
            in1 => \N__25930\,
            in2 => \N__14414\,
            in3 => \N__15617\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_0_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__24257\,
            in1 => \N__21467\,
            in2 => \N__24027\,
            in3 => \N__24280\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25215\,
            ce => 'H',
            sr => \N__24788\
        );

    \ppm_encoder_1.PPM_STATE_1_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24284\,
            in3 => \N__24019\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25215\,
            ce => 'H',
            sr => \N__24788\
        );

    \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__20026\,
            in1 => \N__16127\,
            in2 => \N__23676\,
            in3 => \N__14513\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_0_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000000110010"
        )
    port map (
            in0 => \N__19497\,
            in1 => \N__19694\,
            in2 => \N__14411\,
            in3 => \N__15530\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25209\,
            ce => 'H',
            sr => \N__24794\
        );

    \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20025\,
            in1 => \N__14514\,
            in2 => \N__23677\,
            in3 => \N__16125\,
            lcout => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23683\,
            in1 => \_gnd_net_\,
            in2 => \N__22752\,
            in3 => \N__20024\,
            lcout => \ppm_encoder_1.un1_init_pulses_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22138\,
            in1 => \N__14515\,
            in2 => \N__23678\,
            in3 => \N__16126\,
            lcout => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_2_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__19496\,
            in1 => \N__14474\,
            in2 => \N__15782\,
            in3 => \N__19695\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25209\,
            ce => 'H',
            sr => \N__24794\
        );

    \ppm_encoder_1.init_pulses_RNIANUS_2_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22137\,
            in1 => \N__22683\,
            in2 => \_gnd_net_\,
            in3 => \N__23682\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_2\,
            ltout => \ppm_encoder_1.un1_init_pulses_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI5V123_2_LC_8_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14465\,
            in3 => \N__14462\,
            lcout => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_11_LC_8_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19692\,
            in1 => \N__14456\,
            in2 => \N__19551\,
            in3 => \N__15890\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25204\,
            ce => 'H',
            sr => \N__24798\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_8_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22548\,
            in1 => \N__23686\,
            in2 => \_gnd_net_\,
            in3 => \N__22787\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23684\,
            in1 => \_gnd_net_\,
            in2 => \N__22823\,
            in3 => \N__22549\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_12_LC_8_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__19550\,
            in1 => \N__14435\,
            in2 => \N__19706\,
            in3 => \N__15881\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25204\,
            ce => 'H',
            sr => \N__24798\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_12_LC_8_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23687\,
            in1 => \_gnd_net_\,
            in2 => \N__22824\,
            in3 => \N__22458\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_8_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22459\,
            in1 => \N__23685\,
            in2 => \_gnd_net_\,
            in3 => \N__22786\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_14_LC_8_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19693\,
            in1 => \N__14567\,
            in2 => \N__19552\,
            in3 => \N__15857\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25204\,
            ce => 'H',
            sr => \N__24798\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_14_LC_8_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22317\,
            in1 => \N__23688\,
            in2 => \_gnd_net_\,
            in3 => \N__22791\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_8_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23692\,
            in1 => \N__16050\,
            in2 => \N__22826\,
            in3 => \N__16146\,
            lcout => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_15_LC_8_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__19576\,
            in1 => \N__14558\,
            in2 => \N__19702\,
            in3 => \N__15833\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25200\,
            ce => 'H',
            sr => \N__24801\
        );

    \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_8_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23690\,
            in1 => \_gnd_net_\,
            in2 => \N__22825\,
            in3 => \N__16051\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_18_LC_8_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19670\,
            in1 => \N__14546\,
            in2 => \N__19583\,
            in3 => \N__16154\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25200\,
            ce => 'H',
            sr => \N__24801\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_8_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22796\,
            in2 => \_gnd_net_\,
            in3 => \N__23691\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_10_LC_8_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__19669\,
            in1 => \N__19575\,
            in2 => \N__14663\,
            in3 => \N__15932\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25200\,
            ce => 'H',
            sr => \N__24801\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_8_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22017\,
            in1 => \N__22792\,
            in2 => \_gnd_net_\,
            in3 => \N__23689\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_16_LC_8_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19561\,
            in1 => \N__19667\,
            in2 => \N__14654\,
            in3 => \N__15824\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25196\,
            ce => 'H',
            sr => \N__24804\
        );

    \ppm_encoder_1.init_pulses_17_LC_8_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__19562\,
            in1 => \N__19668\,
            in2 => \N__15809\,
            in3 => \N__14645\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25196\,
            ce => 'H',
            sr => \N__24804\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_8_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23681\,
            in1 => \_gnd_net_\,
            in2 => \N__22821\,
            in3 => \N__16071\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_4_LC_8_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19666\,
            in1 => \N__14639\,
            in2 => \N__19580\,
            in3 => \N__15701\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25196\,
            ce => 'H',
            sr => \N__24804\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_4_LC_8_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19071\,
            in1 => \N__22772\,
            in2 => \_gnd_net_\,
            in3 => \N__23679\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_8_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23680\,
            in1 => \_gnd_net_\,
            in2 => \N__22820\,
            in3 => \N__19072\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_esr_6_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14627\,
            lcout => uart_pc_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25281\,
            ce => \N__14602\,
            sr => \N__14809\
        );

    \uart_frame_decoder.state_1_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__14671\,
            in1 => \N__14786\,
            in2 => \N__14780\,
            in3 => \N__23913\,
            lcout => \uart_frame_decoder.state_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25276\,
            ce => 'H',
            sr => \N__24742\
        );

    \uart_frame_decoder.state_1_10_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__23914\,
            in1 => \N__14672\,
            in2 => \N__14741\,
            in3 => \N__15318\,
            lcout => \uart_frame_decoder.state_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25276\,
            ce => 'H',
            sr => \N__24742\
        );

    \uart_frame_decoder.state_1_RNIF7PK_9_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14752\,
            in2 => \_gnd_net_\,
            in3 => \N__23821\,
            lcout => \uart_frame_decoder.source_offset4data_1_sqmuxa\,
            ltout => \uart_frame_decoder.source_offset4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNICKVT_9_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14732\,
            in3 => \N__24907\,
            lcout => \uart_frame_decoder.source_offset4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__16202\,
            in1 => \N__15039\,
            in2 => \_gnd_net_\,
            in3 => \N__15080\,
            lcout => \scaler_2.un2_source_data_0_cry_1_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNINMHJ_10_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23820\,
            in2 => \_gnd_net_\,
            in3 => \N__15315\,
            lcout => \uart_frame_decoder.state_1_RNINMHJZ0Z_10\,
            ltout => \uart_frame_decoder.state_1_RNINMHJZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_RNI8GDP1_2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__14729\,
            in1 => \N__14705\,
            in2 => \N__14675\,
            in3 => \N__16622\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_o2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_CH2data_esr_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21094\,
            lcout => \frame_decoder_CH2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25267\,
            ce => \N__17815\,
            sr => \N__24748\
        );

    \uart_frame_decoder.source_CH2data_esr_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20976\,
            lcout => \frame_decoder_CH2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25267\,
            ce => \N__17815\,
            sr => \N__24748\
        );

    \uart_frame_decoder.source_CH2data_esr_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20892\,
            lcout => \frame_decoder_CH2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25267\,
            ce => \N__17815\,
            sr => \N__24748\
        );

    \uart_frame_decoder.source_CH2data_esr_3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20809\,
            lcout => \frame_decoder_CH2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25267\,
            ce => \N__17815\,
            sr => \N__24748\
        );

    \uart_frame_decoder.source_CH2data_esr_4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20720\,
            lcout => \frame_decoder_CH2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25267\,
            ce => \N__17815\,
            sr => \N__24748\
        );

    \uart_frame_decoder.source_CH2data_esr_5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26355\,
            lcout => \frame_decoder_CH2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25267\,
            ce => \N__17815\,
            sr => \N__24748\
        );

    \uart_frame_decoder.source_CH2data_esr_6_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20606\,
            lcout => \frame_decoder_CH2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25267\,
            ce => \N__17815\,
            sr => \N__24748\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15038\,
            in2 => \N__15085\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14864\,
            in2 => \N__14858\,
            in3 => \N__14849\,
            lcout => \scaler_2.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_0\,
            carryout => \scaler_2.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14846\,
            in2 => \N__14840\,
            in3 => \N__14831\,
            lcout => \scaler_2.un3_source_data_0_cry_1_c_RNILSPH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_1\,
            carryout => \scaler_2.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14828\,
            in2 => \N__14822\,
            in3 => \N__14813\,
            lcout => \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_2\,
            carryout => \scaler_2.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14960\,
            in2 => \N__14954\,
            in3 => \N__14945\,
            lcout => \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_3\,
            carryout => \scaler_2.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14942\,
            in2 => \N__14936\,
            in3 => \N__14927\,
            lcout => \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_4\,
            carryout => \scaler_2.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14924\,
            in2 => \N__14918\,
            in3 => \N__14909\,
            lcout => \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_5\,
            carryout => \scaler_2.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17846\,
            in2 => \_gnd_net_\,
            in3 => \N__14906\,
            lcout => \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_6\,
            carryout => \scaler_2.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15134\,
            in2 => \N__21916\,
            in3 => \N__14903\,
            lcout => \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14900\,
            lcout => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI91PK_3_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23792\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14897\,
            lcout => \uart_frame_decoder.source_CH2data_1_sqmuxa\,
            ltout => \uart_frame_decoder.source_CH2data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI6EVT_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14867\,
            in3 => \N__24908\,
            lcout => \uart_frame_decoder.source_CH2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16669\,
            in2 => \_gnd_net_\,
            in3 => \N__21379\,
            lcout => \scaler_3.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.N_520_i_l_ofx_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17860\,
            in2 => \_gnd_net_\,
            in3 => \N__17837\,
            lcout => \scaler_2.N_520_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.source_data_1_esr_5_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16502\,
            in1 => \N__16592\,
            in2 => \_gnd_net_\,
            in3 => \N__16555\,
            lcout => scaler_1_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25246\,
            ce => \N__21142\,
            sr => \N__24760\
        );

    \scaler_2.source_data_1_esr_5_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16201\,
            in1 => \N__15081\,
            in2 => \_gnd_net_\,
            in3 => \N__15047\,
            lcout => scaler_2_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25246\,
            ce => \N__21142\,
            sr => \N__24760\
        );

    \scaler_3.source_data_1_esr_5_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21026\,
            in1 => \N__18069\,
            in2 => \_gnd_net_\,
            in3 => \N__16451\,
            lcout => scaler_3_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25246\,
            ce => \N__21142\,
            sr => \N__24760\
        );

    \scaler_1.source_data_1_4_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110010101100"
        )
    port map (
            in0 => \N__16587\,
            in1 => \N__15097\,
            in2 => \N__20176\,
            in3 => \N__16556\,
            lcout => scaler_1_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25241\,
            ce => 'H',
            sr => \N__24766\
        );

    \scaler_2.source_data_1_4_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__20167\,
            in1 => \N__15086\,
            in2 => \N__15016\,
            in3 => \N__15046\,
            lcout => scaler_2_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25241\,
            ce => 'H',
            sr => \N__24766\
        );

    \scaler_3.source_data_1_4_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__20168\,
            in1 => \N__21025\,
            in2 => \N__16460\,
            in3 => \N__14998\,
            lcout => scaler_3_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25241\,
            ce => 'H',
            sr => \N__24766\
        );

    \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__18074\,
            in1 => \N__16455\,
            in2 => \_gnd_net_\,
            in3 => \N__21018\,
            lcout => \scaler_3.un2_source_data_0_cry_1_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_4_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__20169\,
            in1 => \N__17900\,
            in2 => \N__14977\,
            in3 => \N__17936\,
            lcout => scaler_4_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25241\,
            ce => 'H',
            sr => \N__24766\
        );

    \ppm_encoder_1.rudder_10_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__20279\,
            in1 => \N__18110\,
            in2 => \N__25494\,
            in3 => \N__22042\,
            lcout => \ppm_encoder_1.rudderZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25233\,
            ce => 'H',
            sr => \N__24771\
        );

    \scaler_1.source_data_valid_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20165\,
            lcout => scaler_1_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25233\,
            ce => 'H',
            sr => \N__24771\
        );

    \uart_frame_decoder.source_data_valid_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__15281\,
            in1 => \N__15329\,
            in2 => \N__23787\,
            in3 => \N__20166\,
            lcout => pc_frame_decoder_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25233\,
            ce => 'H',
            sr => \N__24771\
        );

    \uart_frame_decoder.count8_cry_2_c_RNIU1C61_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__15328\,
            in1 => \N__24177\,
            in2 => \N__23818\,
            in3 => \N__15280\,
            lcout => \uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_rdy_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15268\,
            in2 => \_gnd_net_\,
            in3 => \N__15165\,
            lcout => uart_pc_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25233\,
            ce => 'H',
            sr => \N__24771\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16960\,
            in1 => \N__25777\,
            in2 => \_gnd_net_\,
            in3 => \N__16982\,
            lcout => \ppm_encoder_1.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_ctle_14_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25377\,
            in2 => \_gnd_net_\,
            in3 => \N__24911\,
            lcout => \ppm_encoder_1.scaler_1_dv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIG4JI2_11_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__16917\,
            in1 => \N__22531\,
            in2 => \N__18689\,
            in3 => \N__18769\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIALRT5_11_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__15923\,
            in1 => \_gnd_net_\,
            in2 => \N__15137\,
            in3 => \N__15362\,
            lcout => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI03DH2_11_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16936\,
            in1 => \N__15351\,
            in2 => \N__18543\,
            in3 => \N__18452\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25787\,
            in1 => \N__16918\,
            in2 => \_gnd_net_\,
            in3 => \N__16937\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26101\,
            in2 => \N__15356\,
            in3 => \N__15352\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_11_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__15353\,
            in1 => \N__25473\,
            in2 => \N__19217\,
            in3 => \N__19190\,
            lcout => \ppm_encoder_1.aileronZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25226\,
            ce => 'H',
            sr => \N__24778\
        );

    \ppm_encoder_1.throttle_RNIS5KK2_8_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__21640\,
            in1 => \N__18746\,
            in2 => \N__19037\,
            in3 => \N__18674\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIONI96_8_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__17423\,
            in1 => \_gnd_net_\,
            in2 => \N__15341\,
            in3 => \N__15338\,
            lcout => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNICKVN2_8_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__16849\,
            in1 => \N__16876\,
            in2 => \N__18451\,
            in3 => \N__18513\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIU7KK2_9_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__18673\,
            in1 => \N__19133\,
            in2 => \N__18768\,
            in3 => \N__25633\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNITSI96_9_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17372\,
            in2 => \N__15332\,
            in3 => \N__15482\,
            lcout => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIEMVN2_9_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011011101"
        )
    port map (
            in0 => \N__18512\,
            in1 => \N__16903\,
            in2 => \N__25656\,
            in3 => \N__18435\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_9_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__18251\,
            in1 => \N__18275\,
            in2 => \N__25528\,
            in3 => \N__25658\,
            lcout => \ppm_encoder_1.elevatorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25221\,
            ce => 'H',
            sr => \N__24783\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15475\,
            in1 => \N__15456\,
            in2 => \N__23590\,
            in3 => \N__25929\,
            lcout => \ppm_encoder_1.init_pulses_1_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__15436\,
            in1 => \N__15422\,
            in2 => \N__15407\,
            in3 => \N__18429\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__15616\,
            in1 => \N__24927\,
            in2 => \N__26100\,
            in3 => \N__23588\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23503\,
            in2 => \_gnd_net_\,
            in3 => \N__15403\,
            lcout => \ppm_encoder_1.init_pulses_3_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNI62ME2_4_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__15391\,
            in1 => \N__19054\,
            in2 => \N__15374\,
            in3 => \N__18643\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNI8CGI5_4_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__15737\,
            in1 => \_gnd_net_\,
            in2 => \N__15371\,
            in3 => \N__15368\,
            lcout => \ppm_encoder_1.aileron_esr_RNI8CGI5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.N_614_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22233\,
            in1 => \N__15615\,
            in2 => \N__25936\,
            in3 => \N__23499\,
            lcout => \ppm_encoder_1.init_pulses_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNI84ME2_5_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__15568\,
            in1 => \N__22081\,
            in2 => \N__18766\,
            in3 => \N__18656\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIDHGI5_5_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18916\,
            in2 => \N__15590\,
            in3 => \N__15587\,
            lcout => \ppm_encoder_1.aileron_esr_RNIDHGI5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__15580\,
            in1 => \N__18505\,
            in2 => \N__15545\,
            in3 => \N__18431\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25805\,
            in1 => \N__15581\,
            in2 => \_gnd_net_\,
            in3 => \N__15569\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26062\,
            in1 => \_gnd_net_\,
            in2 => \N__15557\,
            in3 => \N__15544\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_5_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15554\,
            lcout => \ppm_encoder_1.aileronZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25210\,
            ce => \N__21731\,
            sr => \N__24795\
        );

    \ppm_encoder_1.init_pulses_RNI8LUS_0_0_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15529\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15514\,
            in2 => \N__15503\,
            in3 => \N__15485\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15797\,
            in2 => \N__15791\,
            in3 => \N__15770\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15767\,
            in2 => \N__15752\,
            in3 => \N__15740\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15736\,
            in2 => \N__15713\,
            in3 => \N__15689\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18917\,
            in2 => \N__15686\,
            in3 => \N__15677\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17083\,
            in2 => \N__17057\,
            in3 => \N__15662\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17162\,
            in2 => \N__17188\,
            in3 => \N__15659\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17419\,
            in2 => \N__15656\,
            in3 => \N__15644\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_8\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17365\,
            in2 => \N__15641\,
            in3 => \N__15629\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17221\,
            in2 => \N__17204\,
            in3 => \N__15926\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15919\,
            in2 => \N__15902\,
            in3 => \N__15884\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17038\,
            in2 => \N__17024\,
            in3 => \N__15875\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17314\,
            in2 => \N__17297\,
            in3 => \N__15860\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18577\,
            in2 => \N__18563\,
            in3 => \N__15851\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15848\,
            in2 => \N__15842\,
            in3 => \N__15827\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15941\,
            in2 => \_gnd_net_\,
            in3 => \N__15818\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_16\,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15815\,
            in2 => \_gnd_net_\,
            in3 => \N__15800\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16094\,
            in2 => \_gnd_net_\,
            in3 => \N__16157\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_2_18_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__22813\,
            in1 => \N__16148\,
            in2 => \N__15978\,
            in3 => \N__23675\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__22910\,
            in1 => \N__26192\,
            in2 => \N__16037\,
            in3 => \N__22886\,
            lcout => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16088\,
            in2 => \_gnd_net_\,
            in3 => \N__24239\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_16_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__15955\,
            in1 => \N__17564\,
            in2 => \N__16019\,
            in3 => \N__23712\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25190\,
            ce => 'H',
            sr => \N__24808\
        );

    \ppm_encoder_1.pulses2count_17_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__23709\,
            in1 => \N__16016\,
            in2 => \N__16076\,
            in3 => \N__17551\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25190\,
            ce => 'H',
            sr => \N__24808\
        );

    \ppm_encoder_1.pulses2count_15_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__16055\,
            in1 => \N__16033\,
            in2 => \N__16018\,
            in3 => \N__23711\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25190\,
            ce => 'H',
            sr => \N__24808\
        );

    \ppm_encoder_1.pulses2count_18_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__23710\,
            in1 => \N__16017\,
            in2 => \N__15986\,
            in3 => \N__17531\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25190\,
            ce => 'H',
            sr => \N__24808\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__15954\,
            in1 => \N__22837\,
            in2 => \_gnd_net_\,
            in3 => \N__23708\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_offset4data_esr_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21107\,
            lcout => \frame_decoder_OFF4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25260\,
            ce => \N__20119\,
            sr => \N__24744\
        );

    \uart_frame_decoder.source_offset4data_esr_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20980\,
            lcout => \frame_decoder_OFF4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25260\,
            ce => \N__20119\,
            sr => \N__24744\
        );

    \uart_frame_decoder.source_offset4data_esr_7_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20535\,
            lcout => \frame_decoder_OFF4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25260\,
            ce => \N__20119\,
            sr => \N__24744\
        );

    \uart_frame_decoder.source_offset4data_esr_3_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20810\,
            lcout => \frame_decoder_OFF4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25260\,
            ce => \N__20119\,
            sr => \N__24744\
        );

    \uart_frame_decoder.source_offset4data_esr_5_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25260\,
            ce => \N__20119\,
            sr => \N__24744\
        );

    \uart_frame_decoder.source_offset4data_esr_6_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20613\,
            lcout => \frame_decoder_OFF4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25260\,
            ce => \N__20119\,
            sr => \N__24744\
        );

    \uart_frame_decoder.source_offset4data_esr_2_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20893\,
            lcout => \frame_decoder_OFF4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25260\,
            ce => \N__20119\,
            sr => \N__24744\
        );

    \scaler_2.un2_source_data_0_cry_1_c_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16190\,
            in2 => \N__16211\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_6_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16165\,
            in2 => \N__16200\,
            in3 => \N__16172\,
            lcout => scaler_2_data_6,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_1\,
            carryout => \scaler_2.un2_source_data_0_cry_2\,
            clk => \N__25253\,
            ce => \N__21137\,
            sr => \N__24749\
        );

    \scaler_2.source_data_1_esr_7_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16327\,
            in2 => \N__16169\,
            in3 => \N__16334\,
            lcout => scaler_2_data_7,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_2\,
            carryout => \scaler_2.un2_source_data_0_cry_3\,
            clk => \N__25253\,
            ce => \N__21137\,
            sr => \N__24749\
        );

    \scaler_2.source_data_1_esr_8_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16312\,
            in2 => \N__16331\,
            in3 => \N__16319\,
            lcout => scaler_2_data_8,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_3\,
            carryout => \scaler_2.un2_source_data_0_cry_4\,
            clk => \N__25253\,
            ce => \N__21137\,
            sr => \N__24749\
        );

    \scaler_2.source_data_1_esr_9_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16297\,
            in2 => \N__16316\,
            in3 => \N__16304\,
            lcout => scaler_2_data_9,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_4\,
            carryout => \scaler_2.un2_source_data_0_cry_5\,
            clk => \N__25253\,
            ce => \N__21137\,
            sr => \N__24749\
        );

    \scaler_2.source_data_1_esr_10_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16282\,
            in2 => \N__16301\,
            in3 => \N__16289\,
            lcout => scaler_2_data_10,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_5\,
            carryout => \scaler_2.un2_source_data_0_cry_6\,
            clk => \N__25253\,
            ce => \N__21137\,
            sr => \N__24749\
        );

    \scaler_2.source_data_1_esr_11_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16267\,
            in2 => \N__16286\,
            in3 => \N__16274\,
            lcout => scaler_2_data_11,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_6\,
            carryout => \scaler_2.un2_source_data_0_cry_7\,
            clk => \N__25253\,
            ce => \N__21137\,
            sr => \N__24749\
        );

    \scaler_2.source_data_1_esr_12_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16256\,
            in2 => \N__16271\,
            in3 => \N__16259\,
            lcout => scaler_2_data_12,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_7\,
            carryout => \scaler_2.un2_source_data_0_cry_8\,
            clk => \N__25253\,
            ce => \N__21137\,
            sr => \N__24749\
        );

    \scaler_2.source_data_1_esr_13_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16255\,
            in2 => \N__16241\,
            in3 => \N__16232\,
            lcout => scaler_2_data_13,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_9\,
            clk => \N__25248\,
            ce => \N__21138\,
            sr => \N__24753\
        );

    \scaler_2.source_data_1_esr_14_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16229\,
            lcout => scaler_2_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25248\,
            ce => \N__21138\,
            sr => \N__24753\
        );

    \scaler_4.source_data_1_esr_5_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20441\,
            in1 => \N__17896\,
            in2 => \_gnd_net_\,
            in3 => \N__17935\,
            lcout => scaler_4_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25248\,
            ce => \N__21138\,
            sr => \N__24753\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21017\,
            in2 => \N__16459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20909\,
            in2 => \N__16427\,
            in3 => \N__16415\,
            lcout => \scaler_3.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_0\,
            carryout => \scaler_3.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20822\,
            in2 => \N__16412\,
            in3 => \N__16400\,
            lcout => \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_1\,
            carryout => \scaler_3.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16397\,
            in2 => \N__20741\,
            in3 => \N__16388\,
            lcout => \scaler_3.un3_source_data_0_cry_2_c_RNIR08I\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_2\,
            carryout => \scaler_3.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16385\,
            in2 => \N__20645\,
            in3 => \N__16376\,
            lcout => \scaler_3.un3_source_data_0_cry_3_c_RNIU49I\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_3\,
            carryout => \scaler_3.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26279\,
            in2 => \N__16373\,
            in3 => \N__16358\,
            lcout => \scaler_3.un3_source_data_0_cry_4_c_RNI19AI\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_4\,
            carryout => \scaler_3.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16355\,
            in2 => \N__20549\,
            in3 => \N__16346\,
            lcout => \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_5\,
            carryout => \scaler_3.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16343\,
            in2 => \_gnd_net_\,
            in3 => \N__16337\,
            lcout => \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_6\,
            carryout => \scaler_3.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16658\,
            in2 => \N__21922\,
            in3 => \N__16700\,
            lcout => \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16697\,
            lcout => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_0_c_inv_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21893\,
            in1 => \N__16690\,
            in2 => \_gnd_net_\,
            in3 => \N__16610\,
            lcout => \uart_frame_decoder.count8_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.N_532_i_l_ofx_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16676\,
            in2 => \_gnd_net_\,
            in3 => \N__21383\,
            lcout => \scaler_3.N_532_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_0_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__16611\,
            in1 => \N__16652\,
            in2 => \_gnd_net_\,
            in3 => \N__16640\,
            lcout => \uart_frame_decoder.count8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__16511\,
            in1 => \N__16591\,
            in2 => \_gnd_net_\,
            in3 => \N__16554\,
            lcout => \scaler_1.un2_source_data_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un2_source_data_0_cry_1_c_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16503\,
            in2 => \N__16520\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \scaler_1.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.source_data_1_esr_6_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16474\,
            in2 => \N__16510\,
            in3 => \N__16481\,
            lcout => scaler_1_data_6,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_1\,
            carryout => \scaler_1.un2_source_data_0_cry_2\,
            clk => \N__25231\,
            ce => \N__21141\,
            sr => \N__24767\
        );

    \scaler_1.source_data_1_esr_7_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16822\,
            in2 => \N__16478\,
            in3 => \N__16463\,
            lcout => scaler_1_data_7,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_2\,
            carryout => \scaler_1.un2_source_data_0_cry_3\,
            clk => \N__25231\,
            ce => \N__21141\,
            sr => \N__24767\
        );

    \scaler_1.source_data_1_esr_8_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16804\,
            in2 => \N__16826\,
            in3 => \N__16811\,
            lcout => scaler_1_data_8,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_3\,
            carryout => \scaler_1.un2_source_data_0_cry_4\,
            clk => \N__25231\,
            ce => \N__21141\,
            sr => \N__24767\
        );

    \scaler_1.source_data_1_esr_9_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16786\,
            in2 => \N__16808\,
            in3 => \N__16793\,
            lcout => scaler_1_data_9,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_4\,
            carryout => \scaler_1.un2_source_data_0_cry_5\,
            clk => \N__25231\,
            ce => \N__21141\,
            sr => \N__24767\
        );

    \scaler_1.source_data_1_esr_10_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16768\,
            in2 => \N__16790\,
            in3 => \N__16775\,
            lcout => scaler_1_data_10,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_5\,
            carryout => \scaler_1.un2_source_data_0_cry_6\,
            clk => \N__25231\,
            ce => \N__21141\,
            sr => \N__24767\
        );

    \scaler_1.source_data_1_esr_11_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16750\,
            in2 => \N__16772\,
            in3 => \N__16757\,
            lcout => scaler_1_data_11,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_6\,
            carryout => \scaler_1.un2_source_data_0_cry_7\,
            clk => \N__25231\,
            ce => \N__21141\,
            sr => \N__24767\
        );

    \scaler_1.source_data_1_esr_12_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16735\,
            in2 => \N__16754\,
            in3 => \N__16739\,
            lcout => scaler_1_data_12,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_7\,
            carryout => \scaler_1.un2_source_data_0_cry_8\,
            clk => \N__25231\,
            ce => \N__21141\,
            sr => \N__24767\
        );

    \scaler_1.source_data_1_esr_13_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16736\,
            in2 => \N__16718\,
            in3 => \N__16706\,
            lcout => scaler_1_data_13,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \scaler_1.un2_source_data_0_cry_9\,
            clk => \N__25227\,
            ce => \N__21143\,
            sr => \N__24772\
        );

    \scaler_1.source_data_1_esr_14_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16703\,
            lcout => scaler_1_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25227\,
            ce => \N__21143\,
            sr => \N__24772\
        );

    \ppm_encoder_1.aileron_8_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__19325\,
            in1 => \N__19304\,
            in2 => \N__16850\,
            in3 => \N__25424\,
            lcout => \ppm_encoder_1.aileronZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25222\,
            ce => 'H',
            sr => \N__24776\
        );

    \ppm_encoder_1.rudder_8_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__25430\,
            in1 => \N__20351\,
            in2 => \N__19032\,
            in3 => \N__18125\,
            lcout => \ppm_encoder_1.rudderZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25222\,
            ce => 'H',
            sr => \N__24776\
        );

    \ppm_encoder_1.aileron_9_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__19285\,
            in1 => \N__19265\,
            in2 => \N__16904\,
            in3 => \N__25425\,
            lcout => \ppm_encoder_1.aileronZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25222\,
            ce => 'H',
            sr => \N__24776\
        );

    \ppm_encoder_1.elevator_11_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__18197\,
            in1 => \N__18176\,
            in2 => \N__25495\,
            in3 => \N__16935\,
            lcout => \ppm_encoder_1.elevatorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25222\,
            ce => 'H',
            sr => \N__24776\
        );

    \ppm_encoder_1.elevator_8_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__18284\,
            in1 => \N__18302\,
            in2 => \N__16877\,
            in3 => \N__25429\,
            lcout => \ppm_encoder_1.elevatorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25222\,
            ce => 'H',
            sr => \N__24776\
        );

    \ppm_encoder_1.throttle_11_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21275\,
            in1 => \N__21257\,
            in2 => \N__25496\,
            in3 => \N__16919\,
            lcout => \ppm_encoder_1.throttleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25222\,
            ce => 'H',
            sr => \N__24776\
        );

    \ppm_encoder_1.throttle_7_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__21299\,
            in1 => \N__21317\,
            in2 => \N__17147\,
            in3 => \N__25434\,
            lcout => \ppm_encoder_1.throttleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25222\,
            ce => 'H',
            sr => \N__24776\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26099\,
            in1 => \N__25610\,
            in2 => \_gnd_net_\,
            in3 => \N__16899\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_9_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25897\,
            in2 => \N__16880\,
            in3 => \N__19112\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25218\,
            ce => \N__26175\,
            sr => \N__24779\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25794\,
            in1 => \N__21641\,
            in2 => \_gnd_net_\,
            in3 => \N__16872\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26092\,
            in1 => \_gnd_net_\,
            in2 => \N__16853\,
            in3 => \N__16845\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_8_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25898\,
            in1 => \_gnd_net_\,
            in2 => \N__17048\,
            in3 => \N__18974\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25218\,
            ce => \N__26175\,
            sr => \N__24779\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26091\,
            in1 => \N__17126\,
            in2 => \_gnd_net_\,
            in3 => \N__17102\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNII6JI2_12_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16953\,
            in1 => \N__22444\,
            in2 => \N__18773\,
            in3 => \N__18690\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIFQRT5_12_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__17045\,
            in1 => \_gnd_net_\,
            in2 => \N__17027\,
            in3 => \N__17009\,
            lcout => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI25DH2_12_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16974\,
            in1 => \N__16992\,
            in2 => \N__18536\,
            in3 => \N__18444\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26073\,
            in1 => \N__17003\,
            in2 => \_gnd_net_\,
            in3 => \N__16993\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_12_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__16994\,
            in1 => \N__25477\,
            in2 => \N__19877\,
            in3 => \N__19850\,
            lcout => \ppm_encoder_1.aileronZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25212\,
            ce => 'H',
            sr => \N__24784\
        );

    \ppm_encoder_1.elevator_12_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__16975\,
            in1 => \N__18896\,
            in2 => \N__25529\,
            in3 => \N__18875\,
            lcout => \ppm_encoder_1.elevatorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25212\,
            ce => 'H',
            sr => \N__24784\
        );

    \ppm_encoder_1.throttle_12_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__21242\,
            in1 => \N__21218\,
            in2 => \N__16961\,
            in3 => \N__25481\,
            lcout => \ppm_encoder_1.throttleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25212\,
            ce => 'H',
            sr => \N__24784\
        );

    \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__19092\,
            in2 => \N__18765\,
            in3 => \N__18687\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIJII96_7_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17189\,
            in2 => \N__17165\,
            in3 => \N__17153\,
            lcout => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIAIVN2_7_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__17115\,
            in1 => \N__17097\,
            in2 => \N__18530\,
            in3 => \N__18430\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25747\,
            in1 => \N__17146\,
            in2 => \_gnd_net_\,
            in3 => \N__17116\,
            lcout => \ppm_encoder_1.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_7_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011100100"
        )
    port map (
            in0 => \N__25522\,
            in1 => \N__17117\,
            in2 => \N__18320\,
            in3 => \N__18341\,
            lcout => \ppm_encoder_1.elevatorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25206\,
            ce => 'H',
            sr => \N__24789\
        );

    \ppm_encoder_1.aileron_7_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011100100"
        )
    port map (
            in0 => \N__25521\,
            in1 => \N__17098\,
            in2 => \N__19364\,
            in3 => \N__19337\,
            lcout => \ppm_encoder_1.aileronZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25206\,
            ce => 'H',
            sr => \N__24789\
        );

    \ppm_encoder_1.rudder_7_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__19093\,
            in1 => \N__18140\,
            in2 => \N__20399\,
            in3 => \N__25523\,
            lcout => \ppm_encoder_1.rudderZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25206\,
            ce => 'H',
            sr => \N__24789\
        );

    \ppm_encoder_1.throttle_RNIO1KK2_6_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__17235\,
            in1 => \N__26233\,
            in2 => \N__18767\,
            in3 => \N__18672\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIEDI96_6_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__17084\,
            in1 => \_gnd_net_\,
            in2 => \N__17060\,
            in3 => \N__17255\,
            lcout => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI8GVN2_6_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__17247\,
            in1 => \N__22569\,
            in2 => \N__18531\,
            in3 => \N__18436\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25785\,
            in1 => \N__17236\,
            in2 => \_gnd_net_\,
            in3 => \N__17248\,
            lcout => \ppm_encoder_1.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_6_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__22570\,
            in1 => \N__25516\,
            in2 => \_gnd_net_\,
            in3 => \N__19396\,
            lcout => \ppm_encoder_1.aileronZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25202\,
            ce => 'H',
            sr => \N__24796\
        );

    \ppm_encoder_1.elevator_6_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__17249\,
            in1 => \_gnd_net_\,
            in2 => \N__25548\,
            in3 => \N__18362\,
            lcout => \ppm_encoder_1.elevatorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25202\,
            ce => 'H',
            sr => \N__24796\
        );

    \ppm_encoder_1.throttle_6_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__21335\,
            in1 => \N__25520\,
            in2 => \_gnd_net_\,
            in3 => \N__17237\,
            lcout => \ppm_encoder_1.throttleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25202\,
            ce => 'H',
            sr => \N__24796\
        );

    \ppm_encoder_1.throttle_RNIE2JI2_10_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__21550\,
            in1 => \N__22054\,
            in2 => \N__18781\,
            in3 => \N__18691\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI5GRT5_10_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17225\,
            in2 => \N__17207\,
            in3 => \N__17195\,
            lcout => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIU0DH2_10_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__17325\,
            in1 => \N__17337\,
            in2 => \N__18544\,
            in3 => \N__18454\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25786\,
            in1 => \N__21551\,
            in2 => \_gnd_net_\,
            in3 => \N__17326\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26011\,
            in2 => \N__17342\,
            in3 => \N__17338\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_10_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__17339\,
            in1 => \N__25554\,
            in2 => \N__19250\,
            in3 => \N__19226\,
            lcout => \ppm_encoder_1.aileronZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25198\,
            ce => 'H',
            sr => \N__24799\
        );

    \ppm_encoder_1.elevator_10_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__17327\,
            in1 => \N__18212\,
            in2 => \N__25559\,
            in3 => \N__18236\,
            lcout => \ppm_encoder_1.elevatorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25198\,
            ce => 'H',
            sr => \N__24799\
        );

    \ppm_encoder_1.throttle_RNIK8JI2_13_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__17265\,
            in1 => \N__22396\,
            in2 => \N__18785\,
            in3 => \N__18692\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIKVRT5_13_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__17315\,
            in1 => \_gnd_net_\,
            in2 => \N__17300\,
            in3 => \N__17288\,
            lcout => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI47DH2_13_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__25321\,
            in1 => \N__17277\,
            in2 => \N__18548\,
            in3 => \N__18455\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17278\,
            in1 => \N__25806\,
            in2 => \_gnd_net_\,
            in3 => \N__17266\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__25322\,
            in1 => \_gnd_net_\,
            in2 => \N__17282\,
            in3 => \N__26048\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_13_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011011110000100"
        )
    port map (
            in0 => \N__18836\,
            in1 => \N__25524\,
            in2 => \N__18863\,
            in3 => \N__17279\,
            lcout => \ppm_encoder_1.elevatorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25194\,
            ce => 'H',
            sr => \N__24802\
        );

    \ppm_encoder_1.throttle_13_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__21985\,
            in1 => \N__21788\,
            in2 => \N__25549\,
            in3 => \N__17267\,
            lcout => \ppm_encoder_1.throttleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25194\,
            ce => 'H',
            sr => \N__24802\
        );

    \ppm_encoder_1.init_pulses_8_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19671\,
            in1 => \N__17441\,
            in2 => \N__19581\,
            in3 => \N__17429\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25192\,
            ce => 'H',
            sr => \N__24805\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001101100"
        )
    port map (
            in0 => \N__23701\,
            in1 => \N__18988\,
            in2 => \N__22838\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__18987\,
            in1 => \N__22814\,
            in2 => \_gnd_net_\,
            in3 => \N__23699\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_9_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19672\,
            in1 => \N__17390\,
            in2 => \N__19582\,
            in3 => \N__17378\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25192\,
            ce => 'H',
            sr => \N__24805\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__22819\,
            in1 => \_gnd_net_\,
            in2 => \N__23714\,
            in3 => \N__19147\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19146\,
            in1 => \N__23700\,
            in2 => \_gnd_net_\,
            in3 => \N__22815\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_1_c_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20039\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_27_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17576\,
            in2 => \N__21955\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_0\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17570\,
            in2 => \N__21949\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_1\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19727\,
            in2 => \N__21952\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_2\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17582\,
            in2 => \N__21950\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_3\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17615\,
            in2 => \N__21953\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_4\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19733\,
            in2 => \N__21951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_5\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17477\,
            in2 => \N__21954\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_6\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17537\,
            in2 => \N__21965\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_28_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21964\,
            in2 => \N__17519\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_8\,
            carryout => \ppm_encoder_1.counter24_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17471\,
            lcout => \ppm_encoder_1.counter24_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__24348\,
            in1 => \N__17468\,
            in2 => \N__17453\,
            in3 => \N__24459\,
            lcout => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__17495\,
            in1 => \N__20096\,
            in2 => \N__19964\,
            in3 => \N__19898\,
            lcout => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23034\,
            in1 => \N__19784\,
            in2 => \N__19763\,
            in3 => \N__22992\,
            lcout => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__17563\,
            in1 => \N__22976\,
            in2 => \N__17552\,
            in3 => \N__22955\,
            lcout => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22933\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19933\,
            in1 => \N__19899\,
            in2 => \N__20102\,
            in3 => \N__21481\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_2_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19900\,
            in1 => \N__24023\,
            in2 => \N__19934\,
            in3 => \N__20100\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_2_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25893\,
            in1 => \N__17510\,
            in2 => \_gnd_net_\,
            in3 => \N__22118\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25185\,
            ce => \N__26177\,
            sr => \N__24811\
        );

    \ppm_encoder_1.pulses2count_esr_10_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17489\,
            in1 => \N__25894\,
            in2 => \_gnd_net_\,
            in3 => \N__22001\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25185\,
            ce => \N__26177\,
            sr => \N__24811\
        );

    \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__17621\,
            in1 => \N__24327\,
            in2 => \N__17591\,
            in3 => \N__24366\,
            lcout => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_11_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17606\,
            in1 => \N__25895\,
            in2 => \_gnd_net_\,
            in3 => \N__22361\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25185\,
            ce => \N__26177\,
            sr => \N__24811\
        );

    \uart_frame_decoder.source_CH4data_esr_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21108\,
            lcout => \frame_decoder_CH4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \uart_frame_decoder.source_CH4data_esr_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20981\,
            lcout => \frame_decoder_CH4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \uart_frame_decoder.source_CH4data_esr_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20872\,
            lcout => \frame_decoder_CH4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \uart_frame_decoder.source_CH4data_esr_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20788\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \uart_frame_decoder.source_CH4data_esr_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20721\,
            lcout => \frame_decoder_CH4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \uart_frame_decoder.source_CH4data_esr_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26332\,
            lcout => \frame_decoder_CH4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \uart_frame_decoder.source_CH4data_esr_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20621\,
            lcout => \frame_decoder_CH4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \uart_frame_decoder.source_CH4data_esr_7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20506\,
            lcout => \frame_decoder_CH4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25261\,
            ce => \N__17948\,
            sr => \N__24745\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17915\,
            in2 => \N__17895\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17723\,
            in2 => \N__17717\,
            in3 => \N__17708\,
            lcout => \scaler_4.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_0\,
            carryout => \scaler_4.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17705\,
            in2 => \N__17699\,
            in3 => \N__17690\,
            lcout => \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_1\,
            carryout => \scaler_4.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17687\,
            in2 => \N__17681\,
            in3 => \N__17672\,
            lcout => \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_2\,
            carryout => \scaler_4.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17669\,
            in2 => \N__20132\,
            in3 => \N__17663\,
            lcout => \scaler_4.un3_source_data_0_cry_3_c_RNI15MI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_3\,
            carryout => \scaler_4.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17660\,
            in2 => \N__17654\,
            in3 => \N__17645\,
            lcout => \scaler_4.un3_source_data_0_cry_4_c_RNI49NI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_4\,
            carryout => \scaler_4.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17642\,
            in2 => \N__17636\,
            in3 => \N__17627\,
            lcout => \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_5\,
            carryout => \scaler_4.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17732\,
            in2 => \_gnd_net_\,
            in3 => \N__17624\,
            lcout => \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_6\,
            carryout => \scaler_4.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17867\,
            in2 => \N__21948\,
            in3 => \N__17954\,
            lcout => \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17951\,
            lcout => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI8GVT_5_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__17773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24909\,
            lcout => \uart_frame_decoder.source_CH4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__20439\,
            in1 => \N__17925\,
            in2 => \_gnd_net_\,
            in3 => \N__17888\,
            lcout => \scaler_4.un2_source_data_0_cry_1_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.N_544_i_l_ofx_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17761\,
            in2 => \_gnd_net_\,
            in3 => \N__17747\,
            lcout => \scaler_4.N_544_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17861\,
            in2 => \_gnd_net_\,
            in3 => \N__17830\,
            lcout => \scaler_2.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_CH2data_esr_7_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20531\,
            lcout => \frame_decoder_CH2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25243\,
            ce => \N__17819\,
            sr => \N__24757\
        );

    \uart_frame_decoder.state_1_RNIB3PK_5_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17798\,
            in2 => \_gnd_net_\,
            in3 => \N__23822\,
            lcout => \uart_frame_decoder.source_CH4data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17762\,
            in2 => \_gnd_net_\,
            in3 => \N__17746\,
            lcout => \scaler_4.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18065\,
            in2 => \N__18089\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.source_data_1_esr_6_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18040\,
            in2 => \N__18073\,
            in3 => \N__18047\,
            lcout => scaler_3_data_6,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_1\,
            carryout => \scaler_3.un2_source_data_0_cry_2\,
            clk => \N__25236\,
            ce => \N__21139\,
            sr => \N__24761\
        );

    \scaler_3.source_data_1_esr_7_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18025\,
            in2 => \N__18044\,
            in3 => \N__18032\,
            lcout => scaler_3_data_7,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_2\,
            carryout => \scaler_3.un2_source_data_0_cry_3\,
            clk => \N__25236\,
            ce => \N__21139\,
            sr => \N__24761\
        );

    \scaler_3.source_data_1_esr_8_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18010\,
            in2 => \N__18029\,
            in3 => \N__18017\,
            lcout => scaler_3_data_8,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_3\,
            carryout => \scaler_3.un2_source_data_0_cry_4\,
            clk => \N__25236\,
            ce => \N__21139\,
            sr => \N__24761\
        );

    \scaler_3.source_data_1_esr_9_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17995\,
            in2 => \N__18014\,
            in3 => \N__18002\,
            lcout => scaler_3_data_9,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_4\,
            carryout => \scaler_3.un2_source_data_0_cry_5\,
            clk => \N__25236\,
            ce => \N__21139\,
            sr => \N__24761\
        );

    \scaler_3.source_data_1_esr_10_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17980\,
            in2 => \N__17999\,
            in3 => \N__17987\,
            lcout => scaler_3_data_10,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_5\,
            carryout => \scaler_3.un2_source_data_0_cry_6\,
            clk => \N__25236\,
            ce => \N__21139\,
            sr => \N__24761\
        );

    \scaler_3.source_data_1_esr_11_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17965\,
            in2 => \N__17984\,
            in3 => \N__17972\,
            lcout => scaler_3_data_11,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_6\,
            carryout => \scaler_3.un2_source_data_0_cry_7\,
            clk => \N__25236\,
            ce => \N__21139\,
            sr => \N__24761\
        );

    \scaler_3.source_data_1_esr_12_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18166\,
            in2 => \N__17969\,
            in3 => \N__17957\,
            lcout => scaler_3_data_12,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_7\,
            carryout => \scaler_3.un2_source_data_0_cry_8\,
            clk => \N__25236\,
            ce => \N__21139\,
            sr => \N__24761\
        );

    \scaler_3.source_data_1_esr_13_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18167\,
            in2 => \N__18155\,
            in3 => \N__18146\,
            lcout => scaler_3_data_13,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_9\,
            clk => \N__25232\,
            ce => \N__21140\,
            sr => \N__24768\
        );

    \scaler_3.source_data_1_esr_14_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18143\,
            lcout => scaler_3_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25232\,
            ce => \N__21140\,
            sr => \N__24768\
        );

    \ppm_encoder_1.un1_rudder_cry_6_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26257\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \ppm_encoder_1.un1_rudder_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20389\,
            in2 => \_gnd_net_\,
            in3 => \N__18128\,
            lcout => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_6\,
            carryout => \ppm_encoder_1.un1_rudder_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20347\,
            in2 => \_gnd_net_\,
            in3 => \N__18116\,
            lcout => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_7\,
            carryout => \ppm_encoder_1.un1_rudder_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20311\,
            in2 => \_gnd_net_\,
            in3 => \N__18113\,
            lcout => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_8\,
            carryout => \ppm_encoder_1.un1_rudder_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20278\,
            in2 => \_gnd_net_\,
            in3 => \N__18098\,
            lcout => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_9\,
            carryout => \ppm_encoder_1.un1_rudder_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21607\,
            in2 => \_gnd_net_\,
            in3 => \N__18095\,
            lcout => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_10\,
            carryout => \ppm_encoder_1.un1_rudder_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21523\,
            in2 => \_gnd_net_\,
            in3 => \N__18092\,
            lcout => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_11\,
            carryout => \ppm_encoder_1.un1_rudder_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21178\,
            in2 => \N__21920\,
            in3 => \N__18368\,
            lcout => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_12\,
            carryout => \ppm_encoder_1.un1_rudder_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_14_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21155\,
            in2 => \_gnd_net_\,
            in3 => \N__18365\,
            lcout => \ppm_encoder_1.rudderZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25223\,
            ce => \N__21738\,
            sr => \N__24777\
        );

    \ppm_encoder_1.un1_elevator_cry_6_c_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18358\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18337\,
            in2 => \_gnd_net_\,
            in3 => \N__18305\,
            lcout => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_6\,
            carryout => \ppm_encoder_1.un1_elevator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18301\,
            in2 => \_gnd_net_\,
            in3 => \N__18278\,
            lcout => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_7\,
            carryout => \ppm_encoder_1.un1_elevator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18268\,
            in2 => \_gnd_net_\,
            in3 => \N__18239\,
            lcout => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_8\,
            carryout => \ppm_encoder_1.un1_elevator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18229\,
            in2 => \_gnd_net_\,
            in3 => \N__18200\,
            lcout => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_9\,
            carryout => \ppm_encoder_1.un1_elevator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18196\,
            in3 => \N__18170\,
            lcout => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_10\,
            carryout => \ppm_encoder_1.un1_elevator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18892\,
            in2 => \_gnd_net_\,
            in3 => \N__18866\,
            lcout => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_11\,
            carryout => \ppm_encoder_1.un1_elevator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21849\,
            in2 => \N__18856\,
            in3 => \N__18824\,
            lcout => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_12\,
            carryout => \ppm_encoder_1.un1_elevator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_esr_14_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18821\,
            in2 => \_gnd_net_\,
            in3 => \N__18809\,
            lcout => \ppm_encoder_1.elevatorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25213\,
            ce => \N__21726\,
            sr => \N__24785\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24256\,
            in2 => \_gnd_net_\,
            in3 => \N__24028\,
            lcout => \ppm_encoder_1.N_143_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_13_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__21182\,
            in1 => \N__18806\,
            in2 => \N__25550\,
            in3 => \N__22389\,
            lcout => \ppm_encoder_1.rudderZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25207\,
            ce => 'H',
            sr => \N__24790\
        );

    \ppm_encoder_1.rudder_9_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__20315\,
            in1 => \N__25533\,
            in2 => \N__18797\,
            in3 => \N__19132\,
            lcout => \ppm_encoder_1.rudderZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25207\,
            ce => 'H',
            sr => \N__24790\
        );

    \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__22294\,
            in1 => \N__21757\,
            in2 => \N__18780\,
            in3 => \N__18688\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__18584\,
            in1 => \_gnd_net_\,
            in2 => \N__18566\,
            in3 => \N__18374\,
            lcout => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__22270\,
            in1 => \N__18535\,
            in2 => \N__19175\,
            in3 => \N__18453\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19174\,
            in1 => \N__25735\,
            in2 => \_gnd_net_\,
            in3 => \N__21758\,
            lcout => \ppm_encoder_1.N_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__23222\,
            in1 => \N__19154\,
            in2 => \N__23277\,
            in3 => \N__19131\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__19411\,
            in1 => \N__23220\,
            in2 => \N__19100\,
            in3 => \N__23258\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__23219\,
            in1 => \N__19079\,
            in2 => \N__23276\,
            in3 => \N__19058\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__19036\,
            in1 => \N__23259\,
            in2 => \N__19001\,
            in3 => \N__23221\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_3_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19703\,
            in1 => \N__18965\,
            in2 => \N__19566\,
            in3 => \N__18953\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25199\,
            ce => 'H',
            sr => \N__24800\
        );

    \ppm_encoder_1.init_pulses_5_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19704\,
            in1 => \N__18941\,
            in2 => \N__19567\,
            in3 => \N__18929\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25199\,
            ce => 'H',
            sr => \N__24800\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001101100"
        )
    port map (
            in0 => \N__22760\,
            in1 => \N__22098\,
            in2 => \N__23693\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23631\,
            in2 => \N__22103\,
            in3 => \N__22759\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_7_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__19705\,
            in1 => \N__19595\,
            in2 => \N__19568\,
            in3 => \N__19430\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25199\,
            ce => 'H',
            sr => \N__24800\
        );

    \ppm_encoder_1.un1_aileron_cry_6_c_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19397\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19360\,
            in2 => \_gnd_net_\,
            in3 => \N__19328\,
            lcout => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_6\,
            carryout => \ppm_encoder_1.un1_aileron_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19324\,
            in2 => \_gnd_net_\,
            in3 => \N__19289\,
            lcout => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_7\,
            carryout => \ppm_encoder_1.un1_aileron_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19286\,
            in2 => \_gnd_net_\,
            in3 => \N__19253\,
            lcout => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_8\,
            carryout => \ppm_encoder_1.un1_aileron_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19246\,
            in2 => \_gnd_net_\,
            in3 => \N__19220\,
            lcout => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_9\,
            carryout => \ppm_encoder_1.un1_aileron_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19213\,
            in2 => \_gnd_net_\,
            in3 => \N__19178\,
            lcout => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_10\,
            carryout => \ppm_encoder_1.un1_aileron_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19873\,
            in2 => \_gnd_net_\,
            in3 => \N__19838\,
            lcout => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_11\,
            carryout => \ppm_encoder_1.un1_aileron_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25591\,
            in2 => \N__21923\,
            in3 => \N__19835\,
            lcout => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_12\,
            carryout => \ppm_encoder_1.un1_aileron_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_14_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19832\,
            in2 => \_gnd_net_\,
            in3 => \N__19814\,
            lcout => \ppm_encoder_1.aileronZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25193\,
            ce => \N__21740\,
            sr => \N__24806\
        );

    \ppm_encoder_1.pulses2count_esr_4_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25884\,
            in1 => \N__19811\,
            in2 => \_gnd_net_\,
            in3 => \N__19796\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25189\,
            ce => \N__26171\,
            sr => \N__24807\
        );

    \ppm_encoder_1.pulses2count_esr_5_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19775\,
            in1 => \N__25885\,
            in2 => \_gnd_net_\,
            in3 => \N__22064\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25189\,
            ce => \N__26171\,
            sr => \N__24807\
        );

    \ppm_encoder_1.pulses2count_esr_13_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25883\,
            in1 => \N__19748\,
            in2 => \_gnd_net_\,
            in3 => \N__22373\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25189\,
            ce => \N__26171\,
            sr => \N__24807\
        );

    \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23318\,
            in1 => \N__22862\,
            in2 => \N__19742\,
            in3 => \N__24440\,
            lcout => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23017\,
            in1 => \N__23348\,
            in2 => \N__23372\,
            in3 => \N__23057\,
            lcout => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__26066\,
            in1 => \N__25781\,
            in2 => \_gnd_net_\,
            in3 => \N__20003\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_1_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25891\,
            in2 => \N__20051\,
            in3 => \N__23063\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25188\,
            ce => \N__26176\,
            sr => \N__24809\
        );

    \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__19925\,
            in1 => \N__24309\,
            in2 => \N__20048\,
            in3 => \N__20009\,
            lcout => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_0_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__23310\,
            in1 => \N__23225\,
            in2 => \_gnd_net_\,
            in3 => \N__20033\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25188\,
            ce => \N__26176\,
            sr => \N__24809\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20002\,
            in2 => \N__25804\,
            in3 => \N__26067\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_3_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22475\,
            in1 => \_gnd_net_\,
            in2 => \N__19967\,
            in3 => \N__25892\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25188\,
            ce => \N__26176\,
            sr => \N__24809\
        );

    \ppm_encoder_1.counter_0_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24311\,
            in2 => \N__19955\,
            in3 => \N__19954\,
            lcout => \ppm_encoder_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_28_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_0\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_1_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19932\,
            in2 => \_gnd_net_\,
            in3 => \N__19904\,
            lcout => \ppm_encoder_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_0\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_1\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_2_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19901\,
            in2 => \_gnd_net_\,
            in3 => \N__19880\,
            lcout => \ppm_encoder_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_1\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_2\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_3_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20101\,
            in2 => \_gnd_net_\,
            in3 => \N__20078\,
            lcout => \ppm_encoder_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_2\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_3\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_4_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22994\,
            in2 => \_gnd_net_\,
            in3 => \N__20075\,
            lcout => \ppm_encoder_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_3\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_4\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_5_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23036\,
            in2 => \_gnd_net_\,
            in3 => \N__20072\,
            lcout => \ppm_encoder_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_4\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_5\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_6_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23056\,
            in2 => \_gnd_net_\,
            in3 => \N__20069\,
            lcout => \ppm_encoder_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_5\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_6\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_7_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23016\,
            in2 => \_gnd_net_\,
            in3 => \N__20066\,
            lcout => \ppm_encoder_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_6\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_7\,
            clk => \N__25186\,
            ce => 'H',
            sr => \N__20201\
        );

    \ppm_encoder_1.counter_8_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24461\,
            in2 => \_gnd_net_\,
            in3 => \N__20063\,
            lcout => \ppm_encoder_1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_29_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_8\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_9_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24350\,
            in2 => \_gnd_net_\,
            in3 => \N__20060\,
            lcout => \ppm_encoder_1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_8\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_9\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_10_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24368\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => \ppm_encoder_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_9\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_10\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_11_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24331\,
            in2 => \_gnd_net_\,
            in3 => \N__20054\,
            lcout => \ppm_encoder_1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_10\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_11\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_12_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24439\,
            in2 => \_gnd_net_\,
            in3 => \N__20222\,
            lcout => \ppm_encoder_1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_11\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_12\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_13_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22861\,
            in2 => \_gnd_net_\,
            in3 => \N__20219\,
            lcout => \ppm_encoder_1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_12\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_13\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_14_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22882\,
            in2 => \_gnd_net_\,
            in3 => \N__20216\,
            lcout => \ppm_encoder_1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_13\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_14\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_15_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22906\,
            in2 => \_gnd_net_\,
            in3 => \N__20213\,
            lcout => \ppm_encoder_1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_14\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_15\,
            clk => \N__25184\,
            ce => 'H',
            sr => \N__20200\
        );

    \ppm_encoder_1.counter_16_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22954\,
            in2 => \_gnd_net_\,
            in3 => \N__20210\,
            lcout => \ppm_encoder_1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_30_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_16\,
            clk => \N__25183\,
            ce => 'H',
            sr => \N__20199\
        );

    \ppm_encoder_1.counter_17_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22975\,
            in2 => \_gnd_net_\,
            in3 => \N__20207\,
            lcout => \ppm_encoder_1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_16\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_17\,
            clk => \N__25183\,
            ce => 'H',
            sr => \N__20199\
        );

    \ppm_encoder_1.counter_18_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22932\,
            in2 => \_gnd_net_\,
            in3 => \N__20204\,
            lcout => \ppm_encoder_1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25183\,
            ce => 'H',
            sr => \N__20199\
        );

    \scaler_1.source_data_1_esr_ctle_14_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20186\,
            in2 => \_gnd_net_\,
            in3 => \N__24895\,
            lcout => pc_frame_decoder_dv_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_offset4data_esr_4_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20729\,
            lcout => \frame_decoder_OFF4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25247\,
            ce => \N__20123\,
            sr => \N__24754\
        );

    \scaler_4.un2_source_data_0_cry_1_c_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20432\,
            in2 => \N__20450\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_6_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20407\,
            in2 => \N__20440\,
            in3 => \N__20414\,
            lcout => scaler_4_data_6,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_1\,
            carryout => \scaler_4.un2_source_data_0_cry_2\,
            clk => \N__25242\,
            ce => \N__21135\,
            sr => \N__24758\
        );

    \scaler_4.source_data_1_esr_7_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20359\,
            in2 => \N__20411\,
            in3 => \N__20366\,
            lcout => scaler_4_data_7,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_2\,
            carryout => \scaler_4.un2_source_data_0_cry_3\,
            clk => \N__25242\,
            ce => \N__21135\,
            sr => \N__24758\
        );

    \scaler_4.source_data_1_esr_8_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20323\,
            in2 => \N__20363\,
            in3 => \N__20330\,
            lcout => scaler_4_data_8,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_3\,
            carryout => \scaler_4.un2_source_data_0_cry_4\,
            clk => \N__25242\,
            ce => \N__21135\,
            sr => \N__24758\
        );

    \scaler_4.source_data_1_esr_9_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20287\,
            in2 => \N__20327\,
            in3 => \N__20294\,
            lcout => scaler_4_data_9,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_4\,
            carryout => \scaler_4.un2_source_data_0_cry_5\,
            clk => \N__25242\,
            ce => \N__21135\,
            sr => \N__24758\
        );

    \scaler_4.source_data_1_esr_10_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20248\,
            in2 => \N__20291\,
            in3 => \N__20255\,
            lcout => scaler_4_data_10,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_5\,
            carryout => \scaler_4.un2_source_data_0_cry_6\,
            clk => \N__25242\,
            ce => \N__21135\,
            sr => \N__24758\
        );

    \scaler_4.source_data_1_esr_11_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20233\,
            in2 => \N__20252\,
            in3 => \N__20240\,
            lcout => scaler_4_data_11,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_6\,
            carryout => \scaler_4.un2_source_data_0_cry_7\,
            clk => \N__25242\,
            ce => \N__21135\,
            sr => \N__24758\
        );

    \scaler_4.source_data_1_esr_12_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21202\,
            in2 => \N__20237\,
            in3 => \N__20225\,
            lcout => scaler_4_data_12,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_7\,
            carryout => \scaler_4.un2_source_data_0_cry_8\,
            clk => \N__25242\,
            ce => \N__21135\,
            sr => \N__24758\
        );

    \scaler_4.source_data_1_esr_13_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21203\,
            in2 => \N__21191\,
            in3 => \N__21161\,
            lcout => scaler_4_data_13,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_9\,
            clk => \N__25234\,
            ce => \N__21136\,
            sr => \N__24762\
        );

    \scaler_4.source_data_1_esr_14_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21158\,
            lcout => scaler_4_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25234\,
            ce => \N__21136\,
            sr => \N__24762\
        );

    \uart_frame_decoder.source_CH3data_esr_0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21109\,
            lcout => \frame_decoder_CH3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25230\,
            ce => \N__26270\,
            sr => \N__24769\
        );

    \uart_frame_decoder.source_CH3data_esr_1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20990\,
            lcout => \frame_decoder_CH3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25230\,
            ce => \N__26270\,
            sr => \N__24769\
        );

    \uart_frame_decoder.source_CH3data_esr_2_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20900\,
            lcout => \frame_decoder_CH3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25230\,
            ce => \N__26270\,
            sr => \N__24769\
        );

    \uart_frame_decoder.source_CH3data_esr_3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20808\,
            lcout => \frame_decoder_CH3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25230\,
            ce => \N__26270\,
            sr => \N__24769\
        );

    \uart_frame_decoder.source_CH3data_esr_4_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20728\,
            lcout => \frame_decoder_CH3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25230\,
            ce => \N__26270\,
            sr => \N__24769\
        );

    \uart_frame_decoder.source_CH3data_esr_6_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20631\,
            lcout => \frame_decoder_CH3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25230\,
            ce => \N__26270\,
            sr => \N__24769\
        );

    \uart_frame_decoder.source_CH3data_esr_7_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20537\,
            lcout => \frame_decoder_CH3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25230\,
            ce => \N__26270\,
            sr => \N__24769\
        );

    \uart_frame_decoder.state_1_RNI80PK_2_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23866\,
            in2 => \_gnd_net_\,
            in3 => \N__23788\,
            lcout => \uart_frame_decoder.source_CH1data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_c_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21334\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21316\,
            in2 => \_gnd_net_\,
            in3 => \N__21287\,
            lcout => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_6\,
            carryout => \ppm_encoder_1.un1_throttle_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21655\,
            in2 => \_gnd_net_\,
            in3 => \N__21284\,
            lcout => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_7\,
            carryout => \ppm_encoder_1.un1_throttle_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21400\,
            in2 => \_gnd_net_\,
            in3 => \N__21281\,
            lcout => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_8\,
            carryout => \ppm_encoder_1.un1_throttle_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21568\,
            in2 => \_gnd_net_\,
            in3 => \N__21278\,
            lcout => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_9\,
            carryout => \ppm_encoder_1.un1_throttle_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21274\,
            in2 => \_gnd_net_\,
            in3 => \N__21245\,
            lcout => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_10\,
            carryout => \ppm_encoder_1.un1_throttle_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21238\,
            in3 => \N__21206\,
            lcout => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_11\,
            carryout => \ppm_encoder_1.un1_throttle_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21986\,
            in2 => \N__21921\,
            in3 => \N__21773\,
            lcout => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_12\,
            carryout => \ppm_encoder_1.un1_throttle_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_14_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21770\,
            in2 => \_gnd_net_\,
            in3 => \N__21761\,
            lcout => \ppm_encoder_1.throttleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25217\,
            ce => \N__21730\,
            sr => \N__24780\
        );

    \ppm_encoder_1.throttle_8_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21668\,
            in1 => \N__21659\,
            in2 => \N__25547\,
            in3 => \N__21633\,
            lcout => \ppm_encoder_1.throttleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25211\,
            ce => 'H',
            sr => \N__24786\
        );

    \ppm_encoder_1.rudder_11_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21611\,
            in1 => \N__21590\,
            in2 => \N__25544\,
            in3 => \N__22530\,
            lcout => \ppm_encoder_1.rudderZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25205\,
            ce => 'H',
            sr => \N__24791\
        );

    \ppm_encoder_1.throttle_10_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__21581\,
            in1 => \N__21572\,
            in2 => \N__21549\,
            in3 => \N__25505\,
            lcout => \ppm_encoder_1.throttleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25205\,
            ce => 'H',
            sr => \N__24791\
        );

    \ppm_encoder_1.rudder_12_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21527\,
            in1 => \N__21503\,
            in2 => \N__25545\,
            in3 => \N__22443\,
            lcout => \ppm_encoder_1.rudderZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25201\,
            ce => 'H',
            sr => \N__24797\
        );

    \ppm_encoder_1.ppm_output_reg_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111101000100"
        )
    port map (
            in0 => \N__24380\,
            in1 => \N__21491\,
            in2 => \N__21485\,
            in3 => \N__21424\,
            lcout => ppm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25201\,
            ce => 'H',
            sr => \N__24797\
        );

    \ppm_encoder_1.throttle_9_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21413\,
            in1 => \N__21404\,
            in2 => \N__25546\,
            in3 => \N__25632\,
            lcout => \ppm_encoder_1.throttleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25201\,
            ce => 'H',
            sr => \N__24797\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__25732\,
            in1 => \N__22249\,
            in2 => \_gnd_net_\,
            in3 => \N__22194\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_7\,
            ltout => \ppm_encoder_1.pulses2count_9_sn_N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__23223\,
            in1 => \N__22331\,
            in2 => \N__22301\,
            in3 => \N__22298\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26031\,
            in1 => \N__22277\,
            in2 => \_gnd_net_\,
            in3 => \N__22271\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__25733\,
            in1 => \N__24928\,
            in2 => \N__26065\,
            in3 => \N__23698\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__22253\,
            in1 => \N__25734\,
            in2 => \_gnd_net_\,
            in3 => \N__22199\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\,
            ltout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__23251\,
            in1 => \N__23211\,
            in2 => \N__22148\,
            in3 => \N__22145\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__23212\,
            in1 => \N__22102\,
            in2 => \N__23275\,
            in3 => \N__22085\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__22055\,
            in1 => \N__23206\,
            in2 => \N__23299\,
            in3 => \N__22028\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110111010"
        )
    port map (
            in0 => \N__24929\,
            in1 => \N__22841\,
            in2 => \N__23713\,
            in3 => \N__25979\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25978\,
            in1 => \N__22592\,
            in2 => \_gnd_net_\,
            in3 => \N__22580\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23205\,
            in1 => \N__22556\,
            in2 => \_gnd_net_\,
            in3 => \N__22535\,
            lcout => \ppm_encoder_1.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__23308\,
            in1 => \N__23209\,
            in2 => \N__23116\,
            in3 => \N__22502\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23207\,
            in1 => \N__22463\,
            in2 => \_gnd_net_\,
            in3 => \N__22445\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__23109\,
            in1 => \_gnd_net_\,
            in2 => \N__22421\,
            in3 => \N__23301\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101001111"
        )
    port map (
            in0 => \N__23208\,
            in1 => \N__22418\,
            in2 => \N__23311\,
            in3 => \N__22400\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__23108\,
            in1 => \N__23300\,
            in2 => \_gnd_net_\,
            in3 => \N__22367\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101001111"
        )
    port map (
            in0 => \N__23210\,
            in1 => \N__22349\,
            in2 => \N__23312\,
            in3 => \N__26234\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24917\,
            in2 => \_gnd_net_\,
            in3 => \N__23694\,
            lcout => \ppm_encoder_1.N_614_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_7_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23396\,
            in1 => \N__25863\,
            in2 => \_gnd_net_\,
            in3 => \N__23384\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25187\,
            ce => \N__26160\,
            sr => \N__24810\
        );

    \ppm_encoder_1.pulses2count_esr_6_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25862\,
            in1 => \N__23363\,
            in2 => \_gnd_net_\,
            in3 => \N__23354\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25187\,
            ce => \N__26160\,
            sr => \N__24810\
        );

    \ppm_encoder_1.pulses2count_esr_12_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25861\,
            in1 => \N__23342\,
            in2 => \_gnd_net_\,
            in3 => \N__23324\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25187\,
            ce => \N__26160\,
            sr => \N__24810\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__23309\,
            in1 => \N__23224\,
            in2 => \N__23120\,
            in3 => \N__23090\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIUS1G_4_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23055\,
            in1 => \N__23035\,
            in2 => \N__23018\,
            in3 => \N__22993\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNI637H_18_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22974\,
            in1 => \N__22953\,
            in2 => \N__22934\,
            in3 => \N__22905\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIDBJ8_13_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22881\,
            in2 => \_gnd_net_\,
            in3 => \N__22860\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIAEV01_8_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__24467\,
            in1 => \N__24460\,
            in2 => \N__24443\,
            in3 => \N__24438\,
            lcout => \ppm_encoder_1.N_148_17\,
            ltout => \ppm_encoder_1.N_148_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24292\,
            in1 => \N__24406\,
            in2 => \N__24419\,
            in3 => \N__24416\,
            lcout => \ppm_encoder_1.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_1_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24407\,
            in1 => \N__24398\,
            in2 => \N__24392\,
            in3 => \N__24293\,
            lcout => \ppm_encoder_1.N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIK1KG_0_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24367\,
            in1 => \N__24349\,
            in2 => \N__24332\,
            in3 => \N__24310\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__24268\,
            in1 => \N__24252\,
            in2 => \N__24203\,
            in3 => \N__24029\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_2_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23963\,
            in1 => \N__23942\,
            in2 => \N__23867\,
            in3 => \N__23915\,
            lcout => \uart_frame_decoder.state_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25249\,
            ce => 'H',
            sr => \N__24763\
        );

    \uart_frame_decoder.state_1_RNIA2PK_4_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23846\,
            in2 => \_gnd_net_\,
            in3 => \N__23819\,
            lcout => \uart_frame_decoder.source_CH3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI7FVT_4_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24910\,
            lcout => \uart_frame_decoder.source_CH3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_CH3data_esr_5_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26362\,
            lcout => \frame_decoder_CH3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25237\,
            ce => \N__26269\,
            sr => \N__24773\
        );

    \ppm_encoder_1.rudder_6_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__25512\,
            in1 => \N__26258\,
            in2 => \_gnd_net_\,
            in3 => \N__26226\,
            lcout => \ppm_encoder_1.rudderZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25219\,
            ce => 'H',
            sr => \N__24792\
        );

    \ppm_encoder_1.pulses2count_esr_14_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26204\,
            in1 => \N__25896\,
            in2 => \_gnd_net_\,
            in3 => \N__26198\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25203\,
            ce => \N__26167\,
            sr => \N__24803\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__26064\,
            in1 => \N__25795\,
            in2 => \_gnd_net_\,
            in3 => \N__25943\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25796\,
            in1 => \N__25657\,
            in2 => \_gnd_net_\,
            in3 => \N__25634\,
            lcout => \ppm_encoder_1.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_13_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__25598\,
            in1 => \N__25571\,
            in2 => \N__25558\,
            in3 => \N__25320\,
            lcout => \ppm_encoder_1.aileronZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25195\,
            ce => 'H',
            sr => \N__24812\
        );
end \INTERFACE\;
