// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 18 2019 12:11:38

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_pc,
    debug_CH5_31B,
    debug_CH3_20A,
    debug_CH0_16A,
    uart_input_drone,
    ppm_output,
    debug_CH6_5B,
    debug_CH2_18A,
    debug_CH4_2A,
    debug_CH1_0A,
    clk_system);

    input uart_input_pc;
    output debug_CH5_31B;
    output debug_CH3_20A;
    output debug_CH0_16A;
    input uart_input_drone;
    output ppm_output;
    output debug_CH6_5B;
    output debug_CH2_18A;
    output debug_CH4_2A;
    output debug_CH1_0A;
    input clk_system;

    wire N__59697;
    wire N__59683;
    wire N__59682;
    wire N__59681;
    wire N__59674;
    wire N__59673;
    wire N__59672;
    wire N__59665;
    wire N__59664;
    wire N__59663;
    wire N__59656;
    wire N__59655;
    wire N__59654;
    wire N__59647;
    wire N__59646;
    wire N__59645;
    wire N__59638;
    wire N__59637;
    wire N__59636;
    wire N__59629;
    wire N__59628;
    wire N__59627;
    wire N__59620;
    wire N__59619;
    wire N__59618;
    wire N__59611;
    wire N__59610;
    wire N__59609;
    wire N__59602;
    wire N__59601;
    wire N__59600;
    wire N__59583;
    wire N__59580;
    wire N__59577;
    wire N__59574;
    wire N__59573;
    wire N__59572;
    wire N__59569;
    wire N__59566;
    wire N__59563;
    wire N__59560;
    wire N__59557;
    wire N__59554;
    wire N__59551;
    wire N__59546;
    wire N__59543;
    wire N__59538;
    wire N__59535;
    wire N__59532;
    wire N__59529;
    wire N__59528;
    wire N__59527;
    wire N__59520;
    wire N__59517;
    wire N__59514;
    wire N__59511;
    wire N__59508;
    wire N__59505;
    wire N__59502;
    wire N__59501;
    wire N__59500;
    wire N__59497;
    wire N__59492;
    wire N__59487;
    wire N__59484;
    wire N__59481;
    wire N__59478;
    wire N__59475;
    wire N__59472;
    wire N__59469;
    wire N__59466;
    wire N__59463;
    wire N__59460;
    wire N__59459;
    wire N__59458;
    wire N__59455;
    wire N__59452;
    wire N__59449;
    wire N__59446;
    wire N__59443;
    wire N__59436;
    wire N__59433;
    wire N__59430;
    wire N__59427;
    wire N__59426;
    wire N__59425;
    wire N__59418;
    wire N__59415;
    wire N__59412;
    wire N__59409;
    wire N__59406;
    wire N__59403;
    wire N__59400;
    wire N__59397;
    wire N__59396;
    wire N__59395;
    wire N__59392;
    wire N__59387;
    wire N__59382;
    wire N__59379;
    wire N__59376;
    wire N__59373;
    wire N__59370;
    wire N__59367;
    wire N__59364;
    wire N__59361;
    wire N__59360;
    wire N__59359;
    wire N__59352;
    wire N__59349;
    wire N__59346;
    wire N__59343;
    wire N__59340;
    wire N__59337;
    wire N__59336;
    wire N__59335;
    wire N__59334;
    wire N__59333;
    wire N__59332;
    wire N__59331;
    wire N__59330;
    wire N__59329;
    wire N__59328;
    wire N__59327;
    wire N__59326;
    wire N__59325;
    wire N__59324;
    wire N__59323;
    wire N__59322;
    wire N__59321;
    wire N__59320;
    wire N__59319;
    wire N__59318;
    wire N__59317;
    wire N__59316;
    wire N__59315;
    wire N__59314;
    wire N__59313;
    wire N__59312;
    wire N__59311;
    wire N__59310;
    wire N__59309;
    wire N__59308;
    wire N__59307;
    wire N__59306;
    wire N__59305;
    wire N__59304;
    wire N__59303;
    wire N__59302;
    wire N__59301;
    wire N__59300;
    wire N__59299;
    wire N__59298;
    wire N__59297;
    wire N__59296;
    wire N__59295;
    wire N__59294;
    wire N__59293;
    wire N__59292;
    wire N__59291;
    wire N__59290;
    wire N__59289;
    wire N__59288;
    wire N__59287;
    wire N__59286;
    wire N__59285;
    wire N__59284;
    wire N__59283;
    wire N__59282;
    wire N__59281;
    wire N__59280;
    wire N__59279;
    wire N__59278;
    wire N__59277;
    wire N__59276;
    wire N__59275;
    wire N__59274;
    wire N__59273;
    wire N__59272;
    wire N__59271;
    wire N__59270;
    wire N__59269;
    wire N__59268;
    wire N__59267;
    wire N__59266;
    wire N__59265;
    wire N__59264;
    wire N__59263;
    wire N__59262;
    wire N__59261;
    wire N__59260;
    wire N__59259;
    wire N__59258;
    wire N__59257;
    wire N__59256;
    wire N__59255;
    wire N__59254;
    wire N__59253;
    wire N__59252;
    wire N__59251;
    wire N__59250;
    wire N__59249;
    wire N__59248;
    wire N__59247;
    wire N__59246;
    wire N__59245;
    wire N__59244;
    wire N__59243;
    wire N__59242;
    wire N__59241;
    wire N__59240;
    wire N__59239;
    wire N__59238;
    wire N__59237;
    wire N__59236;
    wire N__59235;
    wire N__59234;
    wire N__59233;
    wire N__59232;
    wire N__59231;
    wire N__59230;
    wire N__59229;
    wire N__59228;
    wire N__59227;
    wire N__59226;
    wire N__59225;
    wire N__59224;
    wire N__59223;
    wire N__59222;
    wire N__59221;
    wire N__59220;
    wire N__59219;
    wire N__59218;
    wire N__59217;
    wire N__59216;
    wire N__59215;
    wire N__59214;
    wire N__59213;
    wire N__59212;
    wire N__59211;
    wire N__59210;
    wire N__59209;
    wire N__59208;
    wire N__59207;
    wire N__59206;
    wire N__59205;
    wire N__59204;
    wire N__59203;
    wire N__59202;
    wire N__59201;
    wire N__59200;
    wire N__59199;
    wire N__59198;
    wire N__59197;
    wire N__59196;
    wire N__59195;
    wire N__59194;
    wire N__59193;
    wire N__59192;
    wire N__59191;
    wire N__59190;
    wire N__59189;
    wire N__59188;
    wire N__59187;
    wire N__59186;
    wire N__59185;
    wire N__59184;
    wire N__59183;
    wire N__59182;
    wire N__59181;
    wire N__59180;
    wire N__59179;
    wire N__59178;
    wire N__59177;
    wire N__59176;
    wire N__59175;
    wire N__59174;
    wire N__59173;
    wire N__59172;
    wire N__59171;
    wire N__59170;
    wire N__59169;
    wire N__59168;
    wire N__59167;
    wire N__59166;
    wire N__59165;
    wire N__59164;
    wire N__59163;
    wire N__59162;
    wire N__59161;
    wire N__59160;
    wire N__59159;
    wire N__59158;
    wire N__59157;
    wire N__59156;
    wire N__59155;
    wire N__59154;
    wire N__59153;
    wire N__59152;
    wire N__59151;
    wire N__59150;
    wire N__59149;
    wire N__59148;
    wire N__59147;
    wire N__59146;
    wire N__59145;
    wire N__59144;
    wire N__59143;
    wire N__59142;
    wire N__59141;
    wire N__59140;
    wire N__59139;
    wire N__59138;
    wire N__59137;
    wire N__59136;
    wire N__59135;
    wire N__59134;
    wire N__59133;
    wire N__59132;
    wire N__59131;
    wire N__59130;
    wire N__59129;
    wire N__59128;
    wire N__59127;
    wire N__59126;
    wire N__59125;
    wire N__59124;
    wire N__59123;
    wire N__59122;
    wire N__59121;
    wire N__59120;
    wire N__59119;
    wire N__59118;
    wire N__59117;
    wire N__59116;
    wire N__59115;
    wire N__59114;
    wire N__59113;
    wire N__59112;
    wire N__59111;
    wire N__59110;
    wire N__59109;
    wire N__59108;
    wire N__59107;
    wire N__59106;
    wire N__59105;
    wire N__59104;
    wire N__59103;
    wire N__59102;
    wire N__59101;
    wire N__59100;
    wire N__59099;
    wire N__59098;
    wire N__59097;
    wire N__59096;
    wire N__59095;
    wire N__59094;
    wire N__59093;
    wire N__59092;
    wire N__59091;
    wire N__59090;
    wire N__59089;
    wire N__59088;
    wire N__59087;
    wire N__59086;
    wire N__59085;
    wire N__59084;
    wire N__59083;
    wire N__59082;
    wire N__59081;
    wire N__59080;
    wire N__59079;
    wire N__59078;
    wire N__59077;
    wire N__59076;
    wire N__59075;
    wire N__59074;
    wire N__58545;
    wire N__58542;
    wire N__58539;
    wire N__58538;
    wire N__58537;
    wire N__58536;
    wire N__58535;
    wire N__58534;
    wire N__58531;
    wire N__58528;
    wire N__58525;
    wire N__58524;
    wire N__58523;
    wire N__58520;
    wire N__58517;
    wire N__58514;
    wire N__58511;
    wire N__58508;
    wire N__58507;
    wire N__58504;
    wire N__58503;
    wire N__58502;
    wire N__58499;
    wire N__58496;
    wire N__58495;
    wire N__58494;
    wire N__58491;
    wire N__58486;
    wire N__58483;
    wire N__58480;
    wire N__58477;
    wire N__58474;
    wire N__58471;
    wire N__58468;
    wire N__58465;
    wire N__58462;
    wire N__58459;
    wire N__58456;
    wire N__58455;
    wire N__58450;
    wire N__58449;
    wire N__58446;
    wire N__58443;
    wire N__58440;
    wire N__58435;
    wire N__58432;
    wire N__58423;
    wire N__58420;
    wire N__58417;
    wire N__58414;
    wire N__58411;
    wire N__58408;
    wire N__58405;
    wire N__58402;
    wire N__58395;
    wire N__58392;
    wire N__58389;
    wire N__58386;
    wire N__58383;
    wire N__58378;
    wire N__58375;
    wire N__58370;
    wire N__58359;
    wire N__58358;
    wire N__58357;
    wire N__58356;
    wire N__58355;
    wire N__58354;
    wire N__58353;
    wire N__58352;
    wire N__58351;
    wire N__58350;
    wire N__58349;
    wire N__58348;
    wire N__58347;
    wire N__58346;
    wire N__58345;
    wire N__58344;
    wire N__58343;
    wire N__58342;
    wire N__58341;
    wire N__58340;
    wire N__58339;
    wire N__58338;
    wire N__58337;
    wire N__58336;
    wire N__58335;
    wire N__58334;
    wire N__58333;
    wire N__58332;
    wire N__58331;
    wire N__58330;
    wire N__58329;
    wire N__58328;
    wire N__58327;
    wire N__58326;
    wire N__58325;
    wire N__58324;
    wire N__58323;
    wire N__58322;
    wire N__58321;
    wire N__58320;
    wire N__58319;
    wire N__58314;
    wire N__58305;
    wire N__58300;
    wire N__58295;
    wire N__58286;
    wire N__58281;
    wire N__58276;
    wire N__58265;
    wire N__58262;
    wire N__58257;
    wire N__58252;
    wire N__58247;
    wire N__58232;
    wire N__58229;
    wire N__58226;
    wire N__58223;
    wire N__58220;
    wire N__58219;
    wire N__58218;
    wire N__58217;
    wire N__58216;
    wire N__58215;
    wire N__58214;
    wire N__58213;
    wire N__58212;
    wire N__58211;
    wire N__58210;
    wire N__58209;
    wire N__58208;
    wire N__58207;
    wire N__58206;
    wire N__58205;
    wire N__58204;
    wire N__58203;
    wire N__58202;
    wire N__58201;
    wire N__58200;
    wire N__58199;
    wire N__58198;
    wire N__58197;
    wire N__58196;
    wire N__58195;
    wire N__58194;
    wire N__58193;
    wire N__58192;
    wire N__58191;
    wire N__58190;
    wire N__58189;
    wire N__58188;
    wire N__58187;
    wire N__58186;
    wire N__58185;
    wire N__58184;
    wire N__58183;
    wire N__58182;
    wire N__58181;
    wire N__58180;
    wire N__58179;
    wire N__58176;
    wire N__58173;
    wire N__58170;
    wire N__58167;
    wire N__58164;
    wire N__58161;
    wire N__58158;
    wire N__58155;
    wire N__58152;
    wire N__58149;
    wire N__58146;
    wire N__58143;
    wire N__58140;
    wire N__58137;
    wire N__58134;
    wire N__58131;
    wire N__58128;
    wire N__58011;
    wire N__58008;
    wire N__58005;
    wire N__58004;
    wire N__58001;
    wire N__57998;
    wire N__57997;
    wire N__57994;
    wire N__57991;
    wire N__57988;
    wire N__57981;
    wire N__57980;
    wire N__57977;
    wire N__57974;
    wire N__57969;
    wire N__57966;
    wire N__57965;
    wire N__57964;
    wire N__57963;
    wire N__57962;
    wire N__57961;
    wire N__57960;
    wire N__57959;
    wire N__57958;
    wire N__57957;
    wire N__57956;
    wire N__57955;
    wire N__57954;
    wire N__57953;
    wire N__57952;
    wire N__57951;
    wire N__57950;
    wire N__57949;
    wire N__57948;
    wire N__57909;
    wire N__57906;
    wire N__57903;
    wire N__57902;
    wire N__57901;
    wire N__57900;
    wire N__57897;
    wire N__57896;
    wire N__57895;
    wire N__57894;
    wire N__57891;
    wire N__57890;
    wire N__57889;
    wire N__57888;
    wire N__57887;
    wire N__57886;
    wire N__57885;
    wire N__57884;
    wire N__57883;
    wire N__57882;
    wire N__57881;
    wire N__57880;
    wire N__57879;
    wire N__57878;
    wire N__57877;
    wire N__57876;
    wire N__57875;
    wire N__57872;
    wire N__57871;
    wire N__57870;
    wire N__57869;
    wire N__57868;
    wire N__57867;
    wire N__57866;
    wire N__57865;
    wire N__57864;
    wire N__57863;
    wire N__57862;
    wire N__57861;
    wire N__57860;
    wire N__57859;
    wire N__57858;
    wire N__57857;
    wire N__57856;
    wire N__57855;
    wire N__57854;
    wire N__57853;
    wire N__57852;
    wire N__57851;
    wire N__57850;
    wire N__57849;
    wire N__57848;
    wire N__57847;
    wire N__57846;
    wire N__57845;
    wire N__57844;
    wire N__57843;
    wire N__57842;
    wire N__57841;
    wire N__57838;
    wire N__57837;
    wire N__57836;
    wire N__57835;
    wire N__57834;
    wire N__57833;
    wire N__57832;
    wire N__57831;
    wire N__57830;
    wire N__57829;
    wire N__57828;
    wire N__57827;
    wire N__57824;
    wire N__57821;
    wire N__57818;
    wire N__57811;
    wire N__57808;
    wire N__57799;
    wire N__57794;
    wire N__57787;
    wire N__57782;
    wire N__57775;
    wire N__57770;
    wire N__57767;
    wire N__57760;
    wire N__57757;
    wire N__57754;
    wire N__57751;
    wire N__57746;
    wire N__57743;
    wire N__57740;
    wire N__57737;
    wire N__57734;
    wire N__57727;
    wire N__57724;
    wire N__57719;
    wire N__57716;
    wire N__57713;
    wire N__57710;
    wire N__57707;
    wire N__57704;
    wire N__57701;
    wire N__57698;
    wire N__57695;
    wire N__57690;
    wire N__57687;
    wire N__57684;
    wire N__57681;
    wire N__57678;
    wire N__57675;
    wire N__57672;
    wire N__57669;
    wire N__57666;
    wire N__57663;
    wire N__57660;
    wire N__57657;
    wire N__57654;
    wire N__57651;
    wire N__57650;
    wire N__57649;
    wire N__57648;
    wire N__57647;
    wire N__57646;
    wire N__57645;
    wire N__57644;
    wire N__57643;
    wire N__57642;
    wire N__57641;
    wire N__57640;
    wire N__57639;
    wire N__57638;
    wire N__57637;
    wire N__57636;
    wire N__57635;
    wire N__57634;
    wire N__57633;
    wire N__57632;
    wire N__57631;
    wire N__57630;
    wire N__57629;
    wire N__57628;
    wire N__57627;
    wire N__57626;
    wire N__57625;
    wire N__57624;
    wire N__57623;
    wire N__57622;
    wire N__57621;
    wire N__57620;
    wire N__57619;
    wire N__57618;
    wire N__57617;
    wire N__57616;
    wire N__57615;
    wire N__57614;
    wire N__57613;
    wire N__57612;
    wire N__57611;
    wire N__57610;
    wire N__57609;
    wire N__57608;
    wire N__57607;
    wire N__57606;
    wire N__57605;
    wire N__57604;
    wire N__57603;
    wire N__57602;
    wire N__57601;
    wire N__57600;
    wire N__57599;
    wire N__57598;
    wire N__57597;
    wire N__57596;
    wire N__57595;
    wire N__57594;
    wire N__57593;
    wire N__57592;
    wire N__57591;
    wire N__57590;
    wire N__57589;
    wire N__57588;
    wire N__57587;
    wire N__57586;
    wire N__57585;
    wire N__57584;
    wire N__57583;
    wire N__57582;
    wire N__57581;
    wire N__57580;
    wire N__57579;
    wire N__57578;
    wire N__57577;
    wire N__57576;
    wire N__57575;
    wire N__57574;
    wire N__57573;
    wire N__57572;
    wire N__57571;
    wire N__57570;
    wire N__57569;
    wire N__57568;
    wire N__57567;
    wire N__57566;
    wire N__57565;
    wire N__57564;
    wire N__57563;
    wire N__57562;
    wire N__57561;
    wire N__57560;
    wire N__57559;
    wire N__57558;
    wire N__57557;
    wire N__57556;
    wire N__57555;
    wire N__57554;
    wire N__57553;
    wire N__57552;
    wire N__57551;
    wire N__57550;
    wire N__57549;
    wire N__57548;
    wire N__57547;
    wire N__57546;
    wire N__57545;
    wire N__57544;
    wire N__57543;
    wire N__57542;
    wire N__57541;
    wire N__57540;
    wire N__57539;
    wire N__57538;
    wire N__57537;
    wire N__57536;
    wire N__57535;
    wire N__57534;
    wire N__57533;
    wire N__57532;
    wire N__57531;
    wire N__57530;
    wire N__57529;
    wire N__57528;
    wire N__57527;
    wire N__57526;
    wire N__57525;
    wire N__57524;
    wire N__57523;
    wire N__57522;
    wire N__57521;
    wire N__57520;
    wire N__57519;
    wire N__57518;
    wire N__57517;
    wire N__57516;
    wire N__57515;
    wire N__57514;
    wire N__57513;
    wire N__57512;
    wire N__57511;
    wire N__57510;
    wire N__57509;
    wire N__57508;
    wire N__57507;
    wire N__57506;
    wire N__57505;
    wire N__57504;
    wire N__57503;
    wire N__57502;
    wire N__57501;
    wire N__57500;
    wire N__57499;
    wire N__57498;
    wire N__57497;
    wire N__57496;
    wire N__57493;
    wire N__57490;
    wire N__57487;
    wire N__57484;
    wire N__57481;
    wire N__57478;
    wire N__57475;
    wire N__57472;
    wire N__57469;
    wire N__57466;
    wire N__57463;
    wire N__57460;
    wire N__57457;
    wire N__57454;
    wire N__57451;
    wire N__57448;
    wire N__57445;
    wire N__57442;
    wire N__57439;
    wire N__57436;
    wire N__57433;
    wire N__57430;
    wire N__57427;
    wire N__57424;
    wire N__57421;
    wire N__57418;
    wire N__57415;
    wire N__57412;
    wire N__57409;
    wire N__57406;
    wire N__57403;
    wire N__57400;
    wire N__57397;
    wire N__57394;
    wire N__57391;
    wire N__57388;
    wire N__57385;
    wire N__57382;
    wire N__57379;
    wire N__57376;
    wire N__57373;
    wire N__57370;
    wire N__57367;
    wire N__57364;
    wire N__57361;
    wire N__57358;
    wire N__56955;
    wire N__56952;
    wire N__56949;
    wire N__56946;
    wire N__56943;
    wire N__56940;
    wire N__56939;
    wire N__56936;
    wire N__56935;
    wire N__56932;
    wire N__56929;
    wire N__56926;
    wire N__56923;
    wire N__56920;
    wire N__56915;
    wire N__56912;
    wire N__56909;
    wire N__56904;
    wire N__56901;
    wire N__56898;
    wire N__56895;
    wire N__56894;
    wire N__56893;
    wire N__56890;
    wire N__56887;
    wire N__56884;
    wire N__56881;
    wire N__56878;
    wire N__56875;
    wire N__56868;
    wire N__56865;
    wire N__56862;
    wire N__56859;
    wire N__56856;
    wire N__56853;
    wire N__56850;
    wire N__56849;
    wire N__56848;
    wire N__56841;
    wire N__56838;
    wire N__56835;
    wire N__56832;
    wire N__56829;
    wire N__56826;
    wire N__56823;
    wire N__56822;
    wire N__56819;
    wire N__56816;
    wire N__56815;
    wire N__56812;
    wire N__56809;
    wire N__56806;
    wire N__56803;
    wire N__56800;
    wire N__56797;
    wire N__56794;
    wire N__56787;
    wire N__56784;
    wire N__56781;
    wire N__56778;
    wire N__56775;
    wire N__56774;
    wire N__56773;
    wire N__56770;
    wire N__56765;
    wire N__56762;
    wire N__56759;
    wire N__56756;
    wire N__56753;
    wire N__56750;
    wire N__56747;
    wire N__56744;
    wire N__56741;
    wire N__56736;
    wire N__56733;
    wire N__56730;
    wire N__56727;
    wire N__56724;
    wire N__56723;
    wire N__56720;
    wire N__56717;
    wire N__56714;
    wire N__56711;
    wire N__56710;
    wire N__56705;
    wire N__56702;
    wire N__56699;
    wire N__56696;
    wire N__56693;
    wire N__56690;
    wire N__56687;
    wire N__56682;
    wire N__56679;
    wire N__56676;
    wire N__56673;
    wire N__56672;
    wire N__56671;
    wire N__56664;
    wire N__56661;
    wire N__56658;
    wire N__56655;
    wire N__56652;
    wire N__56649;
    wire N__56648;
    wire N__56647;
    wire N__56640;
    wire N__56637;
    wire N__56634;
    wire N__56631;
    wire N__56628;
    wire N__56627;
    wire N__56626;
    wire N__56619;
    wire N__56616;
    wire N__56613;
    wire N__56610;
    wire N__56609;
    wire N__56608;
    wire N__56607;
    wire N__56604;
    wire N__56603;
    wire N__56600;
    wire N__56599;
    wire N__56598;
    wire N__56597;
    wire N__56594;
    wire N__56593;
    wire N__56592;
    wire N__56589;
    wire N__56586;
    wire N__56583;
    wire N__56580;
    wire N__56577;
    wire N__56574;
    wire N__56571;
    wire N__56568;
    wire N__56565;
    wire N__56564;
    wire N__56561;
    wire N__56558;
    wire N__56553;
    wire N__56544;
    wire N__56541;
    wire N__56538;
    wire N__56535;
    wire N__56532;
    wire N__56529;
    wire N__56522;
    wire N__56515;
    wire N__56508;
    wire N__56507;
    wire N__56506;
    wire N__56503;
    wire N__56500;
    wire N__56497;
    wire N__56494;
    wire N__56491;
    wire N__56488;
    wire N__56487;
    wire N__56486;
    wire N__56483;
    wire N__56480;
    wire N__56479;
    wire N__56476;
    wire N__56473;
    wire N__56470;
    wire N__56467;
    wire N__56466;
    wire N__56465;
    wire N__56464;
    wire N__56461;
    wire N__56458;
    wire N__56455;
    wire N__56454;
    wire N__56451;
    wire N__56448;
    wire N__56445;
    wire N__56442;
    wire N__56441;
    wire N__56440;
    wire N__56437;
    wire N__56434;
    wire N__56433;
    wire N__56428;
    wire N__56425;
    wire N__56422;
    wire N__56417;
    wire N__56412;
    wire N__56409;
    wire N__56406;
    wire N__56403;
    wire N__56400;
    wire N__56397;
    wire N__56394;
    wire N__56389;
    wire N__56388;
    wire N__56385;
    wire N__56384;
    wire N__56381;
    wire N__56378;
    wire N__56375;
    wire N__56368;
    wire N__56363;
    wire N__56360;
    wire N__56357;
    wire N__56354;
    wire N__56345;
    wire N__56334;
    wire N__56331;
    wire N__56328;
    wire N__56325;
    wire N__56324;
    wire N__56321;
    wire N__56318;
    wire N__56313;
    wire N__56312;
    wire N__56311;
    wire N__56308;
    wire N__56305;
    wire N__56304;
    wire N__56301;
    wire N__56298;
    wire N__56295;
    wire N__56292;
    wire N__56289;
    wire N__56286;
    wire N__56285;
    wire N__56284;
    wire N__56279;
    wire N__56278;
    wire N__56275;
    wire N__56272;
    wire N__56271;
    wire N__56270;
    wire N__56267;
    wire N__56266;
    wire N__56263;
    wire N__56260;
    wire N__56257;
    wire N__56252;
    wire N__56249;
    wire N__56246;
    wire N__56243;
    wire N__56242;
    wire N__56239;
    wire N__56236;
    wire N__56233;
    wire N__56230;
    wire N__56225;
    wire N__56224;
    wire N__56221;
    wire N__56220;
    wire N__56217;
    wire N__56214;
    wire N__56211;
    wire N__56208;
    wire N__56203;
    wire N__56200;
    wire N__56197;
    wire N__56194;
    wire N__56191;
    wire N__56186;
    wire N__56183;
    wire N__56174;
    wire N__56163;
    wire N__56160;
    wire N__56157;
    wire N__56154;
    wire N__56153;
    wire N__56150;
    wire N__56147;
    wire N__56142;
    wire N__56141;
    wire N__56140;
    wire N__56139;
    wire N__56136;
    wire N__56133;
    wire N__56132;
    wire N__56129;
    wire N__56126;
    wire N__56125;
    wire N__56124;
    wire N__56121;
    wire N__56118;
    wire N__56115;
    wire N__56112;
    wire N__56111;
    wire N__56110;
    wire N__56107;
    wire N__56106;
    wire N__56105;
    wire N__56102;
    wire N__56099;
    wire N__56096;
    wire N__56093;
    wire N__56090;
    wire N__56087;
    wire N__56084;
    wire N__56081;
    wire N__56078;
    wire N__56075;
    wire N__56074;
    wire N__56073;
    wire N__56070;
    wire N__56067;
    wire N__56064;
    wire N__56061;
    wire N__56058;
    wire N__56053;
    wire N__56050;
    wire N__56047;
    wire N__56046;
    wire N__56043;
    wire N__56040;
    wire N__56037;
    wire N__56034;
    wire N__56031;
    wire N__56028;
    wire N__56025;
    wire N__56020;
    wire N__56017;
    wire N__56016;
    wire N__56013;
    wire N__56010;
    wire N__56007;
    wire N__56002;
    wire N__56001;
    wire N__55998;
    wire N__55995;
    wire N__55990;
    wire N__55983;
    wire N__55980;
    wire N__55971;
    wire N__55968;
    wire N__55965;
    wire N__55950;
    wire N__55947;
    wire N__55944;
    wire N__55943;
    wire N__55940;
    wire N__55937;
    wire N__55932;
    wire N__55931;
    wire N__55928;
    wire N__55927;
    wire N__55926;
    wire N__55923;
    wire N__55922;
    wire N__55919;
    wire N__55916;
    wire N__55913;
    wire N__55910;
    wire N__55907;
    wire N__55904;
    wire N__55903;
    wire N__55900;
    wire N__55899;
    wire N__55898;
    wire N__55895;
    wire N__55892;
    wire N__55889;
    wire N__55886;
    wire N__55883;
    wire N__55880;
    wire N__55877;
    wire N__55876;
    wire N__55875;
    wire N__55872;
    wire N__55867;
    wire N__55864;
    wire N__55859;
    wire N__55856;
    wire N__55853;
    wire N__55850;
    wire N__55847;
    wire N__55846;
    wire N__55845;
    wire N__55842;
    wire N__55839;
    wire N__55836;
    wire N__55835;
    wire N__55832;
    wire N__55825;
    wire N__55822;
    wire N__55819;
    wire N__55818;
    wire N__55817;
    wire N__55814;
    wire N__55811;
    wire N__55806;
    wire N__55803;
    wire N__55794;
    wire N__55789;
    wire N__55786;
    wire N__55773;
    wire N__55770;
    wire N__55767;
    wire N__55766;
    wire N__55763;
    wire N__55760;
    wire N__55755;
    wire N__55754;
    wire N__55751;
    wire N__55750;
    wire N__55749;
    wire N__55746;
    wire N__55743;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55733;
    wire N__55732;
    wire N__55731;
    wire N__55730;
    wire N__55727;
    wire N__55724;
    wire N__55723;
    wire N__55720;
    wire N__55717;
    wire N__55716;
    wire N__55713;
    wire N__55710;
    wire N__55709;
    wire N__55706;
    wire N__55705;
    wire N__55702;
    wire N__55699;
    wire N__55696;
    wire N__55693;
    wire N__55688;
    wire N__55685;
    wire N__55682;
    wire N__55679;
    wire N__55676;
    wire N__55673;
    wire N__55670;
    wire N__55667;
    wire N__55666;
    wire N__55659;
    wire N__55656;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55644;
    wire N__55639;
    wire N__55636;
    wire N__55633;
    wire N__55630;
    wire N__55625;
    wire N__55616;
    wire N__55605;
    wire N__55602;
    wire N__55599;
    wire N__55596;
    wire N__55595;
    wire N__55592;
    wire N__55589;
    wire N__55584;
    wire N__55583;
    wire N__55582;
    wire N__55581;
    wire N__55578;
    wire N__55575;
    wire N__55574;
    wire N__55571;
    wire N__55568;
    wire N__55567;
    wire N__55566;
    wire N__55565;
    wire N__55562;
    wire N__55559;
    wire N__55556;
    wire N__55553;
    wire N__55550;
    wire N__55549;
    wire N__55548;
    wire N__55545;
    wire N__55542;
    wire N__55541;
    wire N__55538;
    wire N__55535;
    wire N__55534;
    wire N__55531;
    wire N__55528;
    wire N__55525;
    wire N__55522;
    wire N__55521;
    wire N__55518;
    wire N__55515;
    wire N__55512;
    wire N__55509;
    wire N__55506;
    wire N__55503;
    wire N__55500;
    wire N__55497;
    wire N__55494;
    wire N__55489;
    wire N__55486;
    wire N__55483;
    wire N__55480;
    wire N__55477;
    wire N__55474;
    wire N__55471;
    wire N__55468;
    wire N__55465;
    wire N__55462;
    wire N__55459;
    wire N__55456;
    wire N__55453;
    wire N__55450;
    wire N__55447;
    wire N__55446;
    wire N__55445;
    wire N__55436;
    wire N__55431;
    wire N__55428;
    wire N__55421;
    wire N__55416;
    wire N__55413;
    wire N__55410;
    wire N__55395;
    wire N__55392;
    wire N__55389;
    wire N__55388;
    wire N__55385;
    wire N__55382;
    wire N__55377;
    wire N__55374;
    wire N__55373;
    wire N__55372;
    wire N__55369;
    wire N__55366;
    wire N__55363;
    wire N__55362;
    wire N__55357;
    wire N__55356;
    wire N__55355;
    wire N__55354;
    wire N__55353;
    wire N__55350;
    wire N__55347;
    wire N__55344;
    wire N__55343;
    wire N__55342;
    wire N__55339;
    wire N__55336;
    wire N__55333;
    wire N__55332;
    wire N__55329;
    wire N__55326;
    wire N__55323;
    wire N__55320;
    wire N__55317;
    wire N__55314;
    wire N__55311;
    wire N__55308;
    wire N__55305;
    wire N__55302;
    wire N__55299;
    wire N__55296;
    wire N__55293;
    wire N__55290;
    wire N__55285;
    wire N__55284;
    wire N__55281;
    wire N__55280;
    wire N__55273;
    wire N__55270;
    wire N__55265;
    wire N__55260;
    wire N__55257;
    wire N__55254;
    wire N__55251;
    wire N__55248;
    wire N__55239;
    wire N__55230;
    wire N__55227;
    wire N__55224;
    wire N__55223;
    wire N__55220;
    wire N__55217;
    wire N__55212;
    wire N__55209;
    wire N__55206;
    wire N__55205;
    wire N__55202;
    wire N__55199;
    wire N__55194;
    wire N__55191;
    wire N__55188;
    wire N__55185;
    wire N__55182;
    wire N__55179;
    wire N__55176;
    wire N__55173;
    wire N__55170;
    wire N__55169;
    wire N__55168;
    wire N__55165;
    wire N__55162;
    wire N__55159;
    wire N__55154;
    wire N__55151;
    wire N__55148;
    wire N__55145;
    wire N__55140;
    wire N__55137;
    wire N__55134;
    wire N__55133;
    wire N__55132;
    wire N__55125;
    wire N__55122;
    wire N__55119;
    wire N__55116;
    wire N__55113;
    wire N__55110;
    wire N__55107;
    wire N__55104;
    wire N__55103;
    wire N__55102;
    wire N__55095;
    wire N__55092;
    wire N__55089;
    wire N__55086;
    wire N__55083;
    wire N__55080;
    wire N__55079;
    wire N__55078;
    wire N__55075;
    wire N__55070;
    wire N__55067;
    wire N__55064;
    wire N__55061;
    wire N__55058;
    wire N__55053;
    wire N__55050;
    wire N__55047;
    wire N__55044;
    wire N__55043;
    wire N__55042;
    wire N__55035;
    wire N__55032;
    wire N__55029;
    wire N__55026;
    wire N__55023;
    wire N__55020;
    wire N__55017;
    wire N__55014;
    wire N__55011;
    wire N__55010;
    wire N__55009;
    wire N__55006;
    wire N__55001;
    wire N__54996;
    wire N__54993;
    wire N__54990;
    wire N__54987;
    wire N__54984;
    wire N__54983;
    wire N__54982;
    wire N__54975;
    wire N__54972;
    wire N__54969;
    wire N__54966;
    wire N__54963;
    wire N__54960;
    wire N__54959;
    wire N__54958;
    wire N__54957;
    wire N__54954;
    wire N__54947;
    wire N__54942;
    wire N__54939;
    wire N__54936;
    wire N__54933;
    wire N__54930;
    wire N__54929;
    wire N__54928;
    wire N__54927;
    wire N__54924;
    wire N__54917;
    wire N__54912;
    wire N__54911;
    wire N__54910;
    wire N__54909;
    wire N__54906;
    wire N__54899;
    wire N__54894;
    wire N__54891;
    wire N__54888;
    wire N__54885;
    wire N__54882;
    wire N__54879;
    wire N__54876;
    wire N__54873;
    wire N__54870;
    wire N__54869;
    wire N__54868;
    wire N__54865;
    wire N__54860;
    wire N__54857;
    wire N__54854;
    wire N__54851;
    wire N__54846;
    wire N__54843;
    wire N__54840;
    wire N__54837;
    wire N__54836;
    wire N__54835;
    wire N__54832;
    wire N__54827;
    wire N__54822;
    wire N__54819;
    wire N__54816;
    wire N__54813;
    wire N__54812;
    wire N__54809;
    wire N__54808;
    wire N__54805;
    wire N__54802;
    wire N__54799;
    wire N__54792;
    wire N__54789;
    wire N__54786;
    wire N__54783;
    wire N__54780;
    wire N__54777;
    wire N__54776;
    wire N__54775;
    wire N__54768;
    wire N__54765;
    wire N__54762;
    wire N__54759;
    wire N__54756;
    wire N__54753;
    wire N__54752;
    wire N__54751;
    wire N__54748;
    wire N__54743;
    wire N__54740;
    wire N__54737;
    wire N__54734;
    wire N__54731;
    wire N__54728;
    wire N__54725;
    wire N__54720;
    wire N__54717;
    wire N__54714;
    wire N__54711;
    wire N__54710;
    wire N__54709;
    wire N__54702;
    wire N__54699;
    wire N__54696;
    wire N__54693;
    wire N__54690;
    wire N__54687;
    wire N__54684;
    wire N__54681;
    wire N__54680;
    wire N__54675;
    wire N__54672;
    wire N__54669;
    wire N__54666;
    wire N__54663;
    wire N__54660;
    wire N__54657;
    wire N__54656;
    wire N__54653;
    wire N__54650;
    wire N__54649;
    wire N__54642;
    wire N__54639;
    wire N__54636;
    wire N__54633;
    wire N__54630;
    wire N__54629;
    wire N__54626;
    wire N__54623;
    wire N__54620;
    wire N__54615;
    wire N__54612;
    wire N__54609;
    wire N__54606;
    wire N__54603;
    wire N__54600;
    wire N__54597;
    wire N__54594;
    wire N__54591;
    wire N__54588;
    wire N__54585;
    wire N__54582;
    wire N__54579;
    wire N__54576;
    wire N__54573;
    wire N__54570;
    wire N__54569;
    wire N__54568;
    wire N__54567;
    wire N__54564;
    wire N__54557;
    wire N__54552;
    wire N__54549;
    wire N__54546;
    wire N__54543;
    wire N__54540;
    wire N__54537;
    wire N__54536;
    wire N__54535;
    wire N__54532;
    wire N__54527;
    wire N__54522;
    wire N__54519;
    wire N__54516;
    wire N__54513;
    wire N__54512;
    wire N__54507;
    wire N__54504;
    wire N__54501;
    wire N__54498;
    wire N__54495;
    wire N__54494;
    wire N__54493;
    wire N__54490;
    wire N__54489;
    wire N__54482;
    wire N__54479;
    wire N__54476;
    wire N__54471;
    wire N__54468;
    wire N__54465;
    wire N__54462;
    wire N__54459;
    wire N__54458;
    wire N__54455;
    wire N__54452;
    wire N__54447;
    wire N__54444;
    wire N__54441;
    wire N__54438;
    wire N__54435;
    wire N__54432;
    wire N__54431;
    wire N__54428;
    wire N__54425;
    wire N__54422;
    wire N__54419;
    wire N__54416;
    wire N__54411;
    wire N__54408;
    wire N__54405;
    wire N__54402;
    wire N__54401;
    wire N__54398;
    wire N__54395;
    wire N__54392;
    wire N__54389;
    wire N__54384;
    wire N__54381;
    wire N__54378;
    wire N__54377;
    wire N__54374;
    wire N__54371;
    wire N__54366;
    wire N__54363;
    wire N__54360;
    wire N__54357;
    wire N__54354;
    wire N__54351;
    wire N__54348;
    wire N__54347;
    wire N__54346;
    wire N__54343;
    wire N__54340;
    wire N__54337;
    wire N__54334;
    wire N__54327;
    wire N__54324;
    wire N__54321;
    wire N__54318;
    wire N__54315;
    wire N__54314;
    wire N__54309;
    wire N__54308;
    wire N__54305;
    wire N__54302;
    wire N__54297;
    wire N__54294;
    wire N__54291;
    wire N__54288;
    wire N__54285;
    wire N__54282;
    wire N__54279;
    wire N__54278;
    wire N__54273;
    wire N__54270;
    wire N__54267;
    wire N__54264;
    wire N__54261;
    wire N__54258;
    wire N__54257;
    wire N__54252;
    wire N__54249;
    wire N__54246;
    wire N__54243;
    wire N__54240;
    wire N__54239;
    wire N__54234;
    wire N__54231;
    wire N__54228;
    wire N__54225;
    wire N__54222;
    wire N__54219;
    wire N__54218;
    wire N__54213;
    wire N__54210;
    wire N__54207;
    wire N__54204;
    wire N__54201;
    wire N__54198;
    wire N__54197;
    wire N__54192;
    wire N__54189;
    wire N__54186;
    wire N__54183;
    wire N__54180;
    wire N__54179;
    wire N__54174;
    wire N__54171;
    wire N__54168;
    wire N__54165;
    wire N__54162;
    wire N__54159;
    wire N__54156;
    wire N__54153;
    wire N__54152;
    wire N__54147;
    wire N__54144;
    wire N__54141;
    wire N__54140;
    wire N__54139;
    wire N__54136;
    wire N__54133;
    wire N__54130;
    wire N__54123;
    wire N__54122;
    wire N__54121;
    wire N__54118;
    wire N__54113;
    wire N__54110;
    wire N__54107;
    wire N__54102;
    wire N__54099;
    wire N__54096;
    wire N__54095;
    wire N__54094;
    wire N__54091;
    wire N__54086;
    wire N__54081;
    wire N__54078;
    wire N__54077;
    wire N__54072;
    wire N__54069;
    wire N__54066;
    wire N__54063;
    wire N__54060;
    wire N__54057;
    wire N__54054;
    wire N__54053;
    wire N__54052;
    wire N__54049;
    wire N__54044;
    wire N__54039;
    wire N__54036;
    wire N__54035;
    wire N__54034;
    wire N__54031;
    wire N__54030;
    wire N__54029;
    wire N__54028;
    wire N__54025;
    wire N__54022;
    wire N__54015;
    wire N__54010;
    wire N__54007;
    wire N__54002;
    wire N__53999;
    wire N__53996;
    wire N__53991;
    wire N__53990;
    wire N__53987;
    wire N__53984;
    wire N__53983;
    wire N__53982;
    wire N__53981;
    wire N__53980;
    wire N__53979;
    wire N__53978;
    wire N__53975;
    wire N__53974;
    wire N__53971;
    wire N__53962;
    wire N__53957;
    wire N__53954;
    wire N__53951;
    wire N__53948;
    wire N__53939;
    wire N__53936;
    wire N__53933;
    wire N__53928;
    wire N__53925;
    wire N__53922;
    wire N__53919;
    wire N__53916;
    wire N__53915;
    wire N__53912;
    wire N__53911;
    wire N__53908;
    wire N__53905;
    wire N__53902;
    wire N__53899;
    wire N__53894;
    wire N__53891;
    wire N__53888;
    wire N__53885;
    wire N__53882;
    wire N__53879;
    wire N__53876;
    wire N__53873;
    wire N__53870;
    wire N__53865;
    wire N__53862;
    wire N__53859;
    wire N__53856;
    wire N__53853;
    wire N__53850;
    wire N__53849;
    wire N__53848;
    wire N__53845;
    wire N__53840;
    wire N__53835;
    wire N__53832;
    wire N__53829;
    wire N__53826;
    wire N__53823;
    wire N__53820;
    wire N__53819;
    wire N__53816;
    wire N__53815;
    wire N__53814;
    wire N__53811;
    wire N__53808;
    wire N__53803;
    wire N__53796;
    wire N__53795;
    wire N__53792;
    wire N__53789;
    wire N__53788;
    wire N__53785;
    wire N__53784;
    wire N__53779;
    wire N__53776;
    wire N__53773;
    wire N__53770;
    wire N__53763;
    wire N__53760;
    wire N__53757;
    wire N__53756;
    wire N__53753;
    wire N__53750;
    wire N__53747;
    wire N__53744;
    wire N__53741;
    wire N__53738;
    wire N__53735;
    wire N__53730;
    wire N__53727;
    wire N__53724;
    wire N__53721;
    wire N__53718;
    wire N__53715;
    wire N__53712;
    wire N__53709;
    wire N__53706;
    wire N__53703;
    wire N__53700;
    wire N__53697;
    wire N__53694;
    wire N__53691;
    wire N__53690;
    wire N__53689;
    wire N__53688;
    wire N__53685;
    wire N__53678;
    wire N__53673;
    wire N__53672;
    wire N__53669;
    wire N__53666;
    wire N__53663;
    wire N__53658;
    wire N__53655;
    wire N__53652;
    wire N__53649;
    wire N__53646;
    wire N__53645;
    wire N__53644;
    wire N__53639;
    wire N__53636;
    wire N__53633;
    wire N__53628;
    wire N__53625;
    wire N__53624;
    wire N__53623;
    wire N__53620;
    wire N__53615;
    wire N__53610;
    wire N__53609;
    wire N__53604;
    wire N__53601;
    wire N__53600;
    wire N__53599;
    wire N__53596;
    wire N__53591;
    wire N__53586;
    wire N__53583;
    wire N__53582;
    wire N__53577;
    wire N__53574;
    wire N__53573;
    wire N__53570;
    wire N__53567;
    wire N__53564;
    wire N__53561;
    wire N__53556;
    wire N__53553;
    wire N__53550;
    wire N__53547;
    wire N__53544;
    wire N__53541;
    wire N__53538;
    wire N__53537;
    wire N__53534;
    wire N__53531;
    wire N__53528;
    wire N__53523;
    wire N__53520;
    wire N__53517;
    wire N__53514;
    wire N__53511;
    wire N__53510;
    wire N__53509;
    wire N__53506;
    wire N__53503;
    wire N__53500;
    wire N__53497;
    wire N__53494;
    wire N__53491;
    wire N__53486;
    wire N__53483;
    wire N__53480;
    wire N__53475;
    wire N__53472;
    wire N__53469;
    wire N__53466;
    wire N__53463;
    wire N__53460;
    wire N__53459;
    wire N__53458;
    wire N__53451;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53439;
    wire N__53436;
    wire N__53435;
    wire N__53432;
    wire N__53431;
    wire N__53428;
    wire N__53425;
    wire N__53420;
    wire N__53415;
    wire N__53412;
    wire N__53409;
    wire N__53406;
    wire N__53405;
    wire N__53402;
    wire N__53401;
    wire N__53398;
    wire N__53397;
    wire N__53396;
    wire N__53393;
    wire N__53390;
    wire N__53387;
    wire N__53386;
    wire N__53383;
    wire N__53380;
    wire N__53379;
    wire N__53376;
    wire N__53371;
    wire N__53370;
    wire N__53367;
    wire N__53364;
    wire N__53361;
    wire N__53360;
    wire N__53357;
    wire N__53354;
    wire N__53351;
    wire N__53350;
    wire N__53349;
    wire N__53346;
    wire N__53343;
    wire N__53340;
    wire N__53337;
    wire N__53334;
    wire N__53331;
    wire N__53326;
    wire N__53325;
    wire N__53324;
    wire N__53321;
    wire N__53318;
    wire N__53315;
    wire N__53312;
    wire N__53309;
    wire N__53306;
    wire N__53303;
    wire N__53300;
    wire N__53297;
    wire N__53294;
    wire N__53291;
    wire N__53288;
    wire N__53283;
    wire N__53280;
    wire N__53275;
    wire N__53266;
    wire N__53253;
    wire N__53250;
    wire N__53249;
    wire N__53246;
    wire N__53243;
    wire N__53240;
    wire N__53237;
    wire N__53232;
    wire N__53229;
    wire N__53228;
    wire N__53225;
    wire N__53224;
    wire N__53221;
    wire N__53218;
    wire N__53215;
    wire N__53212;
    wire N__53211;
    wire N__53206;
    wire N__53205;
    wire N__53204;
    wire N__53201;
    wire N__53198;
    wire N__53195;
    wire N__53192;
    wire N__53189;
    wire N__53186;
    wire N__53185;
    wire N__53184;
    wire N__53181;
    wire N__53178;
    wire N__53173;
    wire N__53170;
    wire N__53167;
    wire N__53164;
    wire N__53161;
    wire N__53156;
    wire N__53149;
    wire N__53142;
    wire N__53141;
    wire N__53136;
    wire N__53133;
    wire N__53130;
    wire N__53129;
    wire N__53126;
    wire N__53123;
    wire N__53118;
    wire N__53117;
    wire N__53114;
    wire N__53111;
    wire N__53108;
    wire N__53105;
    wire N__53102;
    wire N__53099;
    wire N__53094;
    wire N__53091;
    wire N__53088;
    wire N__53085;
    wire N__53082;
    wire N__53081;
    wire N__53080;
    wire N__53073;
    wire N__53070;
    wire N__53067;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53054;
    wire N__53051;
    wire N__53048;
    wire N__53043;
    wire N__53040;
    wire N__53037;
    wire N__53034;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53022;
    wire N__53021;
    wire N__53020;
    wire N__53013;
    wire N__53010;
    wire N__53007;
    wire N__53004;
    wire N__53001;
    wire N__52998;
    wire N__52997;
    wire N__52992;
    wire N__52989;
    wire N__52986;
    wire N__52985;
    wire N__52982;
    wire N__52979;
    wire N__52974;
    wire N__52971;
    wire N__52970;
    wire N__52969;
    wire N__52966;
    wire N__52961;
    wire N__52956;
    wire N__52955;
    wire N__52954;
    wire N__52947;
    wire N__52944;
    wire N__52941;
    wire N__52938;
    wire N__52935;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52923;
    wire N__52920;
    wire N__52917;
    wire N__52914;
    wire N__52911;
    wire N__52908;
    wire N__52905;
    wire N__52904;
    wire N__52899;
    wire N__52896;
    wire N__52893;
    wire N__52890;
    wire N__52889;
    wire N__52886;
    wire N__52883;
    wire N__52878;
    wire N__52877;
    wire N__52874;
    wire N__52871;
    wire N__52868;
    wire N__52865;
    wire N__52860;
    wire N__52857;
    wire N__52854;
    wire N__52851;
    wire N__52848;
    wire N__52845;
    wire N__52844;
    wire N__52839;
    wire N__52836;
    wire N__52833;
    wire N__52830;
    wire N__52827;
    wire N__52824;
    wire N__52821;
    wire N__52820;
    wire N__52815;
    wire N__52812;
    wire N__52811;
    wire N__52806;
    wire N__52803;
    wire N__52800;
    wire N__52797;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52779;
    wire N__52776;
    wire N__52773;
    wire N__52770;
    wire N__52769;
    wire N__52766;
    wire N__52763;
    wire N__52760;
    wire N__52757;
    wire N__52754;
    wire N__52751;
    wire N__52746;
    wire N__52743;
    wire N__52740;
    wire N__52737;
    wire N__52736;
    wire N__52733;
    wire N__52730;
    wire N__52727;
    wire N__52724;
    wire N__52721;
    wire N__52718;
    wire N__52713;
    wire N__52710;
    wire N__52709;
    wire N__52708;
    wire N__52705;
    wire N__52702;
    wire N__52699;
    wire N__52694;
    wire N__52693;
    wire N__52690;
    wire N__52687;
    wire N__52684;
    wire N__52683;
    wire N__52680;
    wire N__52679;
    wire N__52676;
    wire N__52673;
    wire N__52670;
    wire N__52667;
    wire N__52664;
    wire N__52663;
    wire N__52656;
    wire N__52653;
    wire N__52650;
    wire N__52649;
    wire N__52646;
    wire N__52643;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52626;
    wire N__52621;
    wire N__52614;
    wire N__52613;
    wire N__52608;
    wire N__52605;
    wire N__52602;
    wire N__52599;
    wire N__52598;
    wire N__52597;
    wire N__52594;
    wire N__52591;
    wire N__52590;
    wire N__52587;
    wire N__52586;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52576;
    wire N__52573;
    wire N__52570;
    wire N__52565;
    wire N__52562;
    wire N__52559;
    wire N__52556;
    wire N__52553;
    wire N__52546;
    wire N__52543;
    wire N__52542;
    wire N__52541;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52529;
    wire N__52526;
    wire N__52523;
    wire N__52520;
    wire N__52513;
    wire N__52506;
    wire N__52503;
    wire N__52502;
    wire N__52501;
    wire N__52498;
    wire N__52493;
    wire N__52488;
    wire N__52485;
    wire N__52484;
    wire N__52481;
    wire N__52478;
    wire N__52477;
    wire N__52472;
    wire N__52469;
    wire N__52468;
    wire N__52467;
    wire N__52464;
    wire N__52461;
    wire N__52458;
    wire N__52457;
    wire N__52454;
    wire N__52449;
    wire N__52446;
    wire N__52443;
    wire N__52440;
    wire N__52433;
    wire N__52430;
    wire N__52427;
    wire N__52426;
    wire N__52423;
    wire N__52420;
    wire N__52417;
    wire N__52410;
    wire N__52407;
    wire N__52406;
    wire N__52403;
    wire N__52400;
    wire N__52395;
    wire N__52392;
    wire N__52391;
    wire N__52388;
    wire N__52385;
    wire N__52384;
    wire N__52379;
    wire N__52378;
    wire N__52375;
    wire N__52374;
    wire N__52371;
    wire N__52368;
    wire N__52365;
    wire N__52362;
    wire N__52361;
    wire N__52356;
    wire N__52351;
    wire N__52348;
    wire N__52347;
    wire N__52344;
    wire N__52341;
    wire N__52338;
    wire N__52335;
    wire N__52332;
    wire N__52327;
    wire N__52324;
    wire N__52317;
    wire N__52314;
    wire N__52311;
    wire N__52308;
    wire N__52307;
    wire N__52304;
    wire N__52301;
    wire N__52300;
    wire N__52295;
    wire N__52292;
    wire N__52291;
    wire N__52288;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52274;
    wire N__52273;
    wire N__52268;
    wire N__52265;
    wire N__52260;
    wire N__52259;
    wire N__52256;
    wire N__52253;
    wire N__52248;
    wire N__52247;
    wire N__52244;
    wire N__52241;
    wire N__52236;
    wire N__52233;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52221;
    wire N__52218;
    wire N__52217;
    wire N__52216;
    wire N__52213;
    wire N__52208;
    wire N__52203;
    wire N__52200;
    wire N__52197;
    wire N__52194;
    wire N__52191;
    wire N__52188;
    wire N__52185;
    wire N__52182;
    wire N__52179;
    wire N__52176;
    wire N__52173;
    wire N__52170;
    wire N__52167;
    wire N__52166;
    wire N__52163;
    wire N__52160;
    wire N__52157;
    wire N__52154;
    wire N__52149;
    wire N__52146;
    wire N__52143;
    wire N__52140;
    wire N__52137;
    wire N__52134;
    wire N__52131;
    wire N__52128;
    wire N__52127;
    wire N__52124;
    wire N__52121;
    wire N__52118;
    wire N__52115;
    wire N__52110;
    wire N__52107;
    wire N__52104;
    wire N__52101;
    wire N__52098;
    wire N__52095;
    wire N__52092;
    wire N__52089;
    wire N__52086;
    wire N__52083;
    wire N__52082;
    wire N__52079;
    wire N__52076;
    wire N__52071;
    wire N__52068;
    wire N__52065;
    wire N__52062;
    wire N__52059;
    wire N__52056;
    wire N__52053;
    wire N__52050;
    wire N__52047;
    wire N__52044;
    wire N__52041;
    wire N__52038;
    wire N__52035;
    wire N__52032;
    wire N__52029;
    wire N__52028;
    wire N__52025;
    wire N__52022;
    wire N__52017;
    wire N__52014;
    wire N__52011;
    wire N__52008;
    wire N__52005;
    wire N__52002;
    wire N__51999;
    wire N__51996;
    wire N__51993;
    wire N__51990;
    wire N__51987;
    wire N__51984;
    wire N__51981;
    wire N__51978;
    wire N__51977;
    wire N__51974;
    wire N__51971;
    wire N__51968;
    wire N__51965;
    wire N__51962;
    wire N__51959;
    wire N__51954;
    wire N__51951;
    wire N__51948;
    wire N__51945;
    wire N__51942;
    wire N__51941;
    wire N__51938;
    wire N__51935;
    wire N__51932;
    wire N__51929;
    wire N__51926;
    wire N__51923;
    wire N__51918;
    wire N__51915;
    wire N__51912;
    wire N__51909;
    wire N__51906;
    wire N__51905;
    wire N__51902;
    wire N__51899;
    wire N__51896;
    wire N__51893;
    wire N__51890;
    wire N__51887;
    wire N__51882;
    wire N__51879;
    wire N__51876;
    wire N__51873;
    wire N__51870;
    wire N__51869;
    wire N__51866;
    wire N__51863;
    wire N__51860;
    wire N__51857;
    wire N__51854;
    wire N__51851;
    wire N__51846;
    wire N__51843;
    wire N__51842;
    wire N__51837;
    wire N__51834;
    wire N__51833;
    wire N__51830;
    wire N__51827;
    wire N__51826;
    wire N__51823;
    wire N__51820;
    wire N__51817;
    wire N__51810;
    wire N__51809;
    wire N__51806;
    wire N__51803;
    wire N__51800;
    wire N__51797;
    wire N__51794;
    wire N__51789;
    wire N__51786;
    wire N__51783;
    wire N__51780;
    wire N__51779;
    wire N__51776;
    wire N__51773;
    wire N__51772;
    wire N__51769;
    wire N__51766;
    wire N__51763;
    wire N__51756;
    wire N__51753;
    wire N__51750;
    wire N__51747;
    wire N__51744;
    wire N__51741;
    wire N__51740;
    wire N__51737;
    wire N__51734;
    wire N__51731;
    wire N__51728;
    wire N__51725;
    wire N__51722;
    wire N__51717;
    wire N__51714;
    wire N__51711;
    wire N__51708;
    wire N__51705;
    wire N__51704;
    wire N__51701;
    wire N__51698;
    wire N__51695;
    wire N__51692;
    wire N__51689;
    wire N__51686;
    wire N__51681;
    wire N__51678;
    wire N__51675;
    wire N__51672;
    wire N__51669;
    wire N__51666;
    wire N__51665;
    wire N__51662;
    wire N__51659;
    wire N__51654;
    wire N__51651;
    wire N__51648;
    wire N__51645;
    wire N__51642;
    wire N__51639;
    wire N__51636;
    wire N__51633;
    wire N__51630;
    wire N__51627;
    wire N__51624;
    wire N__51621;
    wire N__51620;
    wire N__51617;
    wire N__51614;
    wire N__51611;
    wire N__51608;
    wire N__51603;
    wire N__51600;
    wire N__51597;
    wire N__51594;
    wire N__51591;
    wire N__51588;
    wire N__51585;
    wire N__51582;
    wire N__51579;
    wire N__51576;
    wire N__51575;
    wire N__51572;
    wire N__51569;
    wire N__51566;
    wire N__51563;
    wire N__51558;
    wire N__51555;
    wire N__51552;
    wire N__51549;
    wire N__51548;
    wire N__51545;
    wire N__51542;
    wire N__51537;
    wire N__51536;
    wire N__51535;
    wire N__51528;
    wire N__51525;
    wire N__51524;
    wire N__51523;
    wire N__51520;
    wire N__51515;
    wire N__51510;
    wire N__51507;
    wire N__51506;
    wire N__51503;
    wire N__51500;
    wire N__51495;
    wire N__51492;
    wire N__51489;
    wire N__51486;
    wire N__51483;
    wire N__51482;
    wire N__51479;
    wire N__51476;
    wire N__51473;
    wire N__51468;
    wire N__51465;
    wire N__51462;
    wire N__51459;
    wire N__51456;
    wire N__51453;
    wire N__51452;
    wire N__51451;
    wire N__51450;
    wire N__51449;
    wire N__51448;
    wire N__51445;
    wire N__51442;
    wire N__51437;
    wire N__51436;
    wire N__51433;
    wire N__51432;
    wire N__51431;
    wire N__51428;
    wire N__51427;
    wire N__51426;
    wire N__51419;
    wire N__51416;
    wire N__51415;
    wire N__51412;
    wire N__51411;
    wire N__51410;
    wire N__51409;
    wire N__51406;
    wire N__51405;
    wire N__51404;
    wire N__51401;
    wire N__51400;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51386;
    wire N__51383;
    wire N__51382;
    wire N__51381;
    wire N__51378;
    wire N__51375;
    wire N__51372;
    wire N__51369;
    wire N__51366;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51356;
    wire N__51353;
    wire N__51350;
    wire N__51347;
    wire N__51342;
    wire N__51339;
    wire N__51334;
    wire N__51329;
    wire N__51324;
    wire N__51321;
    wire N__51318;
    wire N__51315;
    wire N__51310;
    wire N__51307;
    wire N__51298;
    wire N__51291;
    wire N__51282;
    wire N__51273;
    wire N__51270;
    wire N__51269;
    wire N__51266;
    wire N__51265;
    wire N__51262;
    wire N__51259;
    wire N__51256;
    wire N__51249;
    wire N__51246;
    wire N__51243;
    wire N__51240;
    wire N__51237;
    wire N__51234;
    wire N__51231;
    wire N__51228;
    wire N__51227;
    wire N__51226;
    wire N__51223;
    wire N__51220;
    wire N__51215;
    wire N__51210;
    wire N__51207;
    wire N__51204;
    wire N__51201;
    wire N__51198;
    wire N__51195;
    wire N__51192;
    wire N__51189;
    wire N__51186;
    wire N__51183;
    wire N__51180;
    wire N__51179;
    wire N__51176;
    wire N__51173;
    wire N__51170;
    wire N__51165;
    wire N__51162;
    wire N__51159;
    wire N__51158;
    wire N__51155;
    wire N__51152;
    wire N__51147;
    wire N__51144;
    wire N__51143;
    wire N__51138;
    wire N__51135;
    wire N__51132;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51122;
    wire N__51119;
    wire N__51116;
    wire N__51113;
    wire N__51110;
    wire N__51105;
    wire N__51102;
    wire N__51099;
    wire N__51096;
    wire N__51093;
    wire N__51090;
    wire N__51087;
    wire N__51084;
    wire N__51081;
    wire N__51078;
    wire N__51075;
    wire N__51072;
    wire N__51069;
    wire N__51066;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51047;
    wire N__51046;
    wire N__51043;
    wire N__51038;
    wire N__51033;
    wire N__51030;
    wire N__51027;
    wire N__51026;
    wire N__51023;
    wire N__51020;
    wire N__51015;
    wire N__51012;
    wire N__51011;
    wire N__51006;
    wire N__51003;
    wire N__51000;
    wire N__50997;
    wire N__50994;
    wire N__50993;
    wire N__50992;
    wire N__50989;
    wire N__50984;
    wire N__50979;
    wire N__50978;
    wire N__50973;
    wire N__50970;
    wire N__50967;
    wire N__50966;
    wire N__50963;
    wire N__50960;
    wire N__50957;
    wire N__50952;
    wire N__50951;
    wire N__50950;
    wire N__50943;
    wire N__50940;
    wire N__50937;
    wire N__50936;
    wire N__50933;
    wire N__50930;
    wire N__50925;
    wire N__50922;
    wire N__50919;
    wire N__50916;
    wire N__50913;
    wire N__50910;
    wire N__50907;
    wire N__50904;
    wire N__50901;
    wire N__50900;
    wire N__50895;
    wire N__50892;
    wire N__50889;
    wire N__50888;
    wire N__50883;
    wire N__50880;
    wire N__50877;
    wire N__50874;
    wire N__50871;
    wire N__50868;
    wire N__50867;
    wire N__50866;
    wire N__50859;
    wire N__50856;
    wire N__50853;
    wire N__50850;
    wire N__50847;
    wire N__50844;
    wire N__50841;
    wire N__50838;
    wire N__50835;
    wire N__50832;
    wire N__50829;
    wire N__50828;
    wire N__50825;
    wire N__50822;
    wire N__50817;
    wire N__50814;
    wire N__50811;
    wire N__50808;
    wire N__50807;
    wire N__50802;
    wire N__50799;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50781;
    wire N__50780;
    wire N__50779;
    wire N__50776;
    wire N__50773;
    wire N__50772;
    wire N__50769;
    wire N__50768;
    wire N__50767;
    wire N__50762;
    wire N__50759;
    wire N__50756;
    wire N__50753;
    wire N__50750;
    wire N__50749;
    wire N__50746;
    wire N__50743;
    wire N__50738;
    wire N__50735;
    wire N__50732;
    wire N__50731;
    wire N__50728;
    wire N__50725;
    wire N__50718;
    wire N__50715;
    wire N__50706;
    wire N__50703;
    wire N__50700;
    wire N__50697;
    wire N__50696;
    wire N__50693;
    wire N__50692;
    wire N__50689;
    wire N__50686;
    wire N__50683;
    wire N__50680;
    wire N__50677;
    wire N__50674;
    wire N__50671;
    wire N__50668;
    wire N__50665;
    wire N__50662;
    wire N__50659;
    wire N__50656;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50631;
    wire N__50628;
    wire N__50625;
    wire N__50624;
    wire N__50623;
    wire N__50622;
    wire N__50619;
    wire N__50612;
    wire N__50611;
    wire N__50610;
    wire N__50609;
    wire N__50608;
    wire N__50607;
    wire N__50606;
    wire N__50605;
    wire N__50602;
    wire N__50599;
    wire N__50596;
    wire N__50583;
    wire N__50580;
    wire N__50577;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50556;
    wire N__50553;
    wire N__50544;
    wire N__50541;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50529;
    wire N__50526;
    wire N__50523;
    wire N__50520;
    wire N__50519;
    wire N__50516;
    wire N__50513;
    wire N__50508;
    wire N__50507;
    wire N__50506;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50494;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50484;
    wire N__50481;
    wire N__50480;
    wire N__50477;
    wire N__50474;
    wire N__50471;
    wire N__50468;
    wire N__50465;
    wire N__50462;
    wire N__50459;
    wire N__50454;
    wire N__50447;
    wire N__50442;
    wire N__50441;
    wire N__50438;
    wire N__50435;
    wire N__50434;
    wire N__50431;
    wire N__50428;
    wire N__50425;
    wire N__50420;
    wire N__50417;
    wire N__50414;
    wire N__50409;
    wire N__50406;
    wire N__50403;
    wire N__50402;
    wire N__50399;
    wire N__50398;
    wire N__50395;
    wire N__50394;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50380;
    wire N__50375;
    wire N__50372;
    wire N__50369;
    wire N__50366;
    wire N__50363;
    wire N__50360;
    wire N__50357;
    wire N__50354;
    wire N__50351;
    wire N__50348;
    wire N__50345;
    wire N__50340;
    wire N__50337;
    wire N__50336;
    wire N__50333;
    wire N__50330;
    wire N__50327;
    wire N__50324;
    wire N__50321;
    wire N__50310;
    wire N__50307;
    wire N__50304;
    wire N__50301;
    wire N__50298;
    wire N__50297;
    wire N__50294;
    wire N__50291;
    wire N__50288;
    wire N__50285;
    wire N__50280;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50268;
    wire N__50265;
    wire N__50262;
    wire N__50259;
    wire N__50256;
    wire N__50253;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50241;
    wire N__50240;
    wire N__50237;
    wire N__50234;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50219;
    wire N__50214;
    wire N__50211;
    wire N__50208;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50196;
    wire N__50193;
    wire N__50190;
    wire N__50187;
    wire N__50184;
    wire N__50181;
    wire N__50178;
    wire N__50175;
    wire N__50172;
    wire N__50169;
    wire N__50166;
    wire N__50163;
    wire N__50160;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50148;
    wire N__50145;
    wire N__50144;
    wire N__50139;
    wire N__50136;
    wire N__50135;
    wire N__50134;
    wire N__50131;
    wire N__50126;
    wire N__50121;
    wire N__50118;
    wire N__50117;
    wire N__50114;
    wire N__50111;
    wire N__50106;
    wire N__50103;
    wire N__50100;
    wire N__50097;
    wire N__50094;
    wire N__50091;
    wire N__50088;
    wire N__50085;
    wire N__50082;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50070;
    wire N__50067;
    wire N__50064;
    wire N__50061;
    wire N__50058;
    wire N__50055;
    wire N__50052;
    wire N__50049;
    wire N__50046;
    wire N__50043;
    wire N__50040;
    wire N__50037;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50024;
    wire N__50021;
    wire N__50020;
    wire N__50017;
    wire N__50016;
    wire N__50015;
    wire N__50014;
    wire N__50011;
    wire N__50008;
    wire N__50005;
    wire N__49998;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49980;
    wire N__49977;
    wire N__49974;
    wire N__49971;
    wire N__49968;
    wire N__49967;
    wire N__49966;
    wire N__49965;
    wire N__49962;
    wire N__49959;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49947;
    wire N__49942;
    wire N__49939;
    wire N__49932;
    wire N__49929;
    wire N__49928;
    wire N__49927;
    wire N__49926;
    wire N__49923;
    wire N__49920;
    wire N__49917;
    wire N__49914;
    wire N__49911;
    wire N__49904;
    wire N__49901;
    wire N__49896;
    wire N__49893;
    wire N__49892;
    wire N__49889;
    wire N__49886;
    wire N__49883;
    wire N__49882;
    wire N__49881;
    wire N__49876;
    wire N__49871;
    wire N__49868;
    wire N__49865;
    wire N__49860;
    wire N__49857;
    wire N__49856;
    wire N__49855;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49843;
    wire N__49842;
    wire N__49835;
    wire N__49832;
    wire N__49827;
    wire N__49824;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49800;
    wire N__49797;
    wire N__49794;
    wire N__49791;
    wire N__49788;
    wire N__49785;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49761;
    wire N__49758;
    wire N__49755;
    wire N__49752;
    wire N__49749;
    wire N__49748;
    wire N__49745;
    wire N__49742;
    wire N__49739;
    wire N__49736;
    wire N__49731;
    wire N__49728;
    wire N__49725;
    wire N__49724;
    wire N__49721;
    wire N__49718;
    wire N__49715;
    wire N__49712;
    wire N__49709;
    wire N__49706;
    wire N__49701;
    wire N__49698;
    wire N__49697;
    wire N__49696;
    wire N__49695;
    wire N__49694;
    wire N__49691;
    wire N__49688;
    wire N__49685;
    wire N__49682;
    wire N__49681;
    wire N__49678;
    wire N__49675;
    wire N__49672;
    wire N__49665;
    wire N__49664;
    wire N__49661;
    wire N__49656;
    wire N__49653;
    wire N__49650;
    wire N__49647;
    wire N__49642;
    wire N__49639;
    wire N__49636;
    wire N__49633;
    wire N__49628;
    wire N__49623;
    wire N__49620;
    wire N__49619;
    wire N__49618;
    wire N__49615;
    wire N__49612;
    wire N__49611;
    wire N__49608;
    wire N__49605;
    wire N__49602;
    wire N__49599;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49585;
    wire N__49580;
    wire N__49577;
    wire N__49572;
    wire N__49569;
    wire N__49568;
    wire N__49565;
    wire N__49564;
    wire N__49561;
    wire N__49556;
    wire N__49551;
    wire N__49548;
    wire N__49545;
    wire N__49542;
    wire N__49541;
    wire N__49538;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49528;
    wire N__49525;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49509;
    wire N__49508;
    wire N__49507;
    wire N__49504;
    wire N__49499;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49460;
    wire N__49457;
    wire N__49454;
    wire N__49451;
    wire N__49448;
    wire N__49445;
    wire N__49442;
    wire N__49439;
    wire N__49436;
    wire N__49431;
    wire N__49428;
    wire N__49427;
    wire N__49424;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49411;
    wire N__49404;
    wire N__49401;
    wire N__49400;
    wire N__49397;
    wire N__49394;
    wire N__49389;
    wire N__49386;
    wire N__49383;
    wire N__49380;
    wire N__49377;
    wire N__49376;
    wire N__49375;
    wire N__49374;
    wire N__49373;
    wire N__49372;
    wire N__49371;
    wire N__49370;
    wire N__49369;
    wire N__49368;
    wire N__49367;
    wire N__49366;
    wire N__49365;
    wire N__49364;
    wire N__49363;
    wire N__49362;
    wire N__49361;
    wire N__49360;
    wire N__49359;
    wire N__49358;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49308;
    wire N__49305;
    wire N__49302;
    wire N__49301;
    wire N__49296;
    wire N__49295;
    wire N__49292;
    wire N__49289;
    wire N__49286;
    wire N__49283;
    wire N__49280;
    wire N__49277;
    wire N__49272;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49251;
    wire N__49248;
    wire N__49245;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49230;
    wire N__49227;
    wire N__49224;
    wire N__49221;
    wire N__49218;
    wire N__49215;
    wire N__49212;
    wire N__49209;
    wire N__49206;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49191;
    wire N__49188;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49143;
    wire N__49140;
    wire N__49137;
    wire N__49134;
    wire N__49131;
    wire N__49128;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49112;
    wire N__49109;
    wire N__49106;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49091;
    wire N__49088;
    wire N__49083;
    wire N__49082;
    wire N__49081;
    wire N__49080;
    wire N__49079;
    wire N__49078;
    wire N__49077;
    wire N__49076;
    wire N__49075;
    wire N__49074;
    wire N__49073;
    wire N__49070;
    wire N__49069;
    wire N__49068;
    wire N__49067;
    wire N__49066;
    wire N__49065;
    wire N__49062;
    wire N__49061;
    wire N__49060;
    wire N__49053;
    wire N__49044;
    wire N__49043;
    wire N__49040;
    wire N__49037;
    wire N__49034;
    wire N__49027;
    wire N__49026;
    wire N__49025;
    wire N__49024;
    wire N__49023;
    wire N__49022;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49014;
    wire N__49013;
    wire N__49008;
    wire N__49005;
    wire N__49000;
    wire N__48999;
    wire N__48998;
    wire N__48997;
    wire N__48996;
    wire N__48995;
    wire N__48994;
    wire N__48991;
    wire N__48990;
    wire N__48989;
    wire N__48988;
    wire N__48987;
    wire N__48986;
    wire N__48977;
    wire N__48972;
    wire N__48967;
    wire N__48956;
    wire N__48953;
    wire N__48950;
    wire N__48945;
    wire N__48936;
    wire N__48935;
    wire N__48932;
    wire N__48931;
    wire N__48928;
    wire N__48923;
    wire N__48914;
    wire N__48909;
    wire N__48904;
    wire N__48895;
    wire N__48888;
    wire N__48873;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48869;
    wire N__48868;
    wire N__48867;
    wire N__48866;
    wire N__48865;
    wire N__48864;
    wire N__48863;
    wire N__48862;
    wire N__48861;
    wire N__48858;
    wire N__48855;
    wire N__48854;
    wire N__48853;
    wire N__48852;
    wire N__48851;
    wire N__48848;
    wire N__48841;
    wire N__48838;
    wire N__48835;
    wire N__48834;
    wire N__48833;
    wire N__48832;
    wire N__48829;
    wire N__48826;
    wire N__48825;
    wire N__48824;
    wire N__48823;
    wire N__48822;
    wire N__48821;
    wire N__48820;
    wire N__48819;
    wire N__48816;
    wire N__48815;
    wire N__48812;
    wire N__48809;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48799;
    wire N__48798;
    wire N__48797;
    wire N__48796;
    wire N__48795;
    wire N__48794;
    wire N__48793;
    wire N__48792;
    wire N__48791;
    wire N__48790;
    wire N__48789;
    wire N__48786;
    wire N__48781;
    wire N__48776;
    wire N__48769;
    wire N__48764;
    wire N__48759;
    wire N__48744;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48740;
    wire N__48739;
    wire N__48738;
    wire N__48737;
    wire N__48736;
    wire N__48735;
    wire N__48730;
    wire N__48723;
    wire N__48718;
    wire N__48715;
    wire N__48710;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48702;
    wire N__48701;
    wire N__48700;
    wire N__48699;
    wire N__48698;
    wire N__48697;
    wire N__48696;
    wire N__48687;
    wire N__48682;
    wire N__48671;
    wire N__48666;
    wire N__48663;
    wire N__48654;
    wire N__48647;
    wire N__48646;
    wire N__48645;
    wire N__48644;
    wire N__48643;
    wire N__48642;
    wire N__48641;
    wire N__48640;
    wire N__48639;
    wire N__48638;
    wire N__48637;
    wire N__48636;
    wire N__48635;
    wire N__48632;
    wire N__48627;
    wire N__48622;
    wire N__48619;
    wire N__48610;
    wire N__48599;
    wire N__48596;
    wire N__48587;
    wire N__48580;
    wire N__48571;
    wire N__48568;
    wire N__48557;
    wire N__48554;
    wire N__48549;
    wire N__48522;
    wire N__48519;
    wire N__48516;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48495;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48471;
    wire N__48468;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48444;
    wire N__48441;
    wire N__48438;
    wire N__48435;
    wire N__48432;
    wire N__48429;
    wire N__48426;
    wire N__48423;
    wire N__48420;
    wire N__48417;
    wire N__48414;
    wire N__48411;
    wire N__48408;
    wire N__48405;
    wire N__48402;
    wire N__48399;
    wire N__48396;
    wire N__48393;
    wire N__48390;
    wire N__48387;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48375;
    wire N__48372;
    wire N__48369;
    wire N__48366;
    wire N__48363;
    wire N__48360;
    wire N__48357;
    wire N__48354;
    wire N__48351;
    wire N__48348;
    wire N__48345;
    wire N__48342;
    wire N__48339;
    wire N__48336;
    wire N__48333;
    wire N__48330;
    wire N__48327;
    wire N__48326;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48314;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48297;
    wire N__48296;
    wire N__48293;
    wire N__48292;
    wire N__48291;
    wire N__48290;
    wire N__48287;
    wire N__48286;
    wire N__48285;
    wire N__48282;
    wire N__48279;
    wire N__48276;
    wire N__48275;
    wire N__48274;
    wire N__48269;
    wire N__48264;
    wire N__48259;
    wire N__48256;
    wire N__48251;
    wire N__48240;
    wire N__48237;
    wire N__48236;
    wire N__48233;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48223;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48204;
    wire N__48201;
    wire N__48198;
    wire N__48195;
    wire N__48192;
    wire N__48189;
    wire N__48186;
    wire N__48183;
    wire N__48180;
    wire N__48177;
    wire N__48174;
    wire N__48171;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48159;
    wire N__48156;
    wire N__48153;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48132;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48120;
    wire N__48117;
    wire N__48114;
    wire N__48111;
    wire N__48108;
    wire N__48105;
    wire N__48102;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48086;
    wire N__48085;
    wire N__48084;
    wire N__48081;
    wire N__48074;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48062;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48047;
    wire N__48044;
    wire N__48041;
    wire N__48036;
    wire N__48035;
    wire N__48032;
    wire N__48029;
    wire N__48026;
    wire N__48025;
    wire N__48022;
    wire N__48021;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48008;
    wire N__48005;
    wire N__47994;
    wire N__47991;
    wire N__47988;
    wire N__47987;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47983;
    wire N__47982;
    wire N__47979;
    wire N__47976;
    wire N__47973;
    wire N__47970;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47946;
    wire N__47945;
    wire N__47942;
    wire N__47939;
    wire N__47936;
    wire N__47933;
    wire N__47930;
    wire N__47927;
    wire N__47924;
    wire N__47921;
    wire N__47916;
    wire N__47913;
    wire N__47912;
    wire N__47909;
    wire N__47906;
    wire N__47905;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47873;
    wire N__47872;
    wire N__47871;
    wire N__47870;
    wire N__47869;
    wire N__47866;
    wire N__47863;
    wire N__47854;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47838;
    wire N__47837;
    wire N__47836;
    wire N__47833;
    wire N__47828;
    wire N__47823;
    wire N__47822;
    wire N__47819;
    wire N__47816;
    wire N__47815;
    wire N__47812;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47796;
    wire N__47793;
    wire N__47790;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47762;
    wire N__47761;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47745;
    wire N__47742;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47731;
    wire N__47728;
    wire N__47725;
    wire N__47722;
    wire N__47715;
    wire N__47712;
    wire N__47711;
    wire N__47710;
    wire N__47709;
    wire N__47706;
    wire N__47705;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47691;
    wire N__47688;
    wire N__47685;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47677;
    wire N__47674;
    wire N__47671;
    wire N__47668;
    wire N__47665;
    wire N__47662;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47652;
    wire N__47649;
    wire N__47644;
    wire N__47641;
    wire N__47636;
    wire N__47631;
    wire N__47622;
    wire N__47621;
    wire N__47620;
    wire N__47619;
    wire N__47618;
    wire N__47617;
    wire N__47614;
    wire N__47611;
    wire N__47600;
    wire N__47597;
    wire N__47592;
    wire N__47589;
    wire N__47586;
    wire N__47583;
    wire N__47582;
    wire N__47581;
    wire N__47580;
    wire N__47579;
    wire N__47578;
    wire N__47577;
    wire N__47564;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47554;
    wire N__47553;
    wire N__47552;
    wire N__47551;
    wire N__47548;
    wire N__47545;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47472;
    wire N__47469;
    wire N__47468;
    wire N__47467;
    wire N__47466;
    wire N__47465;
    wire N__47464;
    wire N__47463;
    wire N__47462;
    wire N__47461;
    wire N__47458;
    wire N__47457;
    wire N__47456;
    wire N__47453;
    wire N__47448;
    wire N__47441;
    wire N__47436;
    wire N__47433;
    wire N__47428;
    wire N__47425;
    wire N__47424;
    wire N__47423;
    wire N__47422;
    wire N__47421;
    wire N__47420;
    wire N__47419;
    wire N__47418;
    wire N__47417;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47394;
    wire N__47387;
    wire N__47384;
    wire N__47381;
    wire N__47378;
    wire N__47375;
    wire N__47372;
    wire N__47369;
    wire N__47352;
    wire N__47351;
    wire N__47350;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47344;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47327;
    wire N__47324;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47318;
    wire N__47317;
    wire N__47316;
    wire N__47315;
    wire N__47308;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47287;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47256;
    wire N__47253;
    wire N__47248;
    wire N__47245;
    wire N__47242;
    wire N__47241;
    wire N__47236;
    wire N__47233;
    wire N__47230;
    wire N__47225;
    wire N__47218;
    wire N__47215;
    wire N__47210;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47189;
    wire N__47188;
    wire N__47181;
    wire N__47178;
    wire N__47177;
    wire N__47174;
    wire N__47173;
    wire N__47172;
    wire N__47171;
    wire N__47170;
    wire N__47169;
    wire N__47166;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47162;
    wire N__47161;
    wire N__47158;
    wire N__47153;
    wire N__47152;
    wire N__47151;
    wire N__47150;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47128;
    wire N__47127;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47115;
    wire N__47110;
    wire N__47109;
    wire N__47106;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47084;
    wire N__47081;
    wire N__47072;
    wire N__47069;
    wire N__47064;
    wire N__47061;
    wire N__47054;
    wire N__47051;
    wire N__47040;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47032;
    wire N__47029;
    wire N__47026;
    wire N__47023;
    wire N__47020;
    wire N__47017;
    wire N__47014;
    wire N__47009;
    wire N__47004;
    wire N__47001;
    wire N__47000;
    wire N__46997;
    wire N__46994;
    wire N__46993;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46953;
    wire N__46952;
    wire N__46951;
    wire N__46948;
    wire N__46945;
    wire N__46942;
    wire N__46937;
    wire N__46932;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46920;
    wire N__46919;
    wire N__46914;
    wire N__46911;
    wire N__46908;
    wire N__46907;
    wire N__46906;
    wire N__46901;
    wire N__46900;
    wire N__46897;
    wire N__46894;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46880;
    wire N__46875;
    wire N__46872;
    wire N__46869;
    wire N__46866;
    wire N__46865;
    wire N__46862;
    wire N__46859;
    wire N__46856;
    wire N__46851;
    wire N__46850;
    wire N__46847;
    wire N__46844;
    wire N__46841;
    wire N__46838;
    wire N__46835;
    wire N__46832;
    wire N__46829;
    wire N__46824;
    wire N__46821;
    wire N__46818;
    wire N__46817;
    wire N__46814;
    wire N__46811;
    wire N__46808;
    wire N__46805;
    wire N__46800;
    wire N__46797;
    wire N__46796;
    wire N__46793;
    wire N__46790;
    wire N__46787;
    wire N__46782;
    wire N__46781;
    wire N__46778;
    wire N__46777;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46764;
    wire N__46763;
    wire N__46762;
    wire N__46759;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46735;
    wire N__46732;
    wire N__46727;
    wire N__46724;
    wire N__46721;
    wire N__46716;
    wire N__46713;
    wire N__46712;
    wire N__46709;
    wire N__46708;
    wire N__46705;
    wire N__46702;
    wire N__46699;
    wire N__46692;
    wire N__46689;
    wire N__46686;
    wire N__46685;
    wire N__46684;
    wire N__46677;
    wire N__46676;
    wire N__46673;
    wire N__46670;
    wire N__46665;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46653;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46595;
    wire N__46592;
    wire N__46587;
    wire N__46586;
    wire N__46585;
    wire N__46578;
    wire N__46575;
    wire N__46574;
    wire N__46573;
    wire N__46572;
    wire N__46571;
    wire N__46570;
    wire N__46569;
    wire N__46568;
    wire N__46567;
    wire N__46566;
    wire N__46565;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46555;
    wire N__46554;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46544;
    wire N__46541;
    wire N__46536;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46520;
    wire N__46513;
    wire N__46510;
    wire N__46505;
    wire N__46502;
    wire N__46501;
    wire N__46498;
    wire N__46495;
    wire N__46492;
    wire N__46485;
    wire N__46480;
    wire N__46477;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46455;
    wire N__46454;
    wire N__46453;
    wire N__46450;
    wire N__46449;
    wire N__46448;
    wire N__46447;
    wire N__46446;
    wire N__46445;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46437;
    wire N__46436;
    wire N__46433;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46407;
    wire N__46404;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46389;
    wire N__46388;
    wire N__46383;
    wire N__46378;
    wire N__46371;
    wire N__46366;
    wire N__46361;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46353;
    wire N__46352;
    wire N__46349;
    wire N__46344;
    wire N__46341;
    wire N__46336;
    wire N__46333;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46318;
    wire N__46313;
    wire N__46302;
    wire N__46301;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46291;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46269;
    wire N__46266;
    wire N__46263;
    wire N__46260;
    wire N__46257;
    wire N__46254;
    wire N__46253;
    wire N__46250;
    wire N__46247;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46232;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46219;
    wire N__46216;
    wire N__46213;
    wire N__46208;
    wire N__46203;
    wire N__46200;
    wire N__46199;
    wire N__46198;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46151;
    wire N__46148;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46127;
    wire N__46126;
    wire N__46123;
    wire N__46118;
    wire N__46113;
    wire N__46112;
    wire N__46109;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46070;
    wire N__46067;
    wire N__46064;
    wire N__46063;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46051;
    wire N__46044;
    wire N__46041;
    wire N__46040;
    wire N__46037;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46022;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46004;
    wire N__46001;
    wire N__45998;
    wire N__45995;
    wire N__45992;
    wire N__45989;
    wire N__45984;
    wire N__45983;
    wire N__45982;
    wire N__45975;
    wire N__45972;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45893;
    wire N__45892;
    wire N__45889;
    wire N__45884;
    wire N__45879;
    wire N__45878;
    wire N__45875;
    wire N__45874;
    wire N__45871;
    wire N__45870;
    wire N__45867;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45779;
    wire N__45778;
    wire N__45775;
    wire N__45772;
    wire N__45769;
    wire N__45766;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45752;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45735;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45701;
    wire N__45700;
    wire N__45699;
    wire N__45698;
    wire N__45697;
    wire N__45696;
    wire N__45695;
    wire N__45694;
    wire N__45691;
    wire N__45688;
    wire N__45675;
    wire N__45672;
    wire N__45663;
    wire N__45662;
    wire N__45661;
    wire N__45658;
    wire N__45653;
    wire N__45648;
    wire N__45645;
    wire N__45644;
    wire N__45643;
    wire N__45638;
    wire N__45635;
    wire N__45632;
    wire N__45627;
    wire N__45626;
    wire N__45625;
    wire N__45618;
    wire N__45615;
    wire N__45614;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45575;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45560;
    wire N__45559;
    wire N__45558;
    wire N__45557;
    wire N__45554;
    wire N__45553;
    wire N__45550;
    wire N__45547;
    wire N__45546;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45536;
    wire N__45533;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45516;
    wire N__45515;
    wire N__45514;
    wire N__45513;
    wire N__45510;
    wire N__45505;
    wire N__45504;
    wire N__45503;
    wire N__45500;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45483;
    wire N__45480;
    wire N__45477;
    wire N__45474;
    wire N__45469;
    wire N__45464;
    wire N__45461;
    wire N__45452;
    wire N__45449;
    wire N__45444;
    wire N__45429;
    wire N__45428;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45413;
    wire N__45410;
    wire N__45405;
    wire N__45404;
    wire N__45403;
    wire N__45402;
    wire N__45401;
    wire N__45400;
    wire N__45399;
    wire N__45398;
    wire N__45397;
    wire N__45396;
    wire N__45395;
    wire N__45394;
    wire N__45391;
    wire N__45390;
    wire N__45389;
    wire N__45388;
    wire N__45387;
    wire N__45386;
    wire N__45385;
    wire N__45382;
    wire N__45381;
    wire N__45380;
    wire N__45377;
    wire N__45376;
    wire N__45375;
    wire N__45374;
    wire N__45373;
    wire N__45372;
    wire N__45371;
    wire N__45370;
    wire N__45367;
    wire N__45364;
    wire N__45363;
    wire N__45362;
    wire N__45359;
    wire N__45358;
    wire N__45355;
    wire N__45354;
    wire N__45351;
    wire N__45348;
    wire N__45345;
    wire N__45344;
    wire N__45343;
    wire N__45342;
    wire N__45341;
    wire N__45340;
    wire N__45337;
    wire N__45334;
    wire N__45333;
    wire N__45330;
    wire N__45325;
    wire N__45322;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45314;
    wire N__45311;
    wire N__45306;
    wire N__45299;
    wire N__45298;
    wire N__45297;
    wire N__45296;
    wire N__45295;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45262;
    wire N__45257;
    wire N__45252;
    wire N__45241;
    wire N__45230;
    wire N__45225;
    wire N__45222;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45204;
    wire N__45203;
    wire N__45202;
    wire N__45201;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45190;
    wire N__45187;
    wire N__45186;
    wire N__45181;
    wire N__45174;
    wire N__45169;
    wire N__45164;
    wire N__45159;
    wire N__45144;
    wire N__45141;
    wire N__45136;
    wire N__45133;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45115;
    wire N__45110;
    wire N__45107;
    wire N__45098;
    wire N__45095;
    wire N__45088;
    wire N__45081;
    wire N__45076;
    wire N__45071;
    wire N__45066;
    wire N__45057;
    wire N__45056;
    wire N__45053;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45033;
    wire N__45032;
    wire N__45029;
    wire N__45026;
    wire N__45025;
    wire N__45022;
    wire N__45017;
    wire N__45012;
    wire N__45011;
    wire N__45008;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44984;
    wire N__44981;
    wire N__44980;
    wire N__44979;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44971;
    wire N__44970;
    wire N__44967;
    wire N__44966;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44952;
    wire N__44951;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44935;
    wire N__44932;
    wire N__44929;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44891;
    wire N__44888;
    wire N__44881;
    wire N__44878;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44858;
    wire N__44855;
    wire N__44854;
    wire N__44847;
    wire N__44844;
    wire N__44843;
    wire N__44840;
    wire N__44837;
    wire N__44832;
    wire N__44831;
    wire N__44830;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44816;
    wire N__44813;
    wire N__44810;
    wire N__44807;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44792;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44771;
    wire N__44766;
    wire N__44765;
    wire N__44762;
    wire N__44759;
    wire N__44756;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44736;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44726;
    wire N__44725;
    wire N__44722;
    wire N__44721;
    wire N__44720;
    wire N__44717;
    wire N__44714;
    wire N__44707;
    wire N__44706;
    wire N__44705;
    wire N__44704;
    wire N__44703;
    wire N__44698;
    wire N__44695;
    wire N__44686;
    wire N__44685;
    wire N__44684;
    wire N__44683;
    wire N__44682;
    wire N__44681;
    wire N__44678;
    wire N__44675;
    wire N__44672;
    wire N__44661;
    wire N__44660;
    wire N__44657;
    wire N__44650;
    wire N__44647;
    wire N__44640;
    wire N__44637;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44612;
    wire N__44609;
    wire N__44606;
    wire N__44603;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44592;
    wire N__44589;
    wire N__44584;
    wire N__44581;
    wire N__44580;
    wire N__44577;
    wire N__44572;
    wire N__44569;
    wire N__44566;
    wire N__44563;
    wire N__44560;
    wire N__44553;
    wire N__44552;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44531;
    wire N__44528;
    wire N__44523;
    wire N__44520;
    wire N__44519;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44496;
    wire N__44493;
    wire N__44492;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44471;
    wire N__44468;
    wire N__44463;
    wire N__44460;
    wire N__44459;
    wire N__44456;
    wire N__44455;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44439;
    wire N__44438;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44417;
    wire N__44414;
    wire N__44411;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44351;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44276;
    wire N__44273;
    wire N__44270;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44237;
    wire N__44234;
    wire N__44231;
    wire N__44226;
    wire N__44225;
    wire N__44220;
    wire N__44217;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44202;
    wire N__44201;
    wire N__44200;
    wire N__44199;
    wire N__44196;
    wire N__44195;
    wire N__44194;
    wire N__44191;
    wire N__44190;
    wire N__44189;
    wire N__44186;
    wire N__44183;
    wire N__44180;
    wire N__44177;
    wire N__44174;
    wire N__44171;
    wire N__44170;
    wire N__44167;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44159;
    wire N__44156;
    wire N__44153;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44126;
    wire N__44125;
    wire N__44124;
    wire N__44123;
    wire N__44120;
    wire N__44117;
    wire N__44108;
    wire N__44101;
    wire N__44096;
    wire N__44093;
    wire N__44088;
    wire N__44073;
    wire N__44072;
    wire N__44071;
    wire N__44070;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44059;
    wire N__44058;
    wire N__44055;
    wire N__44054;
    wire N__44053;
    wire N__44050;
    wire N__44049;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44021;
    wire N__44020;
    wire N__44015;
    wire N__44012;
    wire N__44005;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43980;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43916;
    wire N__43915;
    wire N__43912;
    wire N__43907;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43886;
    wire N__43883;
    wire N__43880;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43865;
    wire N__43864;
    wire N__43857;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43842;
    wire N__43841;
    wire N__43838;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43793;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43745;
    wire N__43744;
    wire N__43743;
    wire N__43740;
    wire N__43733;
    wire N__43728;
    wire N__43725;
    wire N__43724;
    wire N__43723;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43711;
    wire N__43704;
    wire N__43703;
    wire N__43700;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43692;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43677;
    wire N__43668;
    wire N__43667;
    wire N__43664;
    wire N__43661;
    wire N__43660;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43618;
    wire N__43615;
    wire N__43612;
    wire N__43609;
    wire N__43608;
    wire N__43605;
    wire N__43600;
    wire N__43597;
    wire N__43590;
    wire N__43587;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43575;
    wire N__43574;
    wire N__43573;
    wire N__43570;
    wire N__43565;
    wire N__43560;
    wire N__43557;
    wire N__43556;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43538;
    wire N__43537;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43517;
    wire N__43512;
    wire N__43511;
    wire N__43510;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43494;
    wire N__43485;
    wire N__43484;
    wire N__43483;
    wire N__43482;
    wire N__43481;
    wire N__43480;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43468;
    wire N__43463;
    wire N__43460;
    wire N__43449;
    wire N__43446;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43438;
    wire N__43437;
    wire N__43436;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43424;
    wire N__43419;
    wire N__43410;
    wire N__43409;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43389;
    wire N__43388;
    wire N__43387;
    wire N__43384;
    wire N__43383;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43373;
    wire N__43368;
    wire N__43359;
    wire N__43358;
    wire N__43357;
    wire N__43356;
    wire N__43355;
    wire N__43352;
    wire N__43351;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43337;
    wire N__43332;
    wire N__43327;
    wire N__43320;
    wire N__43317;
    wire N__43316;
    wire N__43313;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43289;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43275;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43256;
    wire N__43253;
    wire N__43248;
    wire N__43247;
    wire N__43244;
    wire N__43241;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43216;
    wire N__43211;
    wire N__43208;
    wire N__43205;
    wire N__43200;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43157;
    wire N__43156;
    wire N__43153;
    wire N__43148;
    wire N__43143;
    wire N__43142;
    wire N__43141;
    wire N__43138;
    wire N__43133;
    wire N__43128;
    wire N__43125;
    wire N__43124;
    wire N__43121;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43104;
    wire N__43103;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43083;
    wire N__43082;
    wire N__43079;
    wire N__43074;
    wire N__43071;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43055;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43033;
    wire N__43028;
    wire N__43025;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43011;
    wire N__43010;
    wire N__43007;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42983;
    wire N__42978;
    wire N__42975;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42930;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42916;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42885;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42871;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42854;
    wire N__42849;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42810;
    wire N__42809;
    wire N__42808;
    wire N__42805;
    wire N__42802;
    wire N__42799;
    wire N__42796;
    wire N__42789;
    wire N__42788;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42778;
    wire N__42771;
    wire N__42770;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42747;
    wire N__42746;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42719;
    wire N__42718;
    wire N__42715;
    wire N__42712;
    wire N__42709;
    wire N__42706;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42692;
    wire N__42691;
    wire N__42688;
    wire N__42685;
    wire N__42682;
    wire N__42679;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42635;
    wire N__42634;
    wire N__42633;
    wire N__42632;
    wire N__42629;
    wire N__42628;
    wire N__42627;
    wire N__42622;
    wire N__42617;
    wire N__42614;
    wire N__42611;
    wire N__42610;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42598;
    wire N__42595;
    wire N__42590;
    wire N__42587;
    wire N__42582;
    wire N__42579;
    wire N__42572;
    wire N__42567;
    wire N__42566;
    wire N__42563;
    wire N__42562;
    wire N__42561;
    wire N__42556;
    wire N__42553;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42539;
    wire N__42536;
    wire N__42531;
    wire N__42526;
    wire N__42521;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42491;
    wire N__42488;
    wire N__42485;
    wire N__42480;
    wire N__42477;
    wire N__42476;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42458;
    wire N__42457;
    wire N__42454;
    wire N__42451;
    wire N__42450;
    wire N__42449;
    wire N__42448;
    wire N__42447;
    wire N__42446;
    wire N__42443;
    wire N__42442;
    wire N__42441;
    wire N__42440;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42392;
    wire N__42389;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42367;
    wire N__42366;
    wire N__42365;
    wire N__42364;
    wire N__42363;
    wire N__42356;
    wire N__42353;
    wire N__42352;
    wire N__42347;
    wire N__42340;
    wire N__42337;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42326;
    wire N__42321;
    wire N__42318;
    wire N__42317;
    wire N__42316;
    wire N__42315;
    wire N__42310;
    wire N__42307;
    wire N__42300;
    wire N__42299;
    wire N__42298;
    wire N__42297;
    wire N__42296;
    wire N__42295;
    wire N__42292;
    wire N__42289;
    wire N__42288;
    wire N__42287;
    wire N__42286;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42262;
    wire N__42259;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42241;
    wire N__42238;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42230;
    wire N__42229;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42189;
    wire N__42184;
    wire N__42181;
    wire N__42176;
    wire N__42173;
    wire N__42170;
    wire N__42167;
    wire N__42164;
    wire N__42161;
    wire N__42156;
    wire N__42153;
    wire N__42148;
    wire N__42139;
    wire N__42134;
    wire N__42127;
    wire N__42124;
    wire N__42119;
    wire N__42114;
    wire N__42109;
    wire N__42104;
    wire N__42095;
    wire N__42092;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42077;
    wire N__42076;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42064;
    wire N__42057;
    wire N__42056;
    wire N__42053;
    wire N__42052;
    wire N__42051;
    wire N__42048;
    wire N__42045;
    wire N__42040;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42026;
    wire N__42025;
    wire N__42022;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42010;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41945;
    wire N__41944;
    wire N__41941;
    wire N__41938;
    wire N__41935;
    wire N__41932;
    wire N__41925;
    wire N__41922;
    wire N__41921;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41911;
    wire N__41908;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41873;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41858;
    wire N__41853;
    wire N__41852;
    wire N__41849;
    wire N__41848;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41721;
    wire N__41718;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41550;
    wire N__41547;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41510;
    wire N__41509;
    wire N__41506;
    wire N__41501;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41480;
    wire N__41477;
    wire N__41474;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41462;
    wire N__41461;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41435;
    wire N__41432;
    wire N__41429;
    wire N__41426;
    wire N__41423;
    wire N__41418;
    wire N__41415;
    wire N__41412;
    wire N__41411;
    wire N__41410;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41357;
    wire N__41356;
    wire N__41355;
    wire N__41354;
    wire N__41353;
    wire N__41352;
    wire N__41349;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41332;
    wire N__41329;
    wire N__41328;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41313;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41286;
    wire N__41281;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41224;
    wire N__41217;
    wire N__41214;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41206;
    wire N__41201;
    wire N__41198;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41175;
    wire N__41174;
    wire N__41173;
    wire N__41170;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41148;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41091;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41045;
    wire N__41044;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41010;
    wire N__41009;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40990;
    wire N__40983;
    wire N__40982;
    wire N__40981;
    wire N__40980;
    wire N__40979;
    wire N__40976;
    wire N__40975;
    wire N__40974;
    wire N__40971;
    wire N__40970;
    wire N__40969;
    wire N__40968;
    wire N__40965;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40945;
    wire N__40944;
    wire N__40943;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40924;
    wire N__40919;
    wire N__40914;
    wire N__40909;
    wire N__40906;
    wire N__40897;
    wire N__40894;
    wire N__40891;
    wire N__40882;
    wire N__40875;
    wire N__40872;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40850;
    wire N__40849;
    wire N__40846;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40754;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40721;
    wire N__40718;
    wire N__40715;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40662;
    wire N__40659;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40610;
    wire N__40607;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40577;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40562;
    wire N__40557;
    wire N__40554;
    wire N__40553;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40527;
    wire N__40526;
    wire N__40521;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40506;
    wire N__40503;
    wire N__40502;
    wire N__40497;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40475;
    wire N__40470;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40455;
    wire N__40454;
    wire N__40453;
    wire N__40450;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40434;
    wire N__40431;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40418;
    wire N__40417;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40397;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40364;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40343;
    wire N__40342;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40314;
    wire N__40311;
    wire N__40310;
    wire N__40309;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40292;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40266;
    wire N__40265;
    wire N__40264;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40250;
    wire N__40249;
    wire N__40246;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40230;
    wire N__40227;
    wire N__40226;
    wire N__40225;
    wire N__40222;
    wire N__40217;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40205;
    wire N__40204;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40172;
    wire N__40171;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40149;
    wire N__40148;
    wire N__40145;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40133;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40112;
    wire N__40111;
    wire N__40104;
    wire N__40101;
    wire N__40100;
    wire N__40099;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40071;
    wire N__40068;
    wire N__40065;
    wire N__40064;
    wire N__40063;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40046;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40022;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__40001;
    wire N__40000;
    wire N__39997;
    wire N__39992;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39980;
    wire N__39975;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39965;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39953;
    wire N__39952;
    wire N__39947;
    wire N__39944;
    wire N__39941;
    wire N__39938;
    wire N__39935;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39908;
    wire N__39907;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39890;
    wire N__39887;
    wire N__39884;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39860;
    wire N__39859;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39783;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39749;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39737;
    wire N__39736;
    wire N__39735;
    wire N__39732;
    wire N__39731;
    wire N__39730;
    wire N__39729;
    wire N__39728;
    wire N__39727;
    wire N__39726;
    wire N__39725;
    wire N__39724;
    wire N__39723;
    wire N__39722;
    wire N__39721;
    wire N__39720;
    wire N__39719;
    wire N__39718;
    wire N__39717;
    wire N__39706;
    wire N__39701;
    wire N__39686;
    wire N__39679;
    wire N__39678;
    wire N__39677;
    wire N__39676;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39650;
    wire N__39647;
    wire N__39642;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39607;
    wire N__39600;
    wire N__39599;
    wire N__39596;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39588;
    wire N__39585;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39564;
    wire N__39559;
    wire N__39552;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39542;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39528;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39467;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39410;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39398;
    wire N__39397;
    wire N__39394;
    wire N__39389;
    wire N__39384;
    wire N__39383;
    wire N__39380;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39239;
    wire N__39236;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39194;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39095;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39047;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38993;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38975;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38939;
    wire N__38936;
    wire N__38933;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38876;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38819;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38717;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38553;
    wire N__38552;
    wire N__38551;
    wire N__38546;
    wire N__38543;
    wire N__38540;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38528;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38507;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38490;
    wire N__38487;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38457;
    wire N__38454;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38430;
    wire N__38429;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38396;
    wire N__38393;
    wire N__38390;
    wire N__38387;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38362;
    wire N__38357;
    wire N__38352;
    wire N__38349;
    wire N__38348;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38325;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38303;
    wire N__38298;
    wire N__38295;
    wire N__38294;
    wire N__38293;
    wire N__38290;
    wire N__38285;
    wire N__38280;
    wire N__38279;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38258;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38235;
    wire N__38232;
    wire N__38231;
    wire N__38230;
    wire N__38225;
    wire N__38222;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38202;
    wire N__38201;
    wire N__38196;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38171;
    wire N__38170;
    wire N__38167;
    wire N__38162;
    wire N__38157;
    wire N__38154;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38122;
    wire N__38119;
    wire N__38114;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38102;
    wire N__38099;
    wire N__38096;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38081;
    wire N__38078;
    wire N__38075;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38048;
    wire N__38047;
    wire N__38046;
    wire N__38041;
    wire N__38036;
    wire N__38033;
    wire N__38030;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37995;
    wire N__37994;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37955;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37916;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37813;
    wire N__37808;
    wire N__37805;
    wire N__37802;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37743;
    wire N__37740;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37578;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37559;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37544;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37530;
    wire N__37529;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37514;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37467;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37453;
    wire N__37448;
    wire N__37445;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37388;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37373;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37361;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37307;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37188;
    wire N__37185;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37142;
    wire N__37141;
    wire N__37140;
    wire N__37139;
    wire N__37136;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37110;
    wire N__37105;
    wire N__37102;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37062;
    wire N__37059;
    wire N__37056;
    wire N__37055;
    wire N__37054;
    wire N__37053;
    wire N__37050;
    wire N__37043;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37004;
    wire N__37003;
    wire N__37002;
    wire N__36999;
    wire N__36992;
    wire N__36987;
    wire N__36984;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36949;
    wire N__36948;
    wire N__36943;
    wire N__36942;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36885;
    wire N__36882;
    wire N__36879;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36852;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36731;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36725;
    wire N__36724;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36712;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36690;
    wire N__36687;
    wire N__36686;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36678;
    wire N__36675;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36655;
    wire N__36650;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36626;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36609;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36581;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36565;
    wire N__36562;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36452;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36371;
    wire N__36370;
    wire N__36369;
    wire N__36366;
    wire N__36359;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36315;
    wire N__36312;
    wire N__36311;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36290;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36278;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36263;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36215;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36186;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36153;
    wire N__36152;
    wire N__36149;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36125;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36069;
    wire N__36066;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36058;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35971;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35787;
    wire N__35784;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35730;
    wire N__35727;
    wire N__35724;
    wire N__35721;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35684;
    wire N__35679;
    wire N__35676;
    wire N__35675;
    wire N__35674;
    wire N__35671;
    wire N__35666;
    wire N__35661;
    wire N__35658;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35646;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35634;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35596;
    wire N__35591;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35577;
    wire N__35576;
    wire N__35573;
    wire N__35572;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35564;
    wire N__35561;
    wire N__35560;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35547;
    wire N__35542;
    wire N__35539;
    wire N__35538;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35526;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35502;
    wire N__35499;
    wire N__35498;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35487;
    wire N__35486;
    wire N__35485;
    wire N__35484;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35469;
    wire N__35466;
    wire N__35465;
    wire N__35464;
    wire N__35459;
    wire N__35456;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35430;
    wire N__35427;
    wire N__35426;
    wire N__35423;
    wire N__35422;
    wire N__35421;
    wire N__35420;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35390;
    wire N__35389;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35349;
    wire N__35346;
    wire N__35343;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35330;
    wire N__35327;
    wire N__35326;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35318;
    wire N__35313;
    wire N__35308;
    wire N__35305;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35280;
    wire N__35277;
    wire N__35276;
    wire N__35275;
    wire N__35274;
    wire N__35273;
    wire N__35272;
    wire N__35271;
    wire N__35270;
    wire N__35269;
    wire N__35266;
    wire N__35253;
    wire N__35248;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35230;
    wire N__35225;
    wire N__35220;
    wire N__35219;
    wire N__35216;
    wire N__35213;
    wire N__35210;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35193;
    wire N__35190;
    wire N__35189;
    wire N__35188;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35170;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35153;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35129;
    wire N__35128;
    wire N__35125;
    wire N__35120;
    wire N__35119;
    wire N__35114;
    wire N__35111;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35066;
    wire N__35065;
    wire N__35058;
    wire N__35055;
    wire N__35054;
    wire N__35053;
    wire N__35052;
    wire N__35043;
    wire N__35040;
    wire N__35039;
    wire N__35038;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35026;
    wire N__35023;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire N__35009;
    wire N__35008;
    wire N__35007;
    wire N__35004;
    wire N__35001;
    wire N__34996;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34979;
    wire N__34978;
    wire N__34977;
    wire N__34974;
    wire N__34967;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34703;
    wire N__34698;
    wire N__34695;
    wire N__34694;
    wire N__34693;
    wire N__34692;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34674;
    wire N__34667;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34649;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34580;
    wire N__34579;
    wire N__34576;
    wire N__34571;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34559;
    wire N__34556;
    wire N__34555;
    wire N__34552;
    wire N__34547;
    wire N__34542;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34527;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34512;
    wire N__34509;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34494;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34479;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34467;
    wire N__34464;
    wire N__34463;
    wire N__34458;
    wire N__34455;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34443;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34421;
    wire N__34420;
    wire N__34417;
    wire N__34412;
    wire N__34407;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34395;
    wire N__34394;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34382;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34370;
    wire N__34367;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34354;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34313;
    wire N__34310;
    wire N__34307;
    wire N__34302;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34290;
    wire N__34287;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34275;
    wire N__34274;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34262;
    wire N__34261;
    wire N__34254;
    wire N__34251;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34239;
    wire N__34238;
    wire N__34233;
    wire N__34230;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34218;
    wire N__34217;
    wire N__34214;
    wire N__34209;
    wire N__34206;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34056;
    wire N__34053;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34041;
    wire N__34038;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34026;
    wire N__34023;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34011;
    wire N__34008;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33972;
    wire N__33969;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33944;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33928;
    wire N__33923;
    wire N__33920;
    wire N__33919;
    wire N__33918;
    wire N__33913;
    wire N__33912;
    wire N__33911;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33891;
    wire N__33882;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33874;
    wire N__33869;
    wire N__33866;
    wire N__33861;
    wire N__33860;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33852;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33837;
    wire N__33836;
    wire N__33831;
    wire N__33826;
    wire N__33825;
    wire N__33822;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33807;
    wire N__33798;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33790;
    wire N__33789;
    wire N__33788;
    wire N__33787;
    wire N__33786;
    wire N__33785;
    wire N__33782;
    wire N__33777;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33752;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33723;
    wire N__33722;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33705;
    wire N__33704;
    wire N__33703;
    wire N__33702;
    wire N__33699;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33681;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33648;
    wire N__33645;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33609;
    wire N__33606;
    wire N__33605;
    wire N__33604;
    wire N__33601;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33585;
    wire N__33582;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33536;
    wire N__33535;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33498;
    wire N__33497;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33473;
    wire N__33468;
    wire N__33465;
    wire N__33464;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33428;
    wire N__33425;
    wire N__33424;
    wire N__33421;
    wire N__33420;
    wire N__33417;
    wire N__33412;
    wire N__33409;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33389;
    wire N__33388;
    wire N__33387;
    wire N__33386;
    wire N__33385;
    wire N__33382;
    wire N__33371;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33342;
    wire N__33339;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33331;
    wire N__33330;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33310;
    wire N__33307;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33276;
    wire N__33273;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33249;
    wire N__33246;
    wire N__33245;
    wire N__33242;
    wire N__33241;
    wire N__33238;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33219;
    wire N__33218;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33197;
    wire N__33192;
    wire N__33189;
    wire N__33188;
    wire N__33183;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33143;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33120;
    wire N__33117;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33109;
    wire N__33108;
    wire N__33107;
    wire N__33102;
    wire N__33099;
    wire N__33094;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33012;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32997;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32985;
    wire N__32982;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32945;
    wire N__32942;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32893;
    wire N__32892;
    wire N__32891;
    wire N__32890;
    wire N__32889;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32865;
    wire N__32864;
    wire N__32861;
    wire N__32860;
    wire N__32859;
    wire N__32856;
    wire N__32851;
    wire N__32848;
    wire N__32843;
    wire N__32840;
    wire N__32835;
    wire N__32832;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32820;
    wire N__32819;
    wire N__32818;
    wire N__32817;
    wire N__32816;
    wire N__32807;
    wire N__32798;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32763;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32748;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32733;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32718;
    wire N__32715;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32687;
    wire N__32686;
    wire N__32679;
    wire N__32676;
    wire N__32675;
    wire N__32674;
    wire N__32669;
    wire N__32666;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32625;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32613;
    wire N__32610;
    wire N__32609;
    wire N__32608;
    wire N__32607;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32577;
    wire N__32576;
    wire N__32571;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32555;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32525;
    wire N__32520;
    wire N__32519;
    wire N__32518;
    wire N__32515;
    wire N__32510;
    wire N__32505;
    wire N__32504;
    wire N__32501;
    wire N__32500;
    wire N__32495;
    wire N__32492;
    wire N__32491;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32450;
    wire N__32445;
    wire N__32442;
    wire N__32441;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32378;
    wire N__32377;
    wire N__32372;
    wire N__32369;
    wire N__32364;
    wire N__32361;
    wire N__32360;
    wire N__32359;
    wire N__32352;
    wire N__32349;
    wire N__32348;
    wire N__32347;
    wire N__32344;
    wire N__32339;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32309;
    wire N__32306;
    wire N__32305;
    wire N__32304;
    wire N__32301;
    wire N__32296;
    wire N__32293;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32268;
    wire N__32267;
    wire N__32266;
    wire N__32263;
    wire N__32262;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32243;
    wire N__32240;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32213;
    wire N__32212;
    wire N__32209;
    wire N__32208;
    wire N__32207;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32192;
    wire N__32189;
    wire N__32178;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32156;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32076;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32010;
    wire N__32007;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31971;
    wire N__31968;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31914;
    wire N__31913;
    wire N__31910;
    wire N__31909;
    wire N__31908;
    wire N__31901;
    wire N__31898;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31886;
    wire N__31885;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31869;
    wire N__31866;
    wire N__31865;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31853;
    wire N__31850;
    wire N__31845;
    wire N__31842;
    wire N__31841;
    wire N__31840;
    wire N__31837;
    wire N__31832;
    wire N__31831;
    wire N__31826;
    wire N__31823;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31808;
    wire N__31805;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31790;
    wire N__31785;
    wire N__31784;
    wire N__31783;
    wire N__31782;
    wire N__31781;
    wire N__31780;
    wire N__31779;
    wire N__31778;
    wire N__31777;
    wire N__31776;
    wire N__31775;
    wire N__31774;
    wire N__31773;
    wire N__31772;
    wire N__31771;
    wire N__31768;
    wire N__31767;
    wire N__31766;
    wire N__31765;
    wire N__31764;
    wire N__31763;
    wire N__31762;
    wire N__31759;
    wire N__31754;
    wire N__31747;
    wire N__31742;
    wire N__31741;
    wire N__31740;
    wire N__31739;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31728;
    wire N__31727;
    wire N__31726;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31690;
    wire N__31687;
    wire N__31680;
    wire N__31679;
    wire N__31678;
    wire N__31675;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31663;
    wire N__31656;
    wire N__31655;
    wire N__31650;
    wire N__31647;
    wire N__31634;
    wire N__31629;
    wire N__31626;
    wire N__31621;
    wire N__31618;
    wire N__31613;
    wire N__31608;
    wire N__31605;
    wire N__31596;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31565;
    wire N__31560;
    wire N__31557;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31545;
    wire N__31544;
    wire N__31543;
    wire N__31540;
    wire N__31539;
    wire N__31534;
    wire N__31529;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31484;
    wire N__31483;
    wire N__31482;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31467;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31453;
    wire N__31450;
    wire N__31445;
    wire N__31440;
    wire N__31437;
    wire N__31436;
    wire N__31435;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31419;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31407;
    wire N__31406;
    wire N__31405;
    wire N__31402;
    wire N__31397;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31376;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31359;
    wire N__31358;
    wire N__31357;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31345;
    wire N__31338;
    wire N__31335;
    wire N__31334;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31317;
    wire N__31316;
    wire N__31315;
    wire N__31314;
    wire N__31313;
    wire N__31310;
    wire N__31309;
    wire N__31308;
    wire N__31307;
    wire N__31306;
    wire N__31305;
    wire N__31304;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31292;
    wire N__31291;
    wire N__31290;
    wire N__31287;
    wire N__31280;
    wire N__31275;
    wire N__31270;
    wire N__31269;
    wire N__31264;
    wire N__31261;
    wire N__31256;
    wire N__31253;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31234;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31119;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31109;
    wire N__31104;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31092;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31080;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31068;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31053;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31034;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31010;
    wire N__31005;
    wire N__31002;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30990;
    wire N__30987;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30962;
    wire N__30961;
    wire N__30956;
    wire N__30953;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30854;
    wire N__30851;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30833;
    wire N__30830;
    wire N__30825;
    wire N__30824;
    wire N__30823;
    wire N__30820;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30789;
    wire N__30788;
    wire N__30787;
    wire N__30782;
    wire N__30779;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30686;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30655;
    wire N__30650;
    wire N__30647;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30620;
    wire N__30619;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30598;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30563;
    wire N__30562;
    wire N__30561;
    wire N__30560;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30556;
    wire N__30553;
    wire N__30546;
    wire N__30535;
    wire N__30528;
    wire N__30527;
    wire N__30526;
    wire N__30525;
    wire N__30524;
    wire N__30523;
    wire N__30522;
    wire N__30521;
    wire N__30520;
    wire N__30519;
    wire N__30518;
    wire N__30505;
    wire N__30494;
    wire N__30489;
    wire N__30488;
    wire N__30487;
    wire N__30486;
    wire N__30485;
    wire N__30482;
    wire N__30481;
    wire N__30478;
    wire N__30477;
    wire N__30476;
    wire N__30473;
    wire N__30472;
    wire N__30469;
    wire N__30468;
    wire N__30457;
    wire N__30446;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30411;
    wire N__30408;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30396;
    wire N__30393;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30381;
    wire N__30380;
    wire N__30379;
    wire N__30378;
    wire N__30377;
    wire N__30376;
    wire N__30375;
    wire N__30374;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30344;
    wire N__30341;
    wire N__30340;
    wire N__30339;
    wire N__30338;
    wire N__30337;
    wire N__30336;
    wire N__30335;
    wire N__30334;
    wire N__30333;
    wire N__30330;
    wire N__30329;
    wire N__30328;
    wire N__30327;
    wire N__30326;
    wire N__30323;
    wire N__30314;
    wire N__30305;
    wire N__30302;
    wire N__30295;
    wire N__30292;
    wire N__30279;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30249;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30237;
    wire N__30236;
    wire N__30235;
    wire N__30234;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30224;
    wire N__30219;
    wire N__30212;
    wire N__30201;
    wire N__30198;
    wire N__30197;
    wire N__30194;
    wire N__30193;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30179;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30149;
    wire N__30148;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30090;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30075;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30060;
    wire N__30057;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30045;
    wire N__30044;
    wire N__30043;
    wire N__30040;
    wire N__30033;
    wire N__30030;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30011;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29998;
    wire N__29993;
    wire N__29992;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29978;
    wire N__29973;
    wire N__29972;
    wire N__29969;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29949;
    wire N__29940;
    wire N__29937;
    wire N__29936;
    wire N__29935;
    wire N__29934;
    wire N__29933;
    wire N__29932;
    wire N__29931;
    wire N__29930;
    wire N__29927;
    wire N__29920;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29895;
    wire N__29892;
    wire N__29883;
    wire N__29882;
    wire N__29881;
    wire N__29880;
    wire N__29879;
    wire N__29878;
    wire N__29877;
    wire N__29876;
    wire N__29871;
    wire N__29868;
    wire N__29863;
    wire N__29856;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29549;
    wire N__29548;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29524;
    wire N__29521;
    wire N__29514;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29396;
    wire N__29391;
    wire N__29388;
    wire N__29387;
    wire N__29384;
    wire N__29383;
    wire N__29380;
    wire N__29379;
    wire N__29376;
    wire N__29369;
    wire N__29364;
    wire N__29363;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29351;
    wire N__29348;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29292;
    wire N__29289;
    wire N__29288;
    wire N__29287;
    wire N__29286;
    wire N__29283;
    wire N__29276;
    wire N__29271;
    wire N__29268;
    wire N__29267;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29255;
    wire N__29254;
    wire N__29253;
    wire N__29252;
    wire N__29251;
    wire N__29250;
    wire N__29243;
    wire N__29234;
    wire N__29229;
    wire N__29228;
    wire N__29227;
    wire N__29224;
    wire N__29223;
    wire N__29222;
    wire N__29219;
    wire N__29218;
    wire N__29211;
    wire N__29204;
    wire N__29199;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29136;
    wire N__29135;
    wire N__29134;
    wire N__29131;
    wire N__29126;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29110;
    wire N__29109;
    wire N__29108;
    wire N__29101;
    wire N__29096;
    wire N__29091;
    wire N__29088;
    wire N__29087;
    wire N__29086;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29072;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29036;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28968;
    wire N__28967;
    wire N__28962;
    wire N__28961;
    wire N__28960;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28942;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28918;
    wire N__28911;
    wire N__28910;
    wire N__28907;
    wire N__28906;
    wire N__28905;
    wire N__28904;
    wire N__28903;
    wire N__28902;
    wire N__28901;
    wire N__28900;
    wire N__28899;
    wire N__28896;
    wire N__28891;
    wire N__28888;
    wire N__28881;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28862;
    wire N__28855;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28838;
    wire N__28837;
    wire N__28836;
    wire N__28835;
    wire N__28834;
    wire N__28833;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28825;
    wire N__28824;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28808;
    wire N__28799;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28779;
    wire N__28778;
    wire N__28775;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28731;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28719;
    wire N__28716;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28708;
    wire N__28703;
    wire N__28700;
    wire N__28699;
    wire N__28694;
    wire N__28691;
    wire N__28686;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28633;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28568;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28415;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28391;
    wire N__28390;
    wire N__28389;
    wire N__28388;
    wire N__28383;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28361;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28349;
    wire N__28348;
    wire N__28341;
    wire N__28338;
    wire N__28337;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28301;
    wire N__28300;
    wire N__28297;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28281;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28273;
    wire N__28270;
    wire N__28265;
    wire N__28260;
    wire N__28257;
    wire N__28256;
    wire N__28253;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28226;
    wire N__28225;
    wire N__28222;
    wire N__28217;
    wire N__28214;
    wire N__28211;
    wire N__28206;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28198;
    wire N__28195;
    wire N__28190;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28178;
    wire N__28177;
    wire N__28174;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28152;
    wire N__28151;
    wire N__28150;
    wire N__28149;
    wire N__28148;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28130;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28118;
    wire N__28115;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28103;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28058;
    wire N__28055;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28043;
    wire N__28040;
    wire N__28039;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28014;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28006;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27987;
    wire N__27984;
    wire N__27983;
    wire N__27980;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27909;
    wire N__27906;
    wire N__27905;
    wire N__27904;
    wire N__27901;
    wire N__27900;
    wire N__27897;
    wire N__27896;
    wire N__27895;
    wire N__27888;
    wire N__27883;
    wire N__27880;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27866;
    wire N__27865;
    wire N__27862;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27840;
    wire N__27837;
    wire N__27836;
    wire N__27835;
    wire N__27832;
    wire N__27827;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27815;
    wire N__27814;
    wire N__27811;
    wire N__27806;
    wire N__27801;
    wire N__27798;
    wire N__27797;
    wire N__27796;
    wire N__27793;
    wire N__27788;
    wire N__27783;
    wire N__27782;
    wire N__27781;
    wire N__27778;
    wire N__27773;
    wire N__27768;
    wire N__27767;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27735;
    wire N__27734;
    wire N__27733;
    wire N__27728;
    wire N__27725;
    wire N__27720;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27677;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27647;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27630;
    wire N__27629;
    wire N__27628;
    wire N__27625;
    wire N__27620;
    wire N__27615;
    wire N__27614;
    wire N__27613;
    wire N__27612;
    wire N__27611;
    wire N__27610;
    wire N__27609;
    wire N__27608;
    wire N__27607;
    wire N__27606;
    wire N__27605;
    wire N__27604;
    wire N__27603;
    wire N__27602;
    wire N__27601;
    wire N__27600;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27596;
    wire N__27595;
    wire N__27594;
    wire N__27593;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27528;
    wire N__27525;
    wire N__27524;
    wire N__27523;
    wire N__27522;
    wire N__27517;
    wire N__27512;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27497;
    wire N__27492;
    wire N__27489;
    wire N__27488;
    wire N__27485;
    wire N__27484;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27426;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27414;
    wire N__27413;
    wire N__27412;
    wire N__27411;
    wire N__27410;
    wire N__27409;
    wire N__27396;
    wire N__27395;
    wire N__27394;
    wire N__27393;
    wire N__27390;
    wire N__27383;
    wire N__27378;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27366;
    wire N__27363;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27261;
    wire N__27260;
    wire N__27255;
    wire N__27252;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27204;
    wire N__27201;
    wire N__27200;
    wire N__27199;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27170;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27155;
    wire N__27150;
    wire N__27147;
    wire N__27146;
    wire N__27145;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27117;
    wire N__27114;
    wire N__27107;
    wire N__27102;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27087;
    wire N__27086;
    wire N__27083;
    wire N__27082;
    wire N__27081;
    wire N__27080;
    wire N__27079;
    wire N__27076;
    wire N__27069;
    wire N__27064;
    wire N__27057;
    wire N__27054;
    wire N__27053;
    wire N__27052;
    wire N__27051;
    wire N__27050;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27034;
    wire N__27031;
    wire N__27026;
    wire N__27023;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26988;
    wire N__26987;
    wire N__26984;
    wire N__26979;
    wire N__26976;
    wire N__26975;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26952;
    wire N__26951;
    wire N__26950;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26921;
    wire N__26916;
    wire N__26913;
    wire N__26912;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26864;
    wire N__26863;
    wire N__26860;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26814;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26787;
    wire N__26786;
    wire N__26781;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26759;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26747;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26733;
    wire N__26732;
    wire N__26731;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26708;
    wire N__26703;
    wire N__26700;
    wire N__26699;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26678;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26634;
    wire N__26631;
    wire N__26630;
    wire N__26625;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26581;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26565;
    wire N__26562;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26525;
    wire N__26524;
    wire N__26521;
    wire N__26516;
    wire N__26511;
    wire N__26508;
    wire N__26507;
    wire N__26502;
    wire N__26499;
    wire N__26498;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26481;
    wire N__26480;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26462;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26405;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26387;
    wire N__26386;
    wire N__26383;
    wire N__26378;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26313;
    wire N__26310;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26286;
    wire N__26283;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26271;
    wire N__26270;
    wire N__26269;
    wire N__26266;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26169;
    wire N__26168;
    wire N__26167;
    wire N__26164;
    wire N__26159;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26145;
    wire N__26144;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26132;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26108;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26055;
    wire N__26052;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26040;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26028;
    wire N__26025;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26013;
    wire N__26010;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__25998;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25923;
    wire N__25922;
    wire N__25919;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25899;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25869;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25847;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25796;
    wire N__25793;
    wire N__25792;
    wire N__25789;
    wire N__25788;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25741;
    wire N__25736;
    wire N__25731;
    wire N__25728;
    wire N__25727;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25707;
    wire N__25706;
    wire N__25705;
    wire N__25702;
    wire N__25697;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25647;
    wire N__25644;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25575;
    wire N__25574;
    wire N__25569;
    wire N__25566;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25061;
    wire N__25060;
    wire N__25057;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25028;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24881;
    wire N__24880;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24830;
    wire N__24829;
    wire N__24826;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24770;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24662;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24627;
    wire N__24626;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24609;
    wire N__24608;
    wire N__24605;
    wire N__24604;
    wire N__24601;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24557;
    wire N__24552;
    wire N__24549;
    wire N__24548;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24524;
    wire N__24523;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24506;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24461;
    wire N__24460;
    wire N__24459;
    wire N__24458;
    wire N__24457;
    wire N__24456;
    wire N__24455;
    wire N__24454;
    wire N__24453;
    wire N__24452;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24448;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24392;
    wire N__24391;
    wire N__24390;
    wire N__24389;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24350;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24326;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24275;
    wire N__24272;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24206;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24152;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24119;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24066;
    wire N__24063;
    wire N__24062;
    wire N__24059;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23909;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23874;
    wire N__23871;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23849;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23814;
    wire N__23811;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23796;
    wire N__23795;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23751;
    wire N__23748;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23733;
    wire N__23732;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23669;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23606;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23543;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23492;
    wire N__23487;
    wire N__23484;
    wire N__23483;
    wire N__23478;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23468;
    wire N__23463;
    wire N__23460;
    wire N__23459;
    wire N__23458;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23422;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23387;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23338;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23297;
    wire N__23292;
    wire N__23289;
    wire N__23288;
    wire N__23287;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23264;
    wire N__23259;
    wire N__23256;
    wire N__23255;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23228;
    wire N__23225;
    wire N__23224;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23212;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23195;
    wire N__23194;
    wire N__23193;
    wire N__23192;
    wire N__23191;
    wire N__23186;
    wire N__23181;
    wire N__23176;
    wire N__23173;
    wire N__23166;
    wire N__23163;
    wire N__23162;
    wire N__23161;
    wire N__23160;
    wire N__23157;
    wire N__23156;
    wire N__23153;
    wire N__23152;
    wire N__23147;
    wire N__23142;
    wire N__23137;
    wire N__23130;
    wire N__23127;
    wire N__23126;
    wire N__23121;
    wire N__23120;
    wire N__23119;
    wire N__23118;
    wire N__23115;
    wire N__23108;
    wire N__23107;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23095;
    wire N__23092;
    wire N__23087;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23046;
    wire N__23043;
    wire N__23042;
    wire N__23037;
    wire N__23034;
    wire N__23033;
    wire N__23032;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22992;
    wire N__22991;
    wire N__22986;
    wire N__22983;
    wire N__22982;
    wire N__22977;
    wire N__22974;
    wire N__22973;
    wire N__22972;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22955;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22943;
    wire N__22942;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22919;
    wire N__22918;
    wire N__22917;
    wire N__22914;
    wire N__22913;
    wire N__22908;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22889;
    wire N__22884;
    wire N__22883;
    wire N__22880;
    wire N__22879;
    wire N__22878;
    wire N__22875;
    wire N__22874;
    wire N__22871;
    wire N__22866;
    wire N__22861;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22847;
    wire N__22846;
    wire N__22845;
    wire N__22844;
    wire N__22843;
    wire N__22840;
    wire N__22835;
    wire N__22828;
    wire N__22825;
    wire N__22820;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22793;
    wire N__22788;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22773;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22616;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22598;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22397;
    wire N__22396;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire \Pc2drone_pll_inst.clk_system_pll ;
    wire GNDG0;
    wire VCCG0;
    wire \pid_alt.O_3_10 ;
    wire \pid_alt.O_3_5 ;
    wire \pid_alt.O_3_14 ;
    wire \pid_alt.O_3_15 ;
    wire \pid_alt.O_3_16 ;
    wire \pid_alt.O_3_17 ;
    wire \pid_alt.O_3_18 ;
    wire \pid_alt.O_3_19 ;
    wire \pid_alt.O_3_20 ;
    wire \pid_alt.O_3_21 ;
    wire \pid_alt.O_3_22 ;
    wire \pid_alt.O_3_23 ;
    wire \pid_alt.O_3_6 ;
    wire \pid_alt.O_3_24 ;
    wire \pid_alt.O_3_7 ;
    wire \pid_alt.O_3_9 ;
    wire alt_kd_7;
    wire alt_kd_2;
    wire alt_kd_1;
    wire alt_kd_5;
    wire alt_ki_6;
    wire alt_ki_7;
    wire alt_ki_1;
    wire alt_ki_3;
    wire alt_ki_4;
    wire alt_ki_5;
    wire \pid_alt.O_4_9 ;
    wire \pid_alt.O_4_24 ;
    wire \pid_alt.O_4_23 ;
    wire \pid_alt.O_4_22 ;
    wire \pid_alt.O_4_10 ;
    wire \pid_alt.O_4_14 ;
    wire \pid_alt.O_4_11 ;
    wire \pid_alt.O_4_17 ;
    wire \pid_alt.O_4_16 ;
    wire \pid_alt.O_4_20 ;
    wire \pid_alt.O_4_18 ;
    wire \pid_alt.O_4_19 ;
    wire \pid_alt.O_4_6 ;
    wire \pid_alt.O_4_21 ;
    wire \pid_alt.O_4_13 ;
    wire \pid_alt.O_4_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_ ;
    wire \pid_alt.N_1666_i_1 ;
    wire \pid_alt.N_3_1 ;
    wire \pid_alt.N_1668_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ;
    wire \pid_alt.N_1674_0_cascade_ ;
    wire \pid_alt.N_1666_i_0 ;
    wire \pid_alt.N_3_0 ;
    wire \pid_alt.N_1668_0 ;
    wire \pid_alt.N_5 ;
    wire \pid_alt.N_1672_0 ;
    wire \pid_front.O_0_16 ;
    wire \pid_front.O_0_17 ;
    wire \pid_front.O_0_18 ;
    wire \pid_front.O_0_19 ;
    wire \pid_front.O_0_12 ;
    wire \pid_front.O_0_7 ;
    wire \pid_front.O_0_22 ;
    wire \pid_front.O_0_23 ;
    wire \pid_front.O_0_24 ;
    wire \pid_front.O_0_21 ;
    wire \pid_front.O_0_20 ;
    wire \pid_front.O_0_14 ;
    wire \pid_front.O_0_10 ;
    wire \pid_front.O_0_13 ;
    wire \pid_alt.O_5_6 ;
    wire \pid_alt.O_5_5 ;
    wire \pid_front.O_0_8 ;
    wire \Commands_frame_decoder.source_CH1data8_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8 ;
    wire \pid_alt.O_5_7 ;
    wire \pid_alt.O_5_8 ;
    wire \pid_alt.O_4_8 ;
    wire \pid_alt.O_5_11 ;
    wire \pid_alt.O_5_22 ;
    wire \pid_alt.O_5_15 ;
    wire \pid_alt.O_5_17 ;
    wire \pid_alt.O_5_20 ;
    wire \pid_alt.O_5_18 ;
    wire \pid_alt.O_5_21 ;
    wire \pid_alt.O_5_19 ;
    wire \pid_alt.O_5_14 ;
    wire \pid_alt.O_5_23 ;
    wire \pid_alt.O_5_16 ;
    wire \pid_alt.O_5_12 ;
    wire \pid_alt.O_5_13 ;
    wire \pid_alt.O_5_24 ;
    wire alt_kd_6;
    wire alt_kd_4;
    wire alt_kd_3;
    wire alt_kd_0;
    wire alt_ki_0;
    wire alt_ki_2;
    wire \Commands_frame_decoder.state_RNIQRI31Z0Z_10 ;
    wire \pid_alt.g0_4_0 ;
    wire \Commands_frame_decoder.stateZ0Z_3 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ;
    wire \pid_alt.O_4_5 ;
    wire \pid_alt.O_3_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ;
    wire \pid_alt.error_d_reg_prevZ0Z_5 ;
    wire \pid_alt.error_d_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prevZ0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_6 ;
    wire \pid_alt.error_p_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prevZ0Z_2 ;
    wire \pid_alt.error_d_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_ ;
    wire \pid_alt.O_5_4 ;
    wire \pid_alt.error_p_regZ0Z_0 ;
    wire \pid_alt.N_1666_i ;
    wire \pid_alt.error_p_regZ0Z_1 ;
    wire \pid_alt.error_d_reg_prevZ0Z_1 ;
    wire \pid_alt.N_1666_i_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_axb_2_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prevZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prevZ0Z_12 ;
    wire \pid_alt.error_p_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ;
    wire \pid_alt.error_p_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prevZ0Z_18 ;
    wire \pid_alt.error_d_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ;
    wire bfn_2_19_0_;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire alt_command_0;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire alt_command_1;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire alt_command_2;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire alt_command_3;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire alt_command_4;
    wire \pid_alt.error_8 ;
    wire bfn_2_20_0_;
    wire alt_command_5;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire alt_command_6;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire alt_command_7;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire alt_kp_1;
    wire drone_altitude_i_10;
    wire alt_kp_0;
    wire alt_kp_6;
    wire \pid_alt.O_5_9 ;
    wire \pid_alt.error_p_regZ0Z_5 ;
    wire \pid_alt.O_5_10 ;
    wire \pid_alt.error_p_regZ0Z_6 ;
    wire alt_kp_7;
    wire alt_kp_3;
    wire \pid_alt.O_3_8 ;
    wire \Commands_frame_decoder.state_RNIRSI31Z0Z_11 ;
    wire \pid_alt.O_3_11 ;
    wire \pid_alt.O_3_12 ;
    wire \pid_alt.O_3_13 ;
    wire \pid_alt.O_4_4 ;
    wire \pid_alt.O_4_7 ;
    wire \pid_alt.O_4_15 ;
    wire \pid_alt.N_664_0_g ;
    wire \Commands_frame_decoder.source_CH1data8lt7_0 ;
    wire \pid_alt.error_d_regZ0Z_0 ;
    wire \pid_alt.error_p_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prevZ0Z_3 ;
    wire \pid_alt.error_d_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ;
    wire \pid_alt.error_p_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prevZ0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ;
    wire bfn_3_14_0_;
    wire \pid_alt.error_i_regZ0Z_1 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_alt.error_i_regZ0Z_2 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_alt.error_i_regZ0Z_3 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_alt.error_i_regZ0Z_4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_alt.error_i_regZ0Z_5 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_alt.error_i_regZ0Z_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_alt.error_i_regZ0Z_7 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_alt.error_i_regZ0Z_8 ;
    wire bfn_3_15_0_;
    wire \pid_alt.error_i_regZ0Z_9 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_alt.error_i_regZ0Z_10 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_alt.error_i_regZ0Z_11 ;
    wire \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_alt.error_i_regZ0Z_12 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_alt.error_i_regZ0Z_13 ;
    wire \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_alt.error_i_regZ0Z_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_alt.error_i_regZ0Z_15 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_alt.error_i_regZ0Z_16 ;
    wire bfn_3_16_0_;
    wire \pid_alt.error_i_regZ0Z_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_alt.error_i_regZ0Z_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_alt.error_i_regZ0Z_19 ;
    wire \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_alt.error_i_regZ0Z_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ;
    wire \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ;
    wire bfn_3_17_0_;
    wire \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ;
    wire \pid_alt.un1_pid_prereg_0 ;
    wire \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1 ;
    wire \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_2 ;
    wire \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_5 ;
    wire \pid_alt.un1_pid_prereg_0_cry_6 ;
    wire bfn_3_18_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_7 ;
    wire \pid_alt.un1_pid_prereg_0_cry_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ;
    wire \pid_alt.un1_pid_prereg_0_cry_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ;
    wire \pid_alt.un1_pid_prereg_0_cry_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ;
    wire \pid_alt.un1_pid_prereg_0_cry_12 ;
    wire \pid_alt.un1_pid_prereg_0_cry_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_14 ;
    wire bfn_3_19_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_15 ;
    wire \pid_alt.un1_pid_prereg_0_cry_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_21 ;
    wire \pid_alt.un1_pid_prereg_0_cry_22 ;
    wire bfn_3_20_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_23 ;
    wire \pid_alt.error_p_regZ0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prevZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ;
    wire \dron_frame_decoder_1.drone_altitude_10 ;
    wire alt_kp_2;
    wire alt_kp_5;
    wire \Commands_frame_decoder.stateZ0Z_2 ;
    wire \pid_alt.error_i_regZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_18 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_19 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_20 ;
    wire \pid_alt.m7_e_4_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_16 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_17 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_14 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_15 ;
    wire \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ;
    wire \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ;
    wire \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ;
    wire \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ;
    wire \pid_alt.error_i_acummZ0Z_3 ;
    wire \pid_alt.error_i_acummZ0Z_1 ;
    wire \pid_alt.N_9_0_cascade_ ;
    wire \pid_alt.N_62_mux_cascade_ ;
    wire \pid_alt.error_i_acummZ0Z_0 ;
    wire \pid_alt.error_i_acummZ0Z_4 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3Z0Z_5 ;
    wire \pid_alt.error_i_acummZ0Z_2 ;
    wire \pid_alt.error_i_acummZ0Z_10 ;
    wire \pid_alt.error_i_acummZ0Z_11 ;
    wire \pid_alt.error_i_acummZ0Z_6 ;
    wire \pid_alt.error_i_acummZ0Z_7 ;
    wire \pid_alt.error_i_acummZ0Z_8 ;
    wire \pid_alt.error_i_acummZ0Z_9 ;
    wire \pid_alt.m35_e_2 ;
    wire \pid_alt.error_i_acummZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ;
    wire \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ;
    wire \pid_alt.error_p_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prevZ0Z_10 ;
    wire \pid_alt.error_d_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ;
    wire drone_altitude_i_11;
    wire \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ;
    wire \pid_alt.error_d_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prevZ0Z_9 ;
    wire \pid_alt.error_p_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prevZ0Z_14 ;
    wire \pid_alt.error_d_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ;
    wire \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_8 ;
    wire \pid_alt.error_p_regZ0Z_8 ;
    wire \pid_alt.error_d_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_7 ;
    wire \pid_alt.error_p_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ;
    wire \pid_alt.error_d_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prevZ0Z_16 ;
    wire \pid_alt.error_p_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ;
    wire \pid_alt.un1_pid_prereg_236_1_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_19 ;
    wire \pid_alt.error_d_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ;
    wire \pid_alt.error_p_regZ0Z_20 ;
    wire \pid_alt.error_d_reg_prevZ0Z_20 ;
    wire \pid_alt.error_d_regZ0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ;
    wire \pid_alt.un1_pid_prereg_236_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ;
    wire \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20 ;
    wire \Commands_frame_decoder.stateZ0Z_11 ;
    wire \Commands_frame_decoder.stateZ0Z_12 ;
    wire \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ;
    wire \Commands_frame_decoder.N_416_cascade_ ;
    wire \Commands_frame_decoder.N_382 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_2_2 ;
    wire \Commands_frame_decoder.N_376_2 ;
    wire \Commands_frame_decoder.N_377 ;
    wire \Commands_frame_decoder.N_376_cascade_ ;
    wire \Commands_frame_decoder.N_379 ;
    wire \Commands_frame_decoder.N_416 ;
    wire \Commands_frame_decoder.N_379_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_1 ;
    wire \Commands_frame_decoder.N_412 ;
    wire \Commands_frame_decoder.stateZ0Z_8 ;
    wire \Commands_frame_decoder.state_RNIF38SZ0Z_6 ;
    wire \Commands_frame_decoder.stateZ0Z_9 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_3 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_2 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_7 ;
    wire \pid_alt.m21_e_0_cascade_ ;
    wire \pid_alt.error_i_acumm7lto4 ;
    wire \pid_alt.m35_e_3 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_9 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_8 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_11 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_6 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_1 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_0 ;
    wire \pid_alt.m21_e_8_cascade_ ;
    wire \pid_alt.error_i_acumm7lto12 ;
    wire \pid_alt.m21_e_2 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ;
    wire \pid_alt.error_i_acumm_preregZ0Z_10 ;
    wire \pid_alt.state_0_g_0 ;
    wire \pid_alt.m21_e_9 ;
    wire \pid_alt.m21_e_10 ;
    wire \pid_alt.N_9_0 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNIO7B05Z0Z_21_cascade_ ;
    wire \pid_alt.un1_reset_1_0_i_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_21 ;
    wire \pid_alt.error_i_acumm7lto13 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14 ;
    wire \pid_alt.error_i_acummZ0Z_13 ;
    wire \pid_alt.N_72_i_0 ;
    wire \pid_alt.un1_reset_1_cascade_ ;
    wire \pid_alt.source_pid_9_0_tz_6_cascade_ ;
    wire \pid_alt.source_pid_9_0_tz_6 ;
    wire \pid_alt.pid_preregZ0Z_2 ;
    wire \pid_alt.pid_preregZ0Z_3 ;
    wire \pid_alt.pid_preregZ0Z_1 ;
    wire \pid_alt.N_44_cascade_ ;
    wire \pid_alt.N_46 ;
    wire \pid_alt.pid_preregZ0Z_0 ;
    wire \pid_alt.N_46_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ;
    wire \pid_alt.pid_preregZ0Z_11 ;
    wire \pid_alt.pid_preregZ0Z_9 ;
    wire \pid_alt.pid_preregZ0Z_10 ;
    wire \pid_alt.pid_preregZ0Z_8 ;
    wire \pid_alt.pid_preregZ0Z_7 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_6 ;
    wire \pid_alt.N_90_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ;
    wire \pid_alt.N_43 ;
    wire \pid_alt.N_48 ;
    wire \pid_alt.pid_preregZ0Z_15 ;
    wire \pid_alt.pid_preregZ0Z_23 ;
    wire \pid_alt.pid_preregZ0Z_21 ;
    wire \pid_alt.pid_preregZ0Z_18 ;
    wire \pid_alt.pid_preregZ0Z_22 ;
    wire \pid_alt.pid_preregZ0Z_20 ;
    wire \pid_alt.pid_preregZ0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_19 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ;
    wire \pid_alt.pid_preregZ0Z_14 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_16 ;
    wire \pid_alt.N_90 ;
    wire \pid_alt.N_305_cascade_ ;
    wire \pid_alt.source_pid_9_0_0_4_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_4 ;
    wire \pid_alt.N_44 ;
    wire \pid_alt.pid_preregZ0Z_5 ;
    wire \pid_alt.pid_preregZ0Z_13 ;
    wire \pid_alt.pid_preregZ0Z_24 ;
    wire \pid_alt.N_305 ;
    wire \pid_alt.pid_preregZ0Z_12 ;
    wire \pid_alt.N_72_i_1 ;
    wire \pid_alt.un1_reset_0_i ;
    wire \pid_alt.error_d_reg_prevZ0Z_17 ;
    wire \pid_alt.error_p_regZ0Z_17 ;
    wire \pid_alt.error_d_regZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ;
    wire bfn_7_7_0_;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1 ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.N_144_1_cascade_ ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.N_126_li_cascade_ ;
    wire \uart_pc.N_143 ;
    wire \uart_pc.N_143_cascade_ ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \Commands_frame_decoder.state_ns_i_a2_0_2_0 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ;
    wire \uart_pc.data_rdyc_1 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.N_378 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire \Commands_frame_decoder.stateZ0Z_0 ;
    wire \Commands_frame_decoder.state_ns_0_i_1_1 ;
    wire \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ;
    wire xy_kp_4;
    wire \Commands_frame_decoder.stateZ0Z_7 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_10 ;
    wire alt_kp_4;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_5 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_6 ;
    wire \Commands_frame_decoder.stateZ0Z_4 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire \pid_front.O_0_6 ;
    wire \pid_front.O_0_4 ;
    wire \pid_front.O_0_9 ;
    wire \pid_front.O_0_15 ;
    wire \dron_frame_decoder_1.drone_altitude_11 ;
    wire drone_altitude_15;
    wire drone_altitude_i_4;
    wire drone_altitude_i_5;
    wire drone_altitude_i_6;
    wire \dron_frame_decoder_1.drone_altitude_9 ;
    wire drone_altitude_i_9;
    wire drone_altitude_i_8;
    wire drone_altitude_i_7;
    wire \pid_alt.drone_altitude_i_0 ;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire uart_input_drone_c;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_8_5_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire bfn_8_6_0_;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire \Commands_frame_decoder.un1_state57_iZ0 ;
    wire \uart_pc.state_srsts_i_0_2_cascade_ ;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.un1_state_4_0_cascade_ ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.N_145_cascade_ ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire \uart_drone.timer_Count_RNO_0_0_1_cascade_ ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \uart_pc.un1_state_2_0 ;
    wire debug_CH2_18A_c;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.CO0_cascade_ ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.un1_state_7_0 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.N_152 ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire xy_kp_6;
    wire xy_kp_5;
    wire drone_altitude_0;
    wire \dron_frame_decoder_1.drone_altitude_4 ;
    wire \dron_frame_decoder_1.drone_altitude_5 ;
    wire \dron_frame_decoder_1.drone_altitude_6 ;
    wire \dron_frame_decoder_1.drone_altitude_7 ;
    wire \dron_frame_decoder_1.drone_altitude_8 ;
    wire drone_altitude_14;
    wire drone_altitude_13;
    wire drone_altitude_12;
    wire \dron_frame_decoder_1.N_513_0 ;
    wire \pid_front.error_p_regZ0Z_9 ;
    wire \pid_front.error_d_reg_prevZ0Z_9 ;
    wire \pid_front.N_1459_i ;
    wire \pid_front.O_0_11 ;
    wire \pid_front.N_1451_i_cascade_ ;
    wire \pid_front.error_d_reg_esr_RNINKUFZ0Z_7_cascade_ ;
    wire \pid_front.un1_pid_prereg_70_0 ;
    wire \pid_front.un1_pid_prereg_23 ;
    wire \pid_front.un1_pid_prereg_23_cascade_ ;
    wire \pid_front.un1_pid_prereg_30_cascade_ ;
    wire \pid_front.error_p_regZ0Z_15 ;
    wire \pid_front.error_d_reg_prevZ0Z_15 ;
    wire \pid_front.un1_pid_prereg_29 ;
    wire \pid_front.un1_pid_prereg_29_cascade_ ;
    wire \pid_front.error_p_regZ0Z_14 ;
    wire \pid_front.un1_pid_prereg_24 ;
    wire \pid_front.state_0_0 ;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire \Commands_frame_decoder.state_0_sqmuxa_1_cascade_ ;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.WDT_RNII19A1Z0Z_4_cascade_ ;
    wire \Commands_frame_decoder.WDT8lto15_N_5L7_1 ;
    wire \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.WDT_RNIAERH3Z0Z_12_cascade_ ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.WDT8_0 ;
    wire \uart_drone.N_126_li_cascade_ ;
    wire \uart_drone.N_143_cascade_ ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire bfn_9_8_0_;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \uart_drone.data_rdyc_1 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.countZ0Z_0 ;
    wire \Commands_frame_decoder.stateZ0Z_14 ;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_13 ;
    wire uart_pc_data_rdy;
    wire \dron_frame_decoder_1.state_ns_0_a3_0_1Z0Z_1_cascade_ ;
    wire \dron_frame_decoder_1.N_220 ;
    wire \dron_frame_decoder_1.N_220_cascade_ ;
    wire \dron_frame_decoder_1.N_224 ;
    wire \dron_frame_decoder_1.N_198_cascade_ ;
    wire \dron_frame_decoder_1.N_200 ;
    wire xy_kp_0;
    wire xy_kp_1;
    wire xy_kp_2;
    wire xy_kp_3;
    wire xy_kp_7;
    wire \Commands_frame_decoder.state_RNIG48SZ0Z_7 ;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_0_0_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ;
    wire \dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ;
    wire \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ;
    wire \dron_frame_decoder_1.drone_H_disp_side_9 ;
    wire drone_altitude_1;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire \pid_front.error_p_regZ0Z_8 ;
    wire \pid_front.error_d_reg_prevZ0Z_8 ;
    wire \pid_front.un1_pid_prereg_80_0 ;
    wire \pid_front.N_1455_i ;
    wire \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11_cascade_ ;
    wire \pid_front.un1_pid_prereg_57_cascade_ ;
    wire \pid_front.un1_pid_prereg_48_cascade_ ;
    wire \pid_front.error_d_reg_prevZ0Z_19 ;
    wire \pid_front.error_p_regZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_56 ;
    wire \pid_front.un1_pid_prereg_56_cascade_ ;
    wire \pid_front.un1_pid_prereg_48 ;
    wire \pid_front.N_1471_i ;
    wire \pid_front.error_p_reg_esr_RNIA93NZ0Z_12 ;
    wire \pid_front.error_d_reg_prevZ0Z_12 ;
    wire \pid_front.error_p_regZ0Z_12 ;
    wire \pid_front.un1_pid_prereg_107_0_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI8NB61Z0Z_11 ;
    wire \uart_drone.N_145_cascade_ ;
    wire \uart_drone.un1_state_4_0_cascade_ ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \reset_module_System.reset6_15_cascade_ ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \reset_module_System.reset6_3_cascade_ ;
    wire \reset_module_System.reset6_13 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire debug_CH0_16A_c;
    wire \uart_drone.un1_state_2_0 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \uart_drone.data_rdyc_1_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire \dron_frame_decoder_1.N_263_5 ;
    wire \dron_frame_decoder_1.N_263_5_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire \dron_frame_decoder_1.N_219_4 ;
    wire \dron_frame_decoder_1.N_219_4_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_1_3 ;
    wire scaler_4_data_5;
    wire \pid_front.O_0_5 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_10 ;
    wire \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13_cascade_ ;
    wire \pid_front.pid_prereg_esr_RNICUKFAZ0Z_6_cascade_ ;
    wire \pid_front.un1_reset_0_i_cascade_ ;
    wire \pid_front.un1_reset_0_i_rn_0 ;
    wire \pid_front.m32_1_cascade_ ;
    wire \pid_front.un1_reset_0_i_sn ;
    wire \pid_alt.error_i_acumm7lto5 ;
    wire \pid_alt.N_62_mux ;
    wire \pid_alt.error_i_acummZ0Z_5 ;
    wire \pid_alt.un1_reset_1_0_i ;
    wire \pid_front.un1_pid_prereg_57 ;
    wire \pid_front.error_p_regZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_18 ;
    wire \pid_front.error_p_regZ0Z_13 ;
    wire \pid_front.error_d_reg_prevZ0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ;
    wire \pid_front.pid_prereg_esr_RNI6FQ75Z0Z_23 ;
    wire \pid_front.un1_pid_prereg_42 ;
    wire \pid_front.un1_pid_prereg_47 ;
    wire \pid_front.un1_pid_prereg_42_cascade_ ;
    wire \pid_front.error_p_regZ0Z_16 ;
    wire \pid_front.error_d_reg_prevZ0Z_16 ;
    wire \pid_front.un1_pid_prereg_35 ;
    wire \pid_front.un1_pid_prereg_36_cascade_ ;
    wire \pid_front.un1_pid_prereg_30 ;
    wire \pid_front.error_p_regZ0Z_17 ;
    wire \pid_front.error_d_reg_prevZ0Z_17 ;
    wire \pid_front.un1_pid_prereg_41 ;
    wire \pid_front.un1_pid_prereg_41_cascade_ ;
    wire \pid_front.un1_pid_prereg_36 ;
    wire \pid_front.error_p_regZ0Z_11 ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.CO0 ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.N_144_1 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire bfn_11_7_0_;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire bfn_11_8_0_;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire bfn_11_9_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.reset6_11 ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_11_10_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire bfn_11_11_0_;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.WDT_RNIIVJ1Z0Z_4_cascade_ ;
    wire \dron_frame_decoder_1.WDT10lt14_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.WDT10lto13_1 ;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \dron_frame_decoder_1.N_218 ;
    wire bfn_11_14_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire throttle_order_5;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_11_15_0_;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire throttle_order_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire throttle_order_10;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire bfn_11_17_0_;
    wire \ppm_encoder_1.un1_aileron_cry_0 ;
    wire \ppm_encoder_1.un1_aileron_cry_1 ;
    wire \ppm_encoder_1.un1_aileron_cry_2 ;
    wire \ppm_encoder_1.un1_aileron_cry_3 ;
    wire \ppm_encoder_1.un1_aileron_cry_4 ;
    wire \ppm_encoder_1.un1_aileron_cry_5 ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire bfn_11_18_0_;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire drone_altitude_2;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire drone_altitude_3;
    wire \dron_frame_decoder_1.N_521_0 ;
    wire \pid_alt.error_d_reg_prevZ0Z_0 ;
    wire \pid_alt.error_d_reg_prev_i_0 ;
    wire \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12_cascade_ ;
    wire \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10_cascade_ ;
    wire \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5_cascade_ ;
    wire \pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5 ;
    wire \pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10 ;
    wire \pid_front.error_p_regZ0Z_7 ;
    wire \pid_front.un1_pid_prereg_60_0_cascade_ ;
    wire \pid_front.N_1447_i_cascade_ ;
    wire \pid_front.error_p_regZ0Z_6 ;
    wire \pid_front.error_d_reg_prevZ0Z_6 ;
    wire \pid_front.un1_pid_prereg_50_0_cascade_ ;
    wire \pid_front.error_d_reg_prevZ0Z_7 ;
    wire \pid_front.m26_e_5_cascade_ ;
    wire \pid_front.m26_e_1_cascade_ ;
    wire \pid_front.m26_e_5 ;
    wire \pid_front.pid_prereg_esr_RNIGSMQ1Z0Z_10 ;
    wire \pid_front.m18_s_5 ;
    wire \pid_front.m18_s_4 ;
    wire \pid_front.m9_e_4_cascade_ ;
    wire \pid_front.m9_e_5 ;
    wire \pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20 ;
    wire \pid_front.pid_prereg_esr_RNIVDO51Z0Z_10 ;
    wire \pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12 ;
    wire \pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13 ;
    wire \pid_front.state_0_1 ;
    wire \pid_front.un1_reset_0_i ;
    wire \pid_front.state_RNIVIRQZ0Z_0_cascade_ ;
    wire \pid_front.error_p_regZ0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNI653NZ0Z_10_cascade_ ;
    wire \pid_front.error_d_reg_prevZ0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11 ;
    wire \pid_front.error_p_reg_esr_RNI653NZ0Z_10 ;
    wire \pid_front.N_1463_i ;
    wire \pid_front.error_p_reg_esr_RNIM6G7Z0Z_9 ;
    wire \uart_drone.N_152 ;
    wire \pid_side.state_0_0 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire bfn_12_12_0_;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire frame_decoder_OFF4data_2;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire frame_decoder_OFF4data_3;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire frame_decoder_OFF4data_4;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire frame_decoder_OFF4data_5;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_OFF4data_6;
    wire frame_decoder_CH4data_6;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire bfn_12_13_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire frame_decoder_OFF4data_7;
    wire frame_decoder_CH4data_7;
    wire \scaler_4.N_1849_i_l_ofxZ0 ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire throttle_order_6;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire throttle_order_3;
    wire throttle_order_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_3_THRU_CO ;
    wire throttle_order_4;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire throttle_order_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire throttle_order_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_1_THRU_CO ;
    wire throttle_order_0;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire throttle_order_7;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ;
    wire \pid_front.error_p_regZ0Z_3 ;
    wire \pid_front.un1_pid_prereg_2_cascade_ ;
    wire \pid_front.un1_pid_prereg_0 ;
    wire \pid_front.un1_pid_prereg_2 ;
    wire \pid_front.un1_pid_prereg_0_cascade_ ;
    wire \pid_front.error_d_reg_prevZ0Z_3 ;
    wire drone_H_disp_front_1;
    wire \dron_frame_decoder_1.N_489_0 ;
    wire bfn_12_21_0_;
    wire \pid_front.un1_pid_prereg_cry_0 ;
    wire \pid_front.pid_preregZ0Z_2 ;
    wire \pid_front.un1_pid_prereg_cry_1 ;
    wire \pid_front.error_p_reg_esr_RNIH7Q01Z0Z_1 ;
    wire \pid_front.pid_preregZ0Z_3 ;
    wire \pid_front.un1_pid_prereg_cry_0_0 ;
    wire \pid_front.error_p_reg_esr_RNIJCSGZ0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNICVO11Z0Z_2 ;
    wire \pid_front.pid_preregZ0Z_4 ;
    wire \pid_front.un1_pid_prereg_cry_1_0 ;
    wire \pid_front.pid_preregZ0Z_5 ;
    wire \pid_front.un1_pid_prereg_cry_2 ;
    wire \pid_front.error_p_reg_esr_RNIH8R01Z0Z_5 ;
    wire \pid_front.pid_preregZ0Z_6 ;
    wire \pid_front.un1_pid_prereg_cry_3 ;
    wire \pid_front.error_d_reg_esr_RNIIFUFZ0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNI94TVZ0Z_6 ;
    wire \pid_front.pid_preregZ0Z_7 ;
    wire \pid_front.un1_pid_prereg_cry_4 ;
    wire \pid_front.un1_pid_prereg_cry_5 ;
    wire \pid_front.error_p_reg_esr_RNIJETVZ0Z_7 ;
    wire \pid_front.error_d_reg_esr_RNINKUFZ0Z_7 ;
    wire \pid_front.pid_preregZ0Z_8 ;
    wire bfn_12_22_0_;
    wire \pid_front.error_d_reg_esr_RNISPUFZ0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNITOTVZ0Z_8 ;
    wire \pid_front.pid_preregZ0Z_9 ;
    wire \pid_front.un1_pid_prereg_cry_6 ;
    wire \pid_front.error_d_reg_esr_RNISPQT1Z0Z_10 ;
    wire \pid_front.error_d_reg_esr_RNI1VUFZ0Z_9 ;
    wire \pid_front.pid_preregZ0Z_10 ;
    wire \pid_front.un1_pid_prereg_cry_7 ;
    wire \pid_front.error_d_reg_esr_RNI9NAB3Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10 ;
    wire \pid_front.pid_preregZ0Z_11 ;
    wire \pid_front.un1_pid_prereg_cry_8 ;
    wire \pid_front.error_p_reg_esr_RNIESET1Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNI1E6A4Z0Z_12 ;
    wire \pid_front.pid_preregZ0Z_12 ;
    wire \pid_front.un1_pid_prereg_cry_9 ;
    wire \pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12 ;
    wire \pid_front.error_d_reg_esr_RNIBO6A4Z0Z_12 ;
    wire \pid_front.pid_preregZ0Z_13 ;
    wire \pid_front.un1_pid_prereg_cry_10 ;
    wire \pid_front.error_p_reg_esr_RNIO6FT1Z0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIN47A4Z0Z_12 ;
    wire \pid_front.pid_preregZ0Z_14 ;
    wire \pid_front.un1_pid_prereg_cry_11 ;
    wire \pid_front.error_p_reg_esr_RNI42GP4Z0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13 ;
    wire \pid_front.pid_preregZ0Z_15 ;
    wire \pid_front.un1_pid_prereg_cry_12 ;
    wire \pid_front.un1_pid_prereg_cry_13 ;
    wire \pid_front.error_p_reg_esr_RNI54OC2Z0Z_14 ;
    wire \pid_front.error_p_reg_esr_RNIGEGP4Z0Z_14 ;
    wire \pid_front.pid_preregZ0Z_16 ;
    wire bfn_12_23_0_;
    wire \pid_front.error_p_reg_esr_RNIBAOC2Z0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNISQGP4Z0Z_15 ;
    wire \pid_front.pid_preregZ0Z_17 ;
    wire \pid_front.un1_pid_prereg_cry_14 ;
    wire \pid_front.error_p_reg_esr_RNIHGOC2Z0Z_16 ;
    wire \pid_front.error_p_reg_esr_RNI87HP4Z0Z_16 ;
    wire \pid_front.pid_preregZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_cry_15 ;
    wire \pid_front.error_p_reg_esr_RNINMOC2Z0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNIKJHP4Z0Z_17 ;
    wire \pid_front.pid_preregZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_cry_16 ;
    wire \pid_front.error_p_reg_esr_RNITSOC2Z0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNI57KP4Z0Z_18 ;
    wire \pid_front.pid_preregZ0Z_20 ;
    wire \pid_front.un1_pid_prereg_cry_17 ;
    wire \pid_front.error_p_reg_esr_RNI8ARC2Z0Z_19 ;
    wire \pid_front.error_p_reg_esr_RNIOUOP4Z0Z_19 ;
    wire \pid_front.pid_preregZ0Z_21 ;
    wire \pid_front.un1_pid_prereg_cry_18 ;
    wire \pid_front.error_p_reg_esr_RNI09RP4Z0Z_20 ;
    wire \pid_front.pid_preregZ0Z_22 ;
    wire \pid_front.un1_pid_prereg_cry_19 ;
    wire \pid_front.un1_pid_prereg_cry_20 ;
    wire \pid_front.pid_preregZ0Z_23 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire \pid_front.un1_pid_prereg_axb_21 ;
    wire front_command_7;
    wire \pid_front.error_p_regZ0Z_20 ;
    wire bfn_13_10_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire bfn_13_11_0_;
    wire bfn_13_12_0_;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire bfn_13_13_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire scaler_4_data_14;
    wire \scaler_4.debug_CH3_20A_c_0 ;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire scaler_4_data_7;
    wire \ppm_encoder_1.N_134_0_cascade_ ;
    wire ppm_output_c;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire throttle_order_2;
    wire scaler_4_data_6;
    wire \ppm_encoder_1.un1_aileron_cry_4_THRU_CO ;
    wire bfn_13_16_0_;
    wire \ppm_encoder_1.un1_elevator_cry_0 ;
    wire front_order_2;
    wire \ppm_encoder_1.un1_elevator_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_1 ;
    wire \ppm_encoder_1.un1_elevator_cry_2 ;
    wire front_order_4;
    wire \ppm_encoder_1.un1_elevator_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_3 ;
    wire front_order_5;
    wire \ppm_encoder_1.un1_elevator_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_4 ;
    wire front_order_6;
    wire \ppm_encoder_1.un1_elevator_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_5 ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire front_order_8;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire bfn_13_17_0_;
    wire front_order_9;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire front_order_10;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire front_order_11;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_13 ;
    wire \ppm_encoder_1.N_299 ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire front_order_13;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_7 ;
    wire \pid_front.error_p_regZ0Z_2 ;
    wire \pid_front.error_d_reg_prevZ0Z_2 ;
    wire \pid_front.error_d_reg_esr_RNIOBP11Z0Z_5 ;
    wire \pid_front.un1_pid_prereg_40_0 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ;
    wire \pid_front.error_p_regZ0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ;
    wire \pid_front.error_d_reg_esr_RNIVOSGZ0Z_5 ;
    wire \pid_front.error_d_reg_prevZ0Z_5 ;
    wire \pid_front.error_p_regZ0Z_4 ;
    wire \pid_front.error_d_reg_prevZ0Z_4 ;
    wire \pid_front.un1_pid_prereg_17 ;
    wire \pid_front.un1_pid_prereg_17_cascade_ ;
    wire \pid_front.un1_pid_prereg_3 ;
    wire \pid_front.error_p_reg_esr_RNIPISGZ0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNI4KF7Z0Z_0_cascade_ ;
    wire \pid_front.error_d_reg_esr_RNINGRVZ0Z_1 ;
    wire \pid_front.error_p_regZ0Z_1 ;
    wire \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1_cascade_ ;
    wire \pid_front.un1_pid_prereg ;
    wire drone_H_disp_front_3;
    wire \pid_front.error_p_reg_esr_RNI6MF7Z0Z_1 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIUQTFZ0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prevZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_5 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_4 ;
    wire \pid_front.error_p_regZ0Z_0 ;
    wire \pid_front.error_d_reg_prevZ0Z_0 ;
    wire \pid_front.N_1427_i ;
    wire \dron_frame_decoder_1.drone_H_disp_front_6 ;
    wire drone_H_disp_front_2;
    wire drone_H_disp_front_0;
    wire \pid_front.error_axb_0 ;
    wire bfn_13_23_0_;
    wire \pid_front.error_axbZ0Z_1 ;
    wire \pid_front.error_1 ;
    wire \pid_front.error_cry_0 ;
    wire \pid_front.error_axbZ0Z_2 ;
    wire \pid_front.error_2 ;
    wire \pid_front.error_cry_1 ;
    wire \pid_front.error_axbZ0Z_3 ;
    wire \pid_front.error_3 ;
    wire \pid_front.error_cry_2 ;
    wire drone_H_disp_front_i_4;
    wire front_command_0;
    wire \pid_front.error_4 ;
    wire \pid_front.error_cry_3 ;
    wire drone_H_disp_front_i_5;
    wire front_command_1;
    wire \pid_front.error_5 ;
    wire \pid_front.error_cry_0_0 ;
    wire drone_H_disp_front_i_6;
    wire front_command_2;
    wire \pid_front.error_6 ;
    wire \pid_front.error_cry_1_0 ;
    wire drone_H_disp_front_i_7;
    wire front_command_3;
    wire \pid_front.error_7 ;
    wire \pid_front.error_cry_2_0 ;
    wire \pid_front.error_cry_3_0 ;
    wire drone_H_disp_front_i_8;
    wire front_command_4;
    wire \pid_front.error_8 ;
    wire bfn_13_24_0_;
    wire front_command_5;
    wire \pid_front.error_9 ;
    wire \pid_front.error_cry_4 ;
    wire drone_H_disp_front_i_10;
    wire front_command_6;
    wire \pid_front.error_10 ;
    wire \pid_front.error_cry_5 ;
    wire \pid_front.error_axbZ0Z_7 ;
    wire \pid_front.error_11 ;
    wire \pid_front.error_cry_6 ;
    wire \pid_front.error_axb_8_l_ofx_0 ;
    wire \pid_front.error_12 ;
    wire \pid_front.error_cry_7 ;
    wire drone_H_disp_front_i_12;
    wire \pid_front.error_13 ;
    wire \pid_front.error_cry_8 ;
    wire drone_H_disp_front_i_13;
    wire \pid_front.error_14 ;
    wire \pid_front.error_cry_9 ;
    wire \pid_front.error_cry_10 ;
    wire \pid_front.error_15 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_10 ;
    wire drone_H_disp_front_11;
    wire drone_H_disp_front_12;
    wire drone_H_disp_front_14;
    wire drone_H_disp_front_15;
    wire \dron_frame_decoder_1.drone_H_disp_front_8 ;
    wire \pid_alt.state_0_0 ;
    wire \pid_alt.state_1_0_0 ;
    wire scaler_4_data_9;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire scaler_4_data_8;
    wire scaler_4_data_10;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire scaler_4_data_13;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \pid_alt.N_72_i ;
    wire \pid_alt.stateZ0Z_0 ;
    wire scaler_4_data_11;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire scaler_4_data_12;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.N_298_cascade_ ;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire front_order_12;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_11 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \ppm_encoder_1.N_297_cascade_ ;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire throttle_order_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_9 ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.N_295 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_6 ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.N_292_cascade_ ;
    wire \ppm_encoder_1.un1_aileron_cry_5_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_7 ;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.N_293_cascade_ ;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire front_order_7;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_8 ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire \ppm_encoder_1.N_294_cascade_ ;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_14 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.N_300_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_10_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_10 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire \ppm_encoder_1.N_296_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire drone_H_disp_front_13;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.N_2150_i ;
    wire bfn_14_23_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire bfn_14_24_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_14_25_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.N_419_g ;
    wire debug_CH3_20A_c;
    wire uart_drone_data_rdy;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.N_313_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_12 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ;
    wire \scaler_4.un2_source_data_0 ;
    wire frame_decoder_OFF4data_0;
    wire frame_decoder_CH4data_0;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire side_order_2;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.N_221_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_4 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_5 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0 ;
    wire \ppm_encoder_1.throttle_m_1 ;
    wire \ppm_encoder_1.N_287_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ;
    wire side_order_1;
    wire \ppm_encoder_1.un1_aileron_cry_0_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_1 ;
    wire \ppm_encoder_1.un1_elevator_cry_0_THRU_CO ;
    wire front_order_1;
    wire \ppm_encoder_1.elevatorZ0Z_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire throttle_order_1;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire bfn_15_17_0_;
    wire \ppm_encoder_1.throttle_RNIUINC6Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.elevator_RNIFISN6Z0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.throttle_RNILVOO6Z0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8 ;
    wire bfn_15_18_0_;
    wire \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.elevator_RNIC22D6Z0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.elevator_RNIH72D6Z0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire bfn_15_19_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_18 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_0 ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire bfn_15_21_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire bfn_15_22_0_;
    wire CONSTANT_ONE_NET;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ;
    wire \ppm_encoder_1.N_232_cascade_ ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire \ppm_encoder_1.N_139_17 ;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ;
    wire \ppm_encoder_1.N_139_17_cascade_ ;
    wire \ppm_encoder_1.N_139 ;
    wire \pid_front.un1_pid_prereg_92 ;
    wire \pid_front.un1_pid_prereg_93 ;
    wire \pid_front.error_p_reg_esr_RNIGKTC2Z0Z_20 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \pid_front.error_d_reg_prevZ0Z_20 ;
    wire side_order_10;
    wire side_order_11;
    wire side_order_6;
    wire side_order_7;
    wire side_order_8;
    wire side_order_9;
    wire side_order_0;
    wire side_order_5;
    wire side_order_4;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ;
    wire \ppm_encoder_1.aileronZ0Z_2 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.N_221 ;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.N_232 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIT3R05Z0Z_3 ;
    wire \ppm_encoder_1.N_289 ;
    wire side_order_3;
    wire \ppm_encoder_1.un1_aileron_cry_2_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_3 ;
    wire \ppm_encoder_1.un1_elevator_cry_2_THRU_CO ;
    wire front_order_3;
    wire \ppm_encoder_1.elevatorZ0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_11_mux ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.N_2150_0 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ;
    wire \pid_front.error_d_reg_prevZ0Z_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \pid_side.m32_1 ;
    wire reset_system;
    wire \pid_side.m26_e_5_cascade_ ;
    wire \pid_side.N_11_0_cascade_ ;
    wire \pid_side.pid_prereg_esr_RNILRSP2Z0Z_5 ;
    wire \pid_side.m26_e_5 ;
    wire \pid_side.pid_prereg_esr_RNIGJDR1Z0Z_10_cascade_ ;
    wire \pid_side.m18_s_4 ;
    wire \pid_side.pid_prereg_esr_RNIQBAH2Z0Z_23_cascade_ ;
    wire \pid_side.un1_reset_0_i_sn ;
    wire \pid_side.i19_mux_cascade_ ;
    wire \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12 ;
    wire \pid_side.N_11_0 ;
    wire \pid_side.pid_prereg_esr_RNIEUA9Z0Z_12_cascade_ ;
    wire \pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10 ;
    wire \pid_side.N_82_mux ;
    wire side_order_12;
    wire \ppm_encoder_1.un2_throttle_iv_0_0 ;
    wire \ppm_encoder_1.init_pulses_2_sqmuxa_0 ;
    wire front_order_0;
    wire pid_altitude_dv;
    wire \ppm_encoder_1.elevatorZ0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_10_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_8 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ;
    wire scaler_4_data_4;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.N_314_cascade_ ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_10 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_11 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.elevatorZ0Z_2 ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.N_288 ;
    wire \ppm_encoder_1.N_290 ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ;
    wire \pid_front.error_d_reg_prevZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_153_d ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \pid_front.error_d_reg_prevZ0Z_11 ;
    wire \pid_alt.state_RNIFCSD1Z0Z_0 ;
    wire \pid_alt.N_664_0 ;
    wire \pid_side.pid_preregZ0Z_0 ;
    wire \pid_side.pid_preregZ0Z_1 ;
    wire debug_CH1_0A_c;
    wire \pid_side.stateZ0Z_0 ;
    wire \pid_side.m18_s_5 ;
    wire \pid_side.stateZ0Z_1 ;
    wire \pid_side.un1_reset_0_i_rn_0 ;
    wire \pid_side.m26_e_1 ;
    wire \pid_side.m9_e_4 ;
    wire \pid_side.m9_e_5_cascade_ ;
    wire \pid_side.pid_prereg_esr_RNIFB07Z0Z_20 ;
    wire \pid_side.pid_prereg_esr_RNIFB07Z0Z_20_cascade_ ;
    wire side_order_13;
    wire \pid_side.state_0_1 ;
    wire \pid_side.un1_reset_0_i ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ;
    wire \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ;
    wire bfn_18_15_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire bfn_18_16_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire bfn_18_17_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12 ;
    wire \ppm_encoder_1.PPM_STATE_53_d ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_5 ;
    wire \pid_front.un1_pid_prereg_axb_0 ;
    wire \pid_front.pid_preregZ0Z_0 ;
    wire \pid_front.error_d_reg_prevZ0Z_18 ;
    wire \pid_front.state_0_g_0 ;
    wire \pid_front.O_6 ;
    wire \pid_front.error_d_regZ0Z_2 ;
    wire GB_BUFFER_reset_system_g_THRU_CO;
    wire bfn_20_9_0_;
    wire \pid_side.un1_pid_prereg_cry_0_THRU_CO ;
    wire \pid_side.un1_pid_prereg_cry_0 ;
    wire \pid_side.pid_preregZ0Z_2 ;
    wire \pid_side.un1_pid_prereg_cry_1 ;
    wire \pid_side.pid_preregZ0Z_3 ;
    wire \pid_side.un1_pid_prereg_cry_0_0 ;
    wire \pid_side.pid_preregZ0Z_4 ;
    wire \pid_side.un1_pid_prereg_cry_1_0 ;
    wire \pid_side.pid_preregZ0Z_5 ;
    wire \pid_side.un1_pid_prereg_cry_2 ;
    wire \pid_side.pid_preregZ0Z_6 ;
    wire \pid_side.un1_pid_prereg_cry_3 ;
    wire \pid_side.pid_preregZ0Z_7 ;
    wire \pid_side.un1_pid_prereg_cry_4 ;
    wire \pid_side.un1_pid_prereg_cry_5 ;
    wire \pid_side.pid_preregZ0Z_8 ;
    wire bfn_20_10_0_;
    wire \pid_side.pid_preregZ0Z_9 ;
    wire \pid_side.un1_pid_prereg_cry_6 ;
    wire \pid_side.pid_preregZ0Z_10 ;
    wire \pid_side.un1_pid_prereg_cry_7 ;
    wire \pid_side.pid_preregZ0Z_11 ;
    wire \pid_side.un1_pid_prereg_cry_8 ;
    wire \pid_side.pid_preregZ0Z_12 ;
    wire \pid_side.un1_pid_prereg_cry_9 ;
    wire \pid_side.pid_preregZ0Z_13 ;
    wire \pid_side.un1_pid_prereg_cry_10 ;
    wire \pid_side.pid_preregZ0Z_14 ;
    wire \pid_side.un1_pid_prereg_cry_11 ;
    wire \pid_side.pid_preregZ0Z_15 ;
    wire \pid_side.un1_pid_prereg_cry_12 ;
    wire \pid_side.un1_pid_prereg_cry_13 ;
    wire \pid_side.pid_preregZ0Z_16 ;
    wire bfn_20_11_0_;
    wire \pid_side.pid_preregZ0Z_17 ;
    wire \pid_side.un1_pid_prereg_cry_14 ;
    wire \pid_side.pid_preregZ0Z_18 ;
    wire \pid_side.un1_pid_prereg_cry_15 ;
    wire \pid_side.pid_preregZ0Z_19 ;
    wire \pid_side.un1_pid_prereg_cry_16 ;
    wire \pid_side.pid_preregZ0Z_20 ;
    wire \pid_side.un1_pid_prereg_cry_17 ;
    wire \pid_side.pid_preregZ0Z_21 ;
    wire \pid_side.un1_pid_prereg_cry_18 ;
    wire \pid_side.pid_preregZ0Z_22 ;
    wire \pid_side.un1_pid_prereg_cry_19 ;
    wire \pid_side.un1_pid_prereg_cry_20 ;
    wire \pid_side.pid_preregZ0Z_23 ;
    wire \pid_side.error_d_reg_prev_esr_RNILHF23Z0Z_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNIJV5H1Z0Z_15 ;
    wire \pid_side.un1_pid_prereg_30_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI0PB23Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNI4UC23Z0Z_17 ;
    wire \pid_side.error_d_reg_prev_esr_RNI5I6H1Z0Z_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNIP56H1Z0Z_16 ;
    wire \pid_side.error_d_reg_prevZ0Z_16 ;
    wire \pid_side.un1_pid_prereg_35 ;
    wire \pid_side.un1_pid_prereg_36_cascade_ ;
    wire \pid_side.un1_pid_prereg_30 ;
    wire \pid_side.error_d_reg_prev_esr_RNIC5C23Z0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNI89K23Z0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNIGJM23Z0Z_20 ;
    wire \pid_side.un1_pid_prereg_axb_21 ;
    wire \ppm_encoder_1.N_286 ;
    wire \ppm_encoder_1.aileronZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNIGV8H1Z0Z_19 ;
    wire drone_H_disp_side_1;
    wire uart_drone_data_2;
    wire drone_H_disp_side_2;
    wire drone_H_disp_side_3;
    wire \dron_frame_decoder_1.N_505_0 ;
    wire drone_H_disp_front_i_9;
    wire uart_drone_data_1;
    wire \dron_frame_decoder_1.drone_H_disp_front_9 ;
    wire \dron_frame_decoder_1.N_481_0 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_4 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_6 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_7 ;
    wire \pid_front.stateZ0Z_1 ;
    wire \pid_front.un1_pid_prereg_cry_0_THRU_CO ;
    wire \pid_front.un1_pid_prereg_axb_1 ;
    wire \pid_front.stateZ0Z_0 ;
    wire \pid_front.pid_preregZ0Z_1 ;
    wire side_command_7;
    wire \pid_front.O_7 ;
    wire \pid_front.error_d_regZ0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNI5QI23Z0Z_5 ;
    wire \pid_side.un1_pid_prereg_axb_1 ;
    wire \pid_side.error_p_reg_esr_RNISH6JZ0Z_0_cascade_ ;
    wire \pid_side.error_d_reg_esr_RNIFP9R2Z0Z_1 ;
    wire \pid_side.N_1546_i ;
    wire \pid_side.error_d_reg_prevZ0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1_cascade_ ;
    wire \pid_side.un1_pid_prereg ;
    wire \pid_side.error_d_reg_prevZ0Z_0 ;
    wire \pid_side.un1_pid_prereg_axb_0 ;
    wire \pid_side.error_p_reg_esr_RNIAVKD1Z0Z_1 ;
    wire \pid_side.un1_pid_prereg_18_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13_cascade_ ;
    wire \pid_side.error_d_reg_prevZ0Z_13 ;
    wire \pid_side.error_d_reg_prev_esr_RNI4NA21Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNIDP5H1Z0Z_14 ;
    wire \pid_side.error_d_reg_esr_RNIKMFP2Z0Z_10 ;
    wire \pid_side.N_1582_i ;
    wire \pid_side.N_1582_i_cascade_ ;
    wire \pid_side.error_d_reg_esr_RNI104E2Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNIKCB23Z0Z_13 ;
    wire \pid_side.un1_pid_prereg_23 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ;
    wire \pid_side.un1_pid_prereg_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNIBAGJ2Z0Z_12 ;
    wire \pid_side.un1_pid_prereg_29 ;
    wire \pid_side.error_d_reg_prev_esr_RNIO9BH1Z0Z_20 ;
    wire \pid_side.error_d_reg_prev_esr_RNILJFJ2Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQCA21Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12 ;
    wire \pid_side.N_1590_i_cascade_ ;
    wire \pid_side.error_d_reg_esr_RNIVTFJ2Z0Z_12 ;
    wire \pid_side.un1_pid_prereg_107_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11 ;
    wire \pid_side.error_d_reg_prevZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2VN9Z0Z_12 ;
    wire \pid_side.error_d_reg_prevZ0Z_11 ;
    wire \pid_side.O_2_15 ;
    wire \pid_side.error_p_regZ0Z_11 ;
    wire \ppm_encoder_1.N_291 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ;
    wire \pid_side.un1_pid_prereg_56 ;
    wire \pid_side.error_d_reg_prevZ0Z_19 ;
    wire \pid_side.un1_pid_prereg_57 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire drone_H_disp_side_0;
    wire \pid_side.error_axb_0 ;
    wire bfn_21_17_0_;
    wire \pid_side.error_axbZ0Z_1 ;
    wire \pid_side.error_1 ;
    wire \pid_side.error_cry_0 ;
    wire \pid_side.error_axbZ0Z_2 ;
    wire \pid_side.error_2 ;
    wire \pid_side.error_cry_1 ;
    wire \pid_side.error_axbZ0Z_3 ;
    wire \pid_side.error_3 ;
    wire \pid_side.error_cry_2 ;
    wire drone_H_disp_side_i_4;
    wire side_command_0;
    wire \pid_side.error_4 ;
    wire \pid_side.error_cry_3 ;
    wire drone_H_disp_side_i_5;
    wire side_command_1;
    wire \pid_side.error_5 ;
    wire \pid_side.error_cry_0_0 ;
    wire drone_H_disp_side_i_6;
    wire side_command_2;
    wire \pid_side.error_6 ;
    wire \pid_side.error_cry_1_0 ;
    wire drone_H_disp_side_i_7;
    wire side_command_3;
    wire \pid_side.error_7 ;
    wire \pid_side.error_cry_2_0 ;
    wire \pid_side.error_cry_3_0 ;
    wire drone_H_disp_side_i_8;
    wire side_command_4;
    wire \pid_side.error_8 ;
    wire bfn_21_18_0_;
    wire drone_H_disp_side_i_9;
    wire side_command_5;
    wire \pid_side.error_9 ;
    wire \pid_side.error_cry_4 ;
    wire drone_H_disp_side_i_10;
    wire side_command_6;
    wire \pid_side.error_10 ;
    wire \pid_side.error_cry_5 ;
    wire \pid_side.error_axbZ0Z_7 ;
    wire \pid_side.error_11 ;
    wire \pid_side.error_cry_6 ;
    wire \pid_side.error_axb_8_l_ofxZ0 ;
    wire \pid_side.error_12 ;
    wire \pid_side.error_cry_7 ;
    wire drone_H_disp_side_i_12;
    wire \pid_side.error_13 ;
    wire \pid_side.error_cry_8 ;
    wire drone_H_disp_side_i_13;
    wire \pid_side.error_14 ;
    wire \pid_side.error_cry_9 ;
    wire \pid_side.error_cry_10 ;
    wire \pid_side.error_15 ;
    wire uart_drone_data_3;
    wire drone_H_disp_side_11;
    wire uart_drone_data_4;
    wire drone_H_disp_side_12;
    wire uart_drone_data_5;
    wire drone_H_disp_side_13;
    wire uart_drone_data_7;
    wire drone_H_disp_side_15;
    wire uart_drone_data_0;
    wire \dron_frame_decoder_1.drone_H_disp_side_8 ;
    wire \pid_front.O_10 ;
    wire \pid_front.error_d_regZ0Z_6 ;
    wire \pid_side.error_d_reg_esr_RNI76TK1Z0Z_5 ;
    wire \pid_side.un1_pid_prereg_40_0_cascade_ ;
    wire \pid_side.error_d_reg_esr_RNI86Q93Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ;
    wire \pid_side.un1_pid_prereg_17_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNI10TK1Z0Z_3 ;
    wire \pid_side.error_d_reg_prevZ0Z_4 ;
    wire \pid_side.un1_pid_prereg_17 ;
    wire \pid_side.error_p_reg_esr_RNISPP93Z0Z_2 ;
    wire \pid_side.O_2_9 ;
    wire \pid_side.O_2_4 ;
    wire \pid_side.error_p_regZ0Z_0 ;
    wire \pid_side.state_RNINK4UZ0Z_0 ;
    wire \pid_side.error_p_reg_esr_RNIE47JZ0Z_9 ;
    wire \pid_side.error_d_reg_prevZ0Z_15 ;
    wire \pid_side.un1_pid_prereg_24 ;
    wire \pid_side.un1_pid_prereg_48 ;
    wire \pid_side.un1_pid_prereg_36 ;
    wire \pid_side.error_d_reg_prev_esr_RNIOHC23Z0Z_16 ;
    wire \pid_side.error_d_reg_prevZ0Z_18 ;
    wire \pid_side.un1_pid_prereg_47 ;
    wire \pid_side.un1_pid_prereg_47_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIVB6H1Z0Z_17 ;
    wire \pid_side.error_d_reg_prevZ0Z_10 ;
    wire \pid_side.O_1_4 ;
    wire \pid_side.error_d_regZ0Z_0 ;
    wire \pid_side.O_1_8 ;
    wire \pid_side.error_d_regZ0Z_4 ;
    wire \pid_side.O_1_5 ;
    wire \pid_side.error_d_regZ0Z_1 ;
    wire uart_pc_data_4;
    wire xy_kd_4;
    wire uart_drone_data_6;
    wire drone_H_disp_side_14;
    wire \dron_frame_decoder_1.N_497_0 ;
    wire \pid_front.O_9 ;
    wire \pid_front.error_d_regZ0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNI5PH23Z0Z_1 ;
    wire \pid_side.un1_pid_prereg_2 ;
    wire \pid_side.un1_pid_prereg_2_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIRPSK1Z0Z_2 ;
    wire \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ;
    wire \pid_side.un1_pid_prereg_0 ;
    wire \pid_side.error_d_reg_prevZ0Z_3 ;
    wire \pid_side.un1_pid_prereg_3 ;
    wire \pid_side.error_d_reg_prevZ0Z_2 ;
    wire \pid_side.error_d_reg_prevZ0Z_14 ;
    wire \pid_side.error_p_regZ0Z_5 ;
    wire \pid_side.error_d_reg_prevZ0Z_5 ;
    wire \pid_side.N_1566_i_cascade_ ;
    wire \pid_side.N_1578_i_cascade_ ;
    wire \pid_side.error_d_reg_esr_RNID3MD1Z0Z_9 ;
    wire \pid_side.N_1574_i_cascade_ ;
    wire \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8 ;
    wire \pid_side.un1_pid_prereg_80_0 ;
    wire \pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIL1CR2Z0Z_8 ;
    wire \pid_side.error_d_reg_prevZ0Z_8 ;
    wire \pid_side.error_d_reg_prevZ0Z_9 ;
    wire \pid_side.un1_pid_prereg_41 ;
    wire \pid_side.un1_pid_prereg_42 ;
    wire \pid_side.error_d_reg_prevZ0Z_17 ;
    wire \pid_side.O_1_13 ;
    wire \pid_side.error_d_regZ0Z_9 ;
    wire \pid_side.un1_pid_prereg_93 ;
    wire \pid_side.un1_pid_prereg_92 ;
    wire \pid_front.O_12 ;
    wire \pid_front.error_d_regZ0Z_8 ;
    wire \pid_front.O_16 ;
    wire \pid_front.error_d_regZ0Z_12 ;
    wire \pid_front.O_14 ;
    wire \pid_front.error_d_regZ0Z_10 ;
    wire \pid_side.O_2_8 ;
    wire \pid_side.error_p_regZ0Z_4 ;
    wire \pid_side.O_2_5 ;
    wire \pid_side.error_p_regZ0Z_1 ;
    wire \pid_side.O_2_7 ;
    wire \pid_side.error_p_regZ0Z_3 ;
    wire \pid_side.O_2_22 ;
    wire \pid_side.error_p_regZ0Z_18 ;
    wire \pid_side.O_2_6 ;
    wire \pid_side.error_p_regZ0Z_2 ;
    wire \pid_side.O_2_20 ;
    wire \pid_side.error_p_regZ0Z_16 ;
    wire \pid_side.O_2_21 ;
    wire \pid_side.error_p_regZ0Z_17 ;
    wire \pid_side.O_1_6 ;
    wire \pid_side.error_d_regZ0Z_2 ;
    wire \pid_side.O_2_17 ;
    wire \pid_side.error_p_regZ0Z_13 ;
    wire \pid_side.O_2_12 ;
    wire \pid_side.error_p_regZ0Z_8 ;
    wire \pid_side.O_2_24 ;
    wire \pid_side.error_p_regZ0Z_20 ;
    wire \pid_side.O_2_18 ;
    wire \pid_side.error_p_regZ0Z_14 ;
    wire \pid_side.O_2_14 ;
    wire \pid_side.error_p_regZ0Z_10 ;
    wire \pid_side.O_2_19 ;
    wire \pid_side.error_p_regZ0Z_15 ;
    wire \pid_side.O_2_10 ;
    wire \pid_side.O_2_13 ;
    wire \pid_side.error_p_regZ0Z_9 ;
    wire \pid_side.O_2_11 ;
    wire \pid_side.O_2_23 ;
    wire \pid_side.error_p_regZ0Z_19 ;
    wire \pid_side.O_2_16 ;
    wire \pid_side.error_p_regZ0Z_12 ;
    wire \pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6 ;
    wire \pid_side.un1_pid_prereg_60_0_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNI1DBR2Z0Z_6 ;
    wire \pid_side.N_1570_i_cascade_ ;
    wire \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7 ;
    wire \pid_side.un1_pid_prereg_70_0 ;
    wire \pid_side.error_p_regZ0Z_7 ;
    wire \pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7_cascade_ ;
    wire \pid_side.error_d_reg_prevZ0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNIBNBR2Z0Z_7 ;
    wire \pid_side.error_p_regZ0Z_6 ;
    wire \pid_side.error_d_reg_prevZ0Z_6 ;
    wire \pid_side.un1_pid_prereg_50_0 ;
    wire \pid_side.O_1_15 ;
    wire \pid_side.error_d_regZ0Z_11 ;
    wire \pid_side.O_1_21 ;
    wire \pid_side.error_d_regZ0Z_17 ;
    wire \pid_side.O_1_19 ;
    wire \pid_side.error_d_regZ0Z_15 ;
    wire \pid_side.O_1_12 ;
    wire \pid_side.error_d_regZ0Z_8 ;
    wire \pid_side.O_1_9 ;
    wire \pid_side.error_d_regZ0Z_5 ;
    wire \pid_side.O_1_16 ;
    wire \pid_side.error_d_regZ0Z_12 ;
    wire \pid_side.O_1_18 ;
    wire \pid_side.error_d_regZ0Z_14 ;
    wire \pid_side.O_1_7 ;
    wire \pid_side.error_d_regZ0Z_3 ;
    wire \pid_side.O_1_17 ;
    wire \pid_side.error_d_regZ0Z_13 ;
    wire \pid_side.O_1_14 ;
    wire \pid_side.error_d_regZ0Z_10 ;
    wire \pid_side.O_1_23 ;
    wire \pid_side.error_d_regZ0Z_19 ;
    wire \pid_side.O_1_24 ;
    wire \pid_side.O_1_10 ;
    wire \pid_side.error_d_regZ0Z_6 ;
    wire \pid_side.O_1_22 ;
    wire \pid_side.error_d_regZ0Z_18 ;
    wire \pid_side.O_1_11 ;
    wire \pid_side.error_d_regZ0Z_7 ;
    wire \pid_side.O_1_20 ;
    wire \pid_side.error_d_regZ0Z_16 ;
    wire \pid_side.N_599_0 ;
    wire uart_pc_data_0;
    wire xy_kd_0;
    wire uart_pc_data_1;
    wire xy_kd_1;
    wire uart_pc_data_2;
    wire xy_kd_2;
    wire uart_pc_data_5;
    wire xy_kd_5;
    wire uart_pc_data_6;
    wire xy_kd_6;
    wire uart_pc_data_7;
    wire xy_kd_7;
    wire uart_pc_data_3;
    wire xy_kd_3;
    wire \Commands_frame_decoder.state_RNITUI31Z0Z_13 ;
    wire \pid_side.error_d_regZ0Z_20 ;
    wire \pid_side.error_d_reg_prevZ0Z_20 ;
    wire \pid_side.state_0_g_0 ;
    wire reset_system_g;
    wire \pid_front.O_4 ;
    wire \pid_front.error_d_regZ0Z_0 ;
    wire \pid_front.O_5 ;
    wire \pid_front.error_d_regZ0Z_1 ;
    wire \pid_front.O_17 ;
    wire \pid_front.error_d_regZ0Z_13 ;
    wire \pid_front.O_15 ;
    wire \pid_front.error_d_regZ0Z_11 ;
    wire \pid_front.O_13 ;
    wire \pid_front.error_d_regZ0Z_9 ;
    wire \pid_front.O_20 ;
    wire \pid_front.error_d_regZ0Z_16 ;
    wire \pid_front.O_21 ;
    wire \pid_front.error_d_regZ0Z_17 ;
    wire \pid_front.O_22 ;
    wire \pid_front.error_d_regZ0Z_18 ;
    wire \pid_front.O_23 ;
    wire \pid_front.error_d_regZ0Z_19 ;
    wire \pid_front.O_24 ;
    wire \pid_front.error_d_regZ0Z_20 ;
    wire \pid_front.O_18 ;
    wire \pid_front.error_d_regZ0Z_14 ;
    wire \pid_front.O_8 ;
    wire \pid_front.error_d_regZ0Z_4 ;
    wire \pid_front.O_11 ;
    wire \pid_front.error_d_regZ0Z_7 ;
    wire \pid_front.O_19 ;
    wire \pid_front.error_d_regZ0Z_15 ;
    wire _gnd_net_;
    wire clk_system_pll_g;
    wire \pid_front.N_543_0 ;
    wire N_665_g;

    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .TEST_MODE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVR=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVQ=3'b110;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVF=7'b0111111;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \Pc2drone_pll_inst.Pc2drone_pll_inst_pll  (
            .PLLOUTGLOBAL(),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__42457),
            .PLLOUTCORE(\Pc2drone_pll_inst.clk_system_pll ),
            .LOCK(),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__59697));
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42363),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42326),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__24010,N__24062,N__24100,N__24152,N__24205,N__23542,N__23605,N__23668,N__23731,N__23794,N__23848,N__23908,N__23338,N__23386,N__23422,N__30685}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__24312,N__23946,N__25680,N__29316,N__24303,N__25692,N__23976,N__23958}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,\pid_alt.O_5_24 ,\pid_alt.O_5_23 ,\pid_alt.O_5_22 ,\pid_alt.O_5_21 ,\pid_alt.O_5_20 ,\pid_alt.O_5_19 ,\pid_alt.O_5_18 ,\pid_alt.O_5_17 ,\pid_alt.O_5_16 ,\pid_alt.O_5_15 ,\pid_alt.O_5_14 ,\pid_alt.O_5_13 ,\pid_alt.O_5_12 ,\pid_alt.O_5_11 ,\pid_alt.O_5_10 ,\pid_alt.O_5_9 ,\pid_alt.O_5_8 ,\pid_alt.O_5_7 ,\pid_alt.O_5_6 ,\pid_alt.O_5_5 ,\pid_alt.O_5_4 ,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50}));
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42230),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42229),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66}),
            .ADDSUBBOT(),
            .A({N__24017,N__24058,N__24107,N__24151,N__24206,N__23543,N__23606,N__23669,N__23732,N__23795,N__23849,N__23909,N__23345,N__23387,N__23429,N__30686}),
            .C({dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82}),
            .B({dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__22083,N__22095,N__22041,N__22050,N__22059,N__22632,N__22071,N__22644}),
            .OHOLDTOP(),
            .O({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,\pid_alt.O_4_24 ,\pid_alt.O_4_23 ,\pid_alt.O_4_22 ,\pid_alt.O_4_21 ,\pid_alt.O_4_20 ,\pid_alt.O_4_19 ,\pid_alt.O_4_18 ,\pid_alt.O_4_17 ,\pid_alt.O_4_16 ,\pid_alt.O_4_15 ,\pid_alt.O_4_14 ,\pid_alt.O_4_13 ,\pid_alt.O_4_12 ,\pid_alt.O_4_11 ,\pid_alt.O_4_10 ,\pid_alt.O_4_9 ,\pid_alt.O_4_8 ,\pid_alt.O_4_7 ,\pid_alt.O_4_6 ,\pid_alt.O_4_5 ,\pid_alt.O_4_4 ,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101}));
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_2_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42287),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42286),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .ADDSUBBOT(),
            .A({N__24021,N__24063,N__24111,N__24159,N__24207,N__23550,N__23610,N__23676,N__23733,N__23796,N__23856,N__23916,N__23352,N__23394,N__23436,N__30693}),
            .C({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133}),
            .B({dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,N__21969,N__22686,N__22101,N__22677,N__22668,N__21963,N__21957,N__22656}),
            .OHOLDTOP(),
            .O({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,\pid_alt.O_3_24 ,\pid_alt.O_3_23 ,\pid_alt.O_3_22 ,\pid_alt.O_3_21 ,\pid_alt.O_3_20 ,\pid_alt.O_3_19 ,\pid_alt.O_3_18 ,\pid_alt.O_3_17 ,\pid_alt.O_3_16 ,\pid_alt.O_3_15 ,\pid_alt.O_3_14 ,\pid_alt.O_3_13 ,\pid_alt.O_3_12 ,\pid_alt.O_3_11 ,\pid_alt.O_3_10 ,\pid_alt.O_3_9 ,\pid_alt.O_3_8 ,\pid_alt.O_3_7 ,\pid_alt.O_3_6 ,\pid_alt.O_3_5 ,\pid_alt.O_3_4 ,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}));
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42288),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42237),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168}),
            .ADDSUBBOT(),
            .A({N__39453,N__39498,N__38960,N__39003,N__39051,N__39099,N__39159,N__39210,N__39270,N__39326,N__38634,N__38691,N__38751,N__38802,N__38853,N__38912}),
            .C({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .B({dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,N__31967,N__30758,N__30722,N__29423,N__32006,N__32033,N__32076,N__32111}),
            .OHOLDTOP(),
            .O({dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,\pid_front.O_0_24 ,\pid_front.O_0_23 ,\pid_front.O_0_22 ,\pid_front.O_0_21 ,\pid_front.O_0_20 ,\pid_front.O_0_19 ,\pid_front.O_0_18 ,\pid_front.O_0_17 ,\pid_front.O_0_16 ,\pid_front.O_0_15 ,\pid_front.O_0_14 ,\pid_front.O_0_13 ,\pid_front.O_0_12 ,\pid_front.O_0_11 ,\pid_front.O_0_10 ,\pid_front.O_0_9 ,\pid_front.O_0_8 ,\pid_front.O_0_7 ,\pid_front.O_0_6 ,\pid_front.O_0_5 ,\pid_front.O_0_4 ,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203}));
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42458),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42432),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .ADDSUBBOT(),
            .A({N__52736,N__52769,N__51869,N__51905,N__51941,N__51977,N__52028,N__52082,N__52127,N__52166,N__51575,N__51620,N__51665,N__51704,N__51740,N__51779}),
            .C({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235}),
            .B({dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,N__55388,N__55595,N__55766,N__53249,N__55223,N__55943,N__56153,N__56324}),
            .OHOLDTOP(),
            .O({dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,\pid_side.O_1_24 ,\pid_side.O_1_23 ,\pid_side.O_1_22 ,\pid_side.O_1_21 ,\pid_side.O_1_20 ,\pid_side.O_1_19 ,\pid_side.O_1_18 ,\pid_side.O_1_17 ,\pid_side.O_1_16 ,\pid_side.O_1_15 ,\pid_side.O_1_14 ,\pid_side.O_1_13 ,\pid_side.O_1_12 ,\pid_side.O_1_11 ,\pid_side.O_1_10 ,\pid_side.O_1_9 ,\pid_side.O_1_8 ,\pid_side.O_1_7 ,\pid_side.O_1_6 ,\pid_side.O_1_5 ,\pid_side.O_1_4 ,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254}));
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42228),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42392),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270}),
            .ADDSUBBOT(),
            .A({N__52740,N__52770,N__51873,N__51909,N__51945,N__51981,N__52032,N__52086,N__52131,N__52173,N__51582,N__51627,N__51672,N__51708,N__51744,N__51786}),
            .C({dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286}),
            .B({dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,N__31971,N__30762,N__30729,N__29433,N__32010,N__32043,N__32075,N__32115}),
            .OHOLDTOP(),
            .O({dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,\pid_side.O_2_24 ,\pid_side.O_2_23 ,\pid_side.O_2_22 ,\pid_side.O_2_21 ,\pid_side.O_2_20 ,\pid_side.O_2_19 ,\pid_side.O_2_18 ,\pid_side.O_2_17 ,\pid_side.O_2_16 ,\pid_side.O_2_15 ,\pid_side.O_2_14 ,\pid_side.O_2_13 ,\pid_side.O_2_12 ,\pid_side.O_2_11 ,\pid_side.O_2_10 ,\pid_side.O_2_9 ,\pid_side.O_2_8 ,\pid_side.O_2_7 ,\pid_side.O_2_6 ,\pid_side.O_2_5 ,\pid_side.O_2_4 ,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305}));
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42459),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42285),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .ADDSUBBOT(),
            .A({N__39452,N__39494,N__38961,N__38993,N__39047,N__39095,N__39155,N__39206,N__39266,N__39327,N__38630,N__38684,N__38747,N__38795,N__38849,N__38916}),
            .C({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .B({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,N__55395,N__55605,N__55773,N__53253,N__55230,N__55950,N__56163,N__56334}),
            .OHOLDTOP(),
            .O({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,dangling_wire_352,\pid_front.O_24 ,\pid_front.O_23 ,\pid_front.O_22 ,\pid_front.O_21 ,\pid_front.O_20 ,\pid_front.O_19 ,\pid_front.O_18 ,\pid_front.O_17 ,\pid_front.O_16 ,\pid_front.O_15 ,\pid_front.O_14 ,\pid_front.O_13 ,\pid_front.O_12 ,\pid_front.O_11 ,\pid_front.O_10 ,\pid_front.O_9 ,\pid_front.O_8 ,\pid_front.O_7 ,\pid_front.O_6 ,\pid_front.O_5 ,\pid_front.O_4 ,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356}));
    IO_PAD \Pc2drone_pll_inst.Pc2drone_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__59697),
            .PACKAGEPIN(clk_system));
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__59683),
            .DIN(N__59682),
            .DOUT(N__59681),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__59683),
            .PADOUT(N__59682),
            .PADIN(N__59681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH2_18A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH2_18A_obuf_iopad (
            .OE(N__59674),
            .DIN(N__59673),
            .DOUT(N__59672),
            .PACKAGEPIN(debug_CH2_18A));
    defparam debug_CH2_18A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH2_18A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH2_18A_obuf_preio (
            .PADOEN(N__59674),
            .PADOUT(N__59673),
            .PADIN(N__59672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30354),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH0_16A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH0_16A_obuf_iopad (
            .OE(N__59665),
            .DIN(N__59664),
            .DOUT(N__59663),
            .PACKAGEPIN(debug_CH0_16A));
    defparam debug_CH0_16A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH0_16A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH0_16A_obuf_preio (
            .PADOEN(N__59665),
            .PADOUT(N__59664),
            .PADIN(N__59663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32904),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH1_0A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH1_0A_obuf_iopad (
            .OE(N__59656),
            .DIN(N__59655),
            .DOUT(N__59654),
            .PACKAGEPIN(debug_CH1_0A));
    defparam debug_CH1_0A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH1_0A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH1_0A_obuf_preio (
            .PADOEN(N__59656),
            .PADOUT(N__59655),
            .PADIN(N__59654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__47715),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH5_31B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH5_31B_obuf_iopad (
            .OE(N__59647),
            .DIN(N__59646),
            .DOUT(N__59645),
            .PACKAGEPIN(debug_CH5_31B));
    defparam debug_CH5_31B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH5_31B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH5_31B_obuf_preio (
            .PADOEN(N__59647),
            .PADOUT(N__59646),
            .PADIN(N__59645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH4_2A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH4_2A_obuf_iopad (
            .OE(N__59638),
            .DIN(N__59637),
            .DOUT(N__59636),
            .PACKAGEPIN(debug_CH4_2A));
    defparam debug_CH4_2A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH4_2A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH4_2A_obuf_preio (
            .PADOEN(N__59638),
            .PADOUT(N__59637),
            .PADIN(N__59636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__59629),
            .DIN(N__59628),
            .DOUT(N__59627),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__59629),
            .PADOUT(N__59628),
            .PADIN(N__59627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37641),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH3_20A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH3_20A_obuf_iopad (
            .OE(N__59620),
            .DIN(N__59619),
            .DOUT(N__59618),
            .PACKAGEPIN(debug_CH3_20A));
    defparam debug_CH3_20A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH3_20A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH3_20A_obuf_preio (
            .PADOEN(N__59620),
            .PADOUT(N__59619),
            .PADIN(N__59618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__41031),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH6_5B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH6_5B_obuf_iopad (
            .OE(N__59611),
            .DIN(N__59610),
            .DOUT(N__59609),
            .PACKAGEPIN(debug_CH6_5B));
    defparam debug_CH6_5B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH6_5B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH6_5B_obuf_preio (
            .PADOEN(N__59611),
            .PADOUT(N__59610),
            .PADIN(N__59609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__59602),
            .DIN(N__59601),
            .DOUT(N__59600),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__59602),
            .PADOUT(N__59601),
            .PADIN(N__59600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__14335 (
            .O(N__59583),
            .I(N__59580));
    LocalMux I__14334 (
            .O(N__59580),
            .I(N__59577));
    Odrv4 I__14333 (
            .O(N__59577),
            .I(\pid_front.O_22 ));
    InMux I__14332 (
            .O(N__59574),
            .I(N__59569));
    InMux I__14331 (
            .O(N__59573),
            .I(N__59566));
    InMux I__14330 (
            .O(N__59572),
            .I(N__59563));
    LocalMux I__14329 (
            .O(N__59569),
            .I(N__59560));
    LocalMux I__14328 (
            .O(N__59566),
            .I(N__59557));
    LocalMux I__14327 (
            .O(N__59563),
            .I(N__59554));
    Span12Mux_h I__14326 (
            .O(N__59560),
            .I(N__59551));
    Span12Mux_v I__14325 (
            .O(N__59557),
            .I(N__59546));
    Span12Mux_h I__14324 (
            .O(N__59554),
            .I(N__59546));
    Span12Mux_h I__14323 (
            .O(N__59551),
            .I(N__59543));
    Odrv12 I__14322 (
            .O(N__59546),
            .I(\pid_front.error_d_regZ0Z_18 ));
    Odrv12 I__14321 (
            .O(N__59543),
            .I(\pid_front.error_d_regZ0Z_18 ));
    InMux I__14320 (
            .O(N__59538),
            .I(N__59535));
    LocalMux I__14319 (
            .O(N__59535),
            .I(N__59532));
    Odrv4 I__14318 (
            .O(N__59532),
            .I(\pid_front.O_23 ));
    InMux I__14317 (
            .O(N__59529),
            .I(N__59520));
    InMux I__14316 (
            .O(N__59528),
            .I(N__59520));
    InMux I__14315 (
            .O(N__59527),
            .I(N__59520));
    LocalMux I__14314 (
            .O(N__59520),
            .I(N__59517));
    Span12Mux_h I__14313 (
            .O(N__59517),
            .I(N__59514));
    Odrv12 I__14312 (
            .O(N__59514),
            .I(\pid_front.error_d_regZ0Z_19 ));
    InMux I__14311 (
            .O(N__59511),
            .I(N__59508));
    LocalMux I__14310 (
            .O(N__59508),
            .I(N__59505));
    Odrv4 I__14309 (
            .O(N__59505),
            .I(\pid_front.O_24 ));
    InMux I__14308 (
            .O(N__59502),
            .I(N__59497));
    InMux I__14307 (
            .O(N__59501),
            .I(N__59492));
    InMux I__14306 (
            .O(N__59500),
            .I(N__59492));
    LocalMux I__14305 (
            .O(N__59497),
            .I(N__59487));
    LocalMux I__14304 (
            .O(N__59492),
            .I(N__59487));
    Span4Mux_h I__14303 (
            .O(N__59487),
            .I(N__59484));
    Span4Mux_h I__14302 (
            .O(N__59484),
            .I(N__59481));
    Span4Mux_h I__14301 (
            .O(N__59481),
            .I(N__59478));
    Odrv4 I__14300 (
            .O(N__59478),
            .I(\pid_front.error_d_regZ0Z_20 ));
    InMux I__14299 (
            .O(N__59475),
            .I(N__59472));
    LocalMux I__14298 (
            .O(N__59472),
            .I(N__59469));
    Odrv4 I__14297 (
            .O(N__59469),
            .I(\pid_front.O_18 ));
    InMux I__14296 (
            .O(N__59466),
            .I(N__59463));
    LocalMux I__14295 (
            .O(N__59463),
            .I(N__59460));
    Span4Mux_v I__14294 (
            .O(N__59460),
            .I(N__59455));
    InMux I__14293 (
            .O(N__59459),
            .I(N__59452));
    InMux I__14292 (
            .O(N__59458),
            .I(N__59449));
    Span4Mux_h I__14291 (
            .O(N__59455),
            .I(N__59446));
    LocalMux I__14290 (
            .O(N__59452),
            .I(N__59443));
    LocalMux I__14289 (
            .O(N__59449),
            .I(N__59436));
    Sp12to4 I__14288 (
            .O(N__59446),
            .I(N__59436));
    Span12Mux_h I__14287 (
            .O(N__59443),
            .I(N__59436));
    Odrv12 I__14286 (
            .O(N__59436),
            .I(\pid_front.error_d_regZ0Z_14 ));
    InMux I__14285 (
            .O(N__59433),
            .I(N__59430));
    LocalMux I__14284 (
            .O(N__59430),
            .I(\pid_front.O_8 ));
    InMux I__14283 (
            .O(N__59427),
            .I(N__59418));
    InMux I__14282 (
            .O(N__59426),
            .I(N__59418));
    InMux I__14281 (
            .O(N__59425),
            .I(N__59418));
    LocalMux I__14280 (
            .O(N__59418),
            .I(N__59415));
    Span4Mux_h I__14279 (
            .O(N__59415),
            .I(N__59412));
    Span4Mux_h I__14278 (
            .O(N__59412),
            .I(N__59409));
    Span4Mux_h I__14277 (
            .O(N__59409),
            .I(N__59406));
    Odrv4 I__14276 (
            .O(N__59406),
            .I(\pid_front.error_d_regZ0Z_4 ));
    InMux I__14275 (
            .O(N__59403),
            .I(N__59400));
    LocalMux I__14274 (
            .O(N__59400),
            .I(\pid_front.O_11 ));
    InMux I__14273 (
            .O(N__59397),
            .I(N__59392));
    InMux I__14272 (
            .O(N__59396),
            .I(N__59387));
    InMux I__14271 (
            .O(N__59395),
            .I(N__59387));
    LocalMux I__14270 (
            .O(N__59392),
            .I(N__59382));
    LocalMux I__14269 (
            .O(N__59387),
            .I(N__59382));
    Span4Mux_h I__14268 (
            .O(N__59382),
            .I(N__59379));
    Span4Mux_h I__14267 (
            .O(N__59379),
            .I(N__59376));
    Span4Mux_h I__14266 (
            .O(N__59376),
            .I(N__59373));
    Span4Mux_h I__14265 (
            .O(N__59373),
            .I(N__59370));
    Odrv4 I__14264 (
            .O(N__59370),
            .I(\pid_front.error_d_regZ0Z_7 ));
    InMux I__14263 (
            .O(N__59367),
            .I(N__59364));
    LocalMux I__14262 (
            .O(N__59364),
            .I(\pid_front.O_19 ));
    InMux I__14261 (
            .O(N__59361),
            .I(N__59352));
    InMux I__14260 (
            .O(N__59360),
            .I(N__59352));
    InMux I__14259 (
            .O(N__59359),
            .I(N__59352));
    LocalMux I__14258 (
            .O(N__59352),
            .I(N__59349));
    Span4Mux_v I__14257 (
            .O(N__59349),
            .I(N__59346));
    Sp12to4 I__14256 (
            .O(N__59346),
            .I(N__59343));
    Span12Mux_h I__14255 (
            .O(N__59343),
            .I(N__59340));
    Odrv12 I__14254 (
            .O(N__59340),
            .I(\pid_front.error_d_regZ0Z_15 ));
    ClkMux I__14253 (
            .O(N__59337),
            .I(N__58545));
    ClkMux I__14252 (
            .O(N__59336),
            .I(N__58545));
    ClkMux I__14251 (
            .O(N__59335),
            .I(N__58545));
    ClkMux I__14250 (
            .O(N__59334),
            .I(N__58545));
    ClkMux I__14249 (
            .O(N__59333),
            .I(N__58545));
    ClkMux I__14248 (
            .O(N__59332),
            .I(N__58545));
    ClkMux I__14247 (
            .O(N__59331),
            .I(N__58545));
    ClkMux I__14246 (
            .O(N__59330),
            .I(N__58545));
    ClkMux I__14245 (
            .O(N__59329),
            .I(N__58545));
    ClkMux I__14244 (
            .O(N__59328),
            .I(N__58545));
    ClkMux I__14243 (
            .O(N__59327),
            .I(N__58545));
    ClkMux I__14242 (
            .O(N__59326),
            .I(N__58545));
    ClkMux I__14241 (
            .O(N__59325),
            .I(N__58545));
    ClkMux I__14240 (
            .O(N__59324),
            .I(N__58545));
    ClkMux I__14239 (
            .O(N__59323),
            .I(N__58545));
    ClkMux I__14238 (
            .O(N__59322),
            .I(N__58545));
    ClkMux I__14237 (
            .O(N__59321),
            .I(N__58545));
    ClkMux I__14236 (
            .O(N__59320),
            .I(N__58545));
    ClkMux I__14235 (
            .O(N__59319),
            .I(N__58545));
    ClkMux I__14234 (
            .O(N__59318),
            .I(N__58545));
    ClkMux I__14233 (
            .O(N__59317),
            .I(N__58545));
    ClkMux I__14232 (
            .O(N__59316),
            .I(N__58545));
    ClkMux I__14231 (
            .O(N__59315),
            .I(N__58545));
    ClkMux I__14230 (
            .O(N__59314),
            .I(N__58545));
    ClkMux I__14229 (
            .O(N__59313),
            .I(N__58545));
    ClkMux I__14228 (
            .O(N__59312),
            .I(N__58545));
    ClkMux I__14227 (
            .O(N__59311),
            .I(N__58545));
    ClkMux I__14226 (
            .O(N__59310),
            .I(N__58545));
    ClkMux I__14225 (
            .O(N__59309),
            .I(N__58545));
    ClkMux I__14224 (
            .O(N__59308),
            .I(N__58545));
    ClkMux I__14223 (
            .O(N__59307),
            .I(N__58545));
    ClkMux I__14222 (
            .O(N__59306),
            .I(N__58545));
    ClkMux I__14221 (
            .O(N__59305),
            .I(N__58545));
    ClkMux I__14220 (
            .O(N__59304),
            .I(N__58545));
    ClkMux I__14219 (
            .O(N__59303),
            .I(N__58545));
    ClkMux I__14218 (
            .O(N__59302),
            .I(N__58545));
    ClkMux I__14217 (
            .O(N__59301),
            .I(N__58545));
    ClkMux I__14216 (
            .O(N__59300),
            .I(N__58545));
    ClkMux I__14215 (
            .O(N__59299),
            .I(N__58545));
    ClkMux I__14214 (
            .O(N__59298),
            .I(N__58545));
    ClkMux I__14213 (
            .O(N__59297),
            .I(N__58545));
    ClkMux I__14212 (
            .O(N__59296),
            .I(N__58545));
    ClkMux I__14211 (
            .O(N__59295),
            .I(N__58545));
    ClkMux I__14210 (
            .O(N__59294),
            .I(N__58545));
    ClkMux I__14209 (
            .O(N__59293),
            .I(N__58545));
    ClkMux I__14208 (
            .O(N__59292),
            .I(N__58545));
    ClkMux I__14207 (
            .O(N__59291),
            .I(N__58545));
    ClkMux I__14206 (
            .O(N__59290),
            .I(N__58545));
    ClkMux I__14205 (
            .O(N__59289),
            .I(N__58545));
    ClkMux I__14204 (
            .O(N__59288),
            .I(N__58545));
    ClkMux I__14203 (
            .O(N__59287),
            .I(N__58545));
    ClkMux I__14202 (
            .O(N__59286),
            .I(N__58545));
    ClkMux I__14201 (
            .O(N__59285),
            .I(N__58545));
    ClkMux I__14200 (
            .O(N__59284),
            .I(N__58545));
    ClkMux I__14199 (
            .O(N__59283),
            .I(N__58545));
    ClkMux I__14198 (
            .O(N__59282),
            .I(N__58545));
    ClkMux I__14197 (
            .O(N__59281),
            .I(N__58545));
    ClkMux I__14196 (
            .O(N__59280),
            .I(N__58545));
    ClkMux I__14195 (
            .O(N__59279),
            .I(N__58545));
    ClkMux I__14194 (
            .O(N__59278),
            .I(N__58545));
    ClkMux I__14193 (
            .O(N__59277),
            .I(N__58545));
    ClkMux I__14192 (
            .O(N__59276),
            .I(N__58545));
    ClkMux I__14191 (
            .O(N__59275),
            .I(N__58545));
    ClkMux I__14190 (
            .O(N__59274),
            .I(N__58545));
    ClkMux I__14189 (
            .O(N__59273),
            .I(N__58545));
    ClkMux I__14188 (
            .O(N__59272),
            .I(N__58545));
    ClkMux I__14187 (
            .O(N__59271),
            .I(N__58545));
    ClkMux I__14186 (
            .O(N__59270),
            .I(N__58545));
    ClkMux I__14185 (
            .O(N__59269),
            .I(N__58545));
    ClkMux I__14184 (
            .O(N__59268),
            .I(N__58545));
    ClkMux I__14183 (
            .O(N__59267),
            .I(N__58545));
    ClkMux I__14182 (
            .O(N__59266),
            .I(N__58545));
    ClkMux I__14181 (
            .O(N__59265),
            .I(N__58545));
    ClkMux I__14180 (
            .O(N__59264),
            .I(N__58545));
    ClkMux I__14179 (
            .O(N__59263),
            .I(N__58545));
    ClkMux I__14178 (
            .O(N__59262),
            .I(N__58545));
    ClkMux I__14177 (
            .O(N__59261),
            .I(N__58545));
    ClkMux I__14176 (
            .O(N__59260),
            .I(N__58545));
    ClkMux I__14175 (
            .O(N__59259),
            .I(N__58545));
    ClkMux I__14174 (
            .O(N__59258),
            .I(N__58545));
    ClkMux I__14173 (
            .O(N__59257),
            .I(N__58545));
    ClkMux I__14172 (
            .O(N__59256),
            .I(N__58545));
    ClkMux I__14171 (
            .O(N__59255),
            .I(N__58545));
    ClkMux I__14170 (
            .O(N__59254),
            .I(N__58545));
    ClkMux I__14169 (
            .O(N__59253),
            .I(N__58545));
    ClkMux I__14168 (
            .O(N__59252),
            .I(N__58545));
    ClkMux I__14167 (
            .O(N__59251),
            .I(N__58545));
    ClkMux I__14166 (
            .O(N__59250),
            .I(N__58545));
    ClkMux I__14165 (
            .O(N__59249),
            .I(N__58545));
    ClkMux I__14164 (
            .O(N__59248),
            .I(N__58545));
    ClkMux I__14163 (
            .O(N__59247),
            .I(N__58545));
    ClkMux I__14162 (
            .O(N__59246),
            .I(N__58545));
    ClkMux I__14161 (
            .O(N__59245),
            .I(N__58545));
    ClkMux I__14160 (
            .O(N__59244),
            .I(N__58545));
    ClkMux I__14159 (
            .O(N__59243),
            .I(N__58545));
    ClkMux I__14158 (
            .O(N__59242),
            .I(N__58545));
    ClkMux I__14157 (
            .O(N__59241),
            .I(N__58545));
    ClkMux I__14156 (
            .O(N__59240),
            .I(N__58545));
    ClkMux I__14155 (
            .O(N__59239),
            .I(N__58545));
    ClkMux I__14154 (
            .O(N__59238),
            .I(N__58545));
    ClkMux I__14153 (
            .O(N__59237),
            .I(N__58545));
    ClkMux I__14152 (
            .O(N__59236),
            .I(N__58545));
    ClkMux I__14151 (
            .O(N__59235),
            .I(N__58545));
    ClkMux I__14150 (
            .O(N__59234),
            .I(N__58545));
    ClkMux I__14149 (
            .O(N__59233),
            .I(N__58545));
    ClkMux I__14148 (
            .O(N__59232),
            .I(N__58545));
    ClkMux I__14147 (
            .O(N__59231),
            .I(N__58545));
    ClkMux I__14146 (
            .O(N__59230),
            .I(N__58545));
    ClkMux I__14145 (
            .O(N__59229),
            .I(N__58545));
    ClkMux I__14144 (
            .O(N__59228),
            .I(N__58545));
    ClkMux I__14143 (
            .O(N__59227),
            .I(N__58545));
    ClkMux I__14142 (
            .O(N__59226),
            .I(N__58545));
    ClkMux I__14141 (
            .O(N__59225),
            .I(N__58545));
    ClkMux I__14140 (
            .O(N__59224),
            .I(N__58545));
    ClkMux I__14139 (
            .O(N__59223),
            .I(N__58545));
    ClkMux I__14138 (
            .O(N__59222),
            .I(N__58545));
    ClkMux I__14137 (
            .O(N__59221),
            .I(N__58545));
    ClkMux I__14136 (
            .O(N__59220),
            .I(N__58545));
    ClkMux I__14135 (
            .O(N__59219),
            .I(N__58545));
    ClkMux I__14134 (
            .O(N__59218),
            .I(N__58545));
    ClkMux I__14133 (
            .O(N__59217),
            .I(N__58545));
    ClkMux I__14132 (
            .O(N__59216),
            .I(N__58545));
    ClkMux I__14131 (
            .O(N__59215),
            .I(N__58545));
    ClkMux I__14130 (
            .O(N__59214),
            .I(N__58545));
    ClkMux I__14129 (
            .O(N__59213),
            .I(N__58545));
    ClkMux I__14128 (
            .O(N__59212),
            .I(N__58545));
    ClkMux I__14127 (
            .O(N__59211),
            .I(N__58545));
    ClkMux I__14126 (
            .O(N__59210),
            .I(N__58545));
    ClkMux I__14125 (
            .O(N__59209),
            .I(N__58545));
    ClkMux I__14124 (
            .O(N__59208),
            .I(N__58545));
    ClkMux I__14123 (
            .O(N__59207),
            .I(N__58545));
    ClkMux I__14122 (
            .O(N__59206),
            .I(N__58545));
    ClkMux I__14121 (
            .O(N__59205),
            .I(N__58545));
    ClkMux I__14120 (
            .O(N__59204),
            .I(N__58545));
    ClkMux I__14119 (
            .O(N__59203),
            .I(N__58545));
    ClkMux I__14118 (
            .O(N__59202),
            .I(N__58545));
    ClkMux I__14117 (
            .O(N__59201),
            .I(N__58545));
    ClkMux I__14116 (
            .O(N__59200),
            .I(N__58545));
    ClkMux I__14115 (
            .O(N__59199),
            .I(N__58545));
    ClkMux I__14114 (
            .O(N__59198),
            .I(N__58545));
    ClkMux I__14113 (
            .O(N__59197),
            .I(N__58545));
    ClkMux I__14112 (
            .O(N__59196),
            .I(N__58545));
    ClkMux I__14111 (
            .O(N__59195),
            .I(N__58545));
    ClkMux I__14110 (
            .O(N__59194),
            .I(N__58545));
    ClkMux I__14109 (
            .O(N__59193),
            .I(N__58545));
    ClkMux I__14108 (
            .O(N__59192),
            .I(N__58545));
    ClkMux I__14107 (
            .O(N__59191),
            .I(N__58545));
    ClkMux I__14106 (
            .O(N__59190),
            .I(N__58545));
    ClkMux I__14105 (
            .O(N__59189),
            .I(N__58545));
    ClkMux I__14104 (
            .O(N__59188),
            .I(N__58545));
    ClkMux I__14103 (
            .O(N__59187),
            .I(N__58545));
    ClkMux I__14102 (
            .O(N__59186),
            .I(N__58545));
    ClkMux I__14101 (
            .O(N__59185),
            .I(N__58545));
    ClkMux I__14100 (
            .O(N__59184),
            .I(N__58545));
    ClkMux I__14099 (
            .O(N__59183),
            .I(N__58545));
    ClkMux I__14098 (
            .O(N__59182),
            .I(N__58545));
    ClkMux I__14097 (
            .O(N__59181),
            .I(N__58545));
    ClkMux I__14096 (
            .O(N__59180),
            .I(N__58545));
    ClkMux I__14095 (
            .O(N__59179),
            .I(N__58545));
    ClkMux I__14094 (
            .O(N__59178),
            .I(N__58545));
    ClkMux I__14093 (
            .O(N__59177),
            .I(N__58545));
    ClkMux I__14092 (
            .O(N__59176),
            .I(N__58545));
    ClkMux I__14091 (
            .O(N__59175),
            .I(N__58545));
    ClkMux I__14090 (
            .O(N__59174),
            .I(N__58545));
    ClkMux I__14089 (
            .O(N__59173),
            .I(N__58545));
    ClkMux I__14088 (
            .O(N__59172),
            .I(N__58545));
    ClkMux I__14087 (
            .O(N__59171),
            .I(N__58545));
    ClkMux I__14086 (
            .O(N__59170),
            .I(N__58545));
    ClkMux I__14085 (
            .O(N__59169),
            .I(N__58545));
    ClkMux I__14084 (
            .O(N__59168),
            .I(N__58545));
    ClkMux I__14083 (
            .O(N__59167),
            .I(N__58545));
    ClkMux I__14082 (
            .O(N__59166),
            .I(N__58545));
    ClkMux I__14081 (
            .O(N__59165),
            .I(N__58545));
    ClkMux I__14080 (
            .O(N__59164),
            .I(N__58545));
    ClkMux I__14079 (
            .O(N__59163),
            .I(N__58545));
    ClkMux I__14078 (
            .O(N__59162),
            .I(N__58545));
    ClkMux I__14077 (
            .O(N__59161),
            .I(N__58545));
    ClkMux I__14076 (
            .O(N__59160),
            .I(N__58545));
    ClkMux I__14075 (
            .O(N__59159),
            .I(N__58545));
    ClkMux I__14074 (
            .O(N__59158),
            .I(N__58545));
    ClkMux I__14073 (
            .O(N__59157),
            .I(N__58545));
    ClkMux I__14072 (
            .O(N__59156),
            .I(N__58545));
    ClkMux I__14071 (
            .O(N__59155),
            .I(N__58545));
    ClkMux I__14070 (
            .O(N__59154),
            .I(N__58545));
    ClkMux I__14069 (
            .O(N__59153),
            .I(N__58545));
    ClkMux I__14068 (
            .O(N__59152),
            .I(N__58545));
    ClkMux I__14067 (
            .O(N__59151),
            .I(N__58545));
    ClkMux I__14066 (
            .O(N__59150),
            .I(N__58545));
    ClkMux I__14065 (
            .O(N__59149),
            .I(N__58545));
    ClkMux I__14064 (
            .O(N__59148),
            .I(N__58545));
    ClkMux I__14063 (
            .O(N__59147),
            .I(N__58545));
    ClkMux I__14062 (
            .O(N__59146),
            .I(N__58545));
    ClkMux I__14061 (
            .O(N__59145),
            .I(N__58545));
    ClkMux I__14060 (
            .O(N__59144),
            .I(N__58545));
    ClkMux I__14059 (
            .O(N__59143),
            .I(N__58545));
    ClkMux I__14058 (
            .O(N__59142),
            .I(N__58545));
    ClkMux I__14057 (
            .O(N__59141),
            .I(N__58545));
    ClkMux I__14056 (
            .O(N__59140),
            .I(N__58545));
    ClkMux I__14055 (
            .O(N__59139),
            .I(N__58545));
    ClkMux I__14054 (
            .O(N__59138),
            .I(N__58545));
    ClkMux I__14053 (
            .O(N__59137),
            .I(N__58545));
    ClkMux I__14052 (
            .O(N__59136),
            .I(N__58545));
    ClkMux I__14051 (
            .O(N__59135),
            .I(N__58545));
    ClkMux I__14050 (
            .O(N__59134),
            .I(N__58545));
    ClkMux I__14049 (
            .O(N__59133),
            .I(N__58545));
    ClkMux I__14048 (
            .O(N__59132),
            .I(N__58545));
    ClkMux I__14047 (
            .O(N__59131),
            .I(N__58545));
    ClkMux I__14046 (
            .O(N__59130),
            .I(N__58545));
    ClkMux I__14045 (
            .O(N__59129),
            .I(N__58545));
    ClkMux I__14044 (
            .O(N__59128),
            .I(N__58545));
    ClkMux I__14043 (
            .O(N__59127),
            .I(N__58545));
    ClkMux I__14042 (
            .O(N__59126),
            .I(N__58545));
    ClkMux I__14041 (
            .O(N__59125),
            .I(N__58545));
    ClkMux I__14040 (
            .O(N__59124),
            .I(N__58545));
    ClkMux I__14039 (
            .O(N__59123),
            .I(N__58545));
    ClkMux I__14038 (
            .O(N__59122),
            .I(N__58545));
    ClkMux I__14037 (
            .O(N__59121),
            .I(N__58545));
    ClkMux I__14036 (
            .O(N__59120),
            .I(N__58545));
    ClkMux I__14035 (
            .O(N__59119),
            .I(N__58545));
    ClkMux I__14034 (
            .O(N__59118),
            .I(N__58545));
    ClkMux I__14033 (
            .O(N__59117),
            .I(N__58545));
    ClkMux I__14032 (
            .O(N__59116),
            .I(N__58545));
    ClkMux I__14031 (
            .O(N__59115),
            .I(N__58545));
    ClkMux I__14030 (
            .O(N__59114),
            .I(N__58545));
    ClkMux I__14029 (
            .O(N__59113),
            .I(N__58545));
    ClkMux I__14028 (
            .O(N__59112),
            .I(N__58545));
    ClkMux I__14027 (
            .O(N__59111),
            .I(N__58545));
    ClkMux I__14026 (
            .O(N__59110),
            .I(N__58545));
    ClkMux I__14025 (
            .O(N__59109),
            .I(N__58545));
    ClkMux I__14024 (
            .O(N__59108),
            .I(N__58545));
    ClkMux I__14023 (
            .O(N__59107),
            .I(N__58545));
    ClkMux I__14022 (
            .O(N__59106),
            .I(N__58545));
    ClkMux I__14021 (
            .O(N__59105),
            .I(N__58545));
    ClkMux I__14020 (
            .O(N__59104),
            .I(N__58545));
    ClkMux I__14019 (
            .O(N__59103),
            .I(N__58545));
    ClkMux I__14018 (
            .O(N__59102),
            .I(N__58545));
    ClkMux I__14017 (
            .O(N__59101),
            .I(N__58545));
    ClkMux I__14016 (
            .O(N__59100),
            .I(N__58545));
    ClkMux I__14015 (
            .O(N__59099),
            .I(N__58545));
    ClkMux I__14014 (
            .O(N__59098),
            .I(N__58545));
    ClkMux I__14013 (
            .O(N__59097),
            .I(N__58545));
    ClkMux I__14012 (
            .O(N__59096),
            .I(N__58545));
    ClkMux I__14011 (
            .O(N__59095),
            .I(N__58545));
    ClkMux I__14010 (
            .O(N__59094),
            .I(N__58545));
    ClkMux I__14009 (
            .O(N__59093),
            .I(N__58545));
    ClkMux I__14008 (
            .O(N__59092),
            .I(N__58545));
    ClkMux I__14007 (
            .O(N__59091),
            .I(N__58545));
    ClkMux I__14006 (
            .O(N__59090),
            .I(N__58545));
    ClkMux I__14005 (
            .O(N__59089),
            .I(N__58545));
    ClkMux I__14004 (
            .O(N__59088),
            .I(N__58545));
    ClkMux I__14003 (
            .O(N__59087),
            .I(N__58545));
    ClkMux I__14002 (
            .O(N__59086),
            .I(N__58545));
    ClkMux I__14001 (
            .O(N__59085),
            .I(N__58545));
    ClkMux I__14000 (
            .O(N__59084),
            .I(N__58545));
    ClkMux I__13999 (
            .O(N__59083),
            .I(N__58545));
    ClkMux I__13998 (
            .O(N__59082),
            .I(N__58545));
    ClkMux I__13997 (
            .O(N__59081),
            .I(N__58545));
    ClkMux I__13996 (
            .O(N__59080),
            .I(N__58545));
    ClkMux I__13995 (
            .O(N__59079),
            .I(N__58545));
    ClkMux I__13994 (
            .O(N__59078),
            .I(N__58545));
    ClkMux I__13993 (
            .O(N__59077),
            .I(N__58545));
    ClkMux I__13992 (
            .O(N__59076),
            .I(N__58545));
    ClkMux I__13991 (
            .O(N__59075),
            .I(N__58545));
    ClkMux I__13990 (
            .O(N__59074),
            .I(N__58545));
    GlobalMux I__13989 (
            .O(N__58545),
            .I(N__58542));
    gio2CtrlBuf I__13988 (
            .O(N__58542),
            .I(clk_system_pll_g));
    CEMux I__13987 (
            .O(N__58539),
            .I(N__58531));
    CEMux I__13986 (
            .O(N__58538),
            .I(N__58528));
    CEMux I__13985 (
            .O(N__58537),
            .I(N__58525));
    CEMux I__13984 (
            .O(N__58536),
            .I(N__58520));
    CEMux I__13983 (
            .O(N__58535),
            .I(N__58517));
    CEMux I__13982 (
            .O(N__58534),
            .I(N__58514));
    LocalMux I__13981 (
            .O(N__58531),
            .I(N__58511));
    LocalMux I__13980 (
            .O(N__58528),
            .I(N__58508));
    LocalMux I__13979 (
            .O(N__58525),
            .I(N__58504));
    CEMux I__13978 (
            .O(N__58524),
            .I(N__58499));
    CEMux I__13977 (
            .O(N__58523),
            .I(N__58496));
    LocalMux I__13976 (
            .O(N__58520),
            .I(N__58491));
    LocalMux I__13975 (
            .O(N__58517),
            .I(N__58486));
    LocalMux I__13974 (
            .O(N__58514),
            .I(N__58486));
    Span4Mux_v I__13973 (
            .O(N__58511),
            .I(N__58483));
    Span4Mux_s3_h I__13972 (
            .O(N__58508),
            .I(N__58480));
    CEMux I__13971 (
            .O(N__58507),
            .I(N__58477));
    Span4Mux_s3_h I__13970 (
            .O(N__58504),
            .I(N__58474));
    CEMux I__13969 (
            .O(N__58503),
            .I(N__58471));
    CEMux I__13968 (
            .O(N__58502),
            .I(N__58468));
    LocalMux I__13967 (
            .O(N__58499),
            .I(N__58465));
    LocalMux I__13966 (
            .O(N__58496),
            .I(N__58462));
    CEMux I__13965 (
            .O(N__58495),
            .I(N__58459));
    CEMux I__13964 (
            .O(N__58494),
            .I(N__58456));
    Span4Mux_s1_h I__13963 (
            .O(N__58491),
            .I(N__58450));
    Span4Mux_v I__13962 (
            .O(N__58486),
            .I(N__58450));
    Span4Mux_v I__13961 (
            .O(N__58483),
            .I(N__58446));
    Span4Mux_v I__13960 (
            .O(N__58480),
            .I(N__58443));
    LocalMux I__13959 (
            .O(N__58477),
            .I(N__58440));
    Span4Mux_h I__13958 (
            .O(N__58474),
            .I(N__58435));
    LocalMux I__13957 (
            .O(N__58471),
            .I(N__58435));
    LocalMux I__13956 (
            .O(N__58468),
            .I(N__58432));
    Span4Mux_s2_h I__13955 (
            .O(N__58465),
            .I(N__58423));
    Span4Mux_s2_h I__13954 (
            .O(N__58462),
            .I(N__58423));
    LocalMux I__13953 (
            .O(N__58459),
            .I(N__58423));
    LocalMux I__13952 (
            .O(N__58456),
            .I(N__58423));
    CEMux I__13951 (
            .O(N__58455),
            .I(N__58420));
    Span4Mux_h I__13950 (
            .O(N__58450),
            .I(N__58417));
    CEMux I__13949 (
            .O(N__58449),
            .I(N__58414));
    Span4Mux_h I__13948 (
            .O(N__58446),
            .I(N__58411));
    Span4Mux_h I__13947 (
            .O(N__58443),
            .I(N__58408));
    Span4Mux_h I__13946 (
            .O(N__58440),
            .I(N__58405));
    Span4Mux_h I__13945 (
            .O(N__58435),
            .I(N__58402));
    Span4Mux_h I__13944 (
            .O(N__58432),
            .I(N__58395));
    Span4Mux_h I__13943 (
            .O(N__58423),
            .I(N__58395));
    LocalMux I__13942 (
            .O(N__58420),
            .I(N__58395));
    Span4Mux_h I__13941 (
            .O(N__58417),
            .I(N__58392));
    LocalMux I__13940 (
            .O(N__58414),
            .I(N__58389));
    Span4Mux_h I__13939 (
            .O(N__58411),
            .I(N__58386));
    Span4Mux_h I__13938 (
            .O(N__58408),
            .I(N__58383));
    Span4Mux_v I__13937 (
            .O(N__58405),
            .I(N__58378));
    Span4Mux_v I__13936 (
            .O(N__58402),
            .I(N__58378));
    Span4Mux_h I__13935 (
            .O(N__58395),
            .I(N__58375));
    Span4Mux_h I__13934 (
            .O(N__58392),
            .I(N__58370));
    Span4Mux_h I__13933 (
            .O(N__58389),
            .I(N__58370));
    Odrv4 I__13932 (
            .O(N__58386),
            .I(\pid_front.N_543_0 ));
    Odrv4 I__13931 (
            .O(N__58383),
            .I(\pid_front.N_543_0 ));
    Odrv4 I__13930 (
            .O(N__58378),
            .I(\pid_front.N_543_0 ));
    Odrv4 I__13929 (
            .O(N__58375),
            .I(\pid_front.N_543_0 ));
    Odrv4 I__13928 (
            .O(N__58370),
            .I(\pid_front.N_543_0 ));
    InMux I__13927 (
            .O(N__58359),
            .I(N__58314));
    InMux I__13926 (
            .O(N__58358),
            .I(N__58314));
    InMux I__13925 (
            .O(N__58357),
            .I(N__58305));
    InMux I__13924 (
            .O(N__58356),
            .I(N__58305));
    InMux I__13923 (
            .O(N__58355),
            .I(N__58305));
    InMux I__13922 (
            .O(N__58354),
            .I(N__58305));
    InMux I__13921 (
            .O(N__58353),
            .I(N__58300));
    InMux I__13920 (
            .O(N__58352),
            .I(N__58300));
    InMux I__13919 (
            .O(N__58351),
            .I(N__58295));
    InMux I__13918 (
            .O(N__58350),
            .I(N__58295));
    InMux I__13917 (
            .O(N__58349),
            .I(N__58286));
    InMux I__13916 (
            .O(N__58348),
            .I(N__58286));
    InMux I__13915 (
            .O(N__58347),
            .I(N__58286));
    InMux I__13914 (
            .O(N__58346),
            .I(N__58286));
    InMux I__13913 (
            .O(N__58345),
            .I(N__58281));
    InMux I__13912 (
            .O(N__58344),
            .I(N__58281));
    InMux I__13911 (
            .O(N__58343),
            .I(N__58276));
    InMux I__13910 (
            .O(N__58342),
            .I(N__58276));
    InMux I__13909 (
            .O(N__58341),
            .I(N__58265));
    InMux I__13908 (
            .O(N__58340),
            .I(N__58265));
    InMux I__13907 (
            .O(N__58339),
            .I(N__58265));
    InMux I__13906 (
            .O(N__58338),
            .I(N__58265));
    InMux I__13905 (
            .O(N__58337),
            .I(N__58265));
    InMux I__13904 (
            .O(N__58336),
            .I(N__58262));
    InMux I__13903 (
            .O(N__58335),
            .I(N__58257));
    InMux I__13902 (
            .O(N__58334),
            .I(N__58257));
    InMux I__13901 (
            .O(N__58333),
            .I(N__58252));
    InMux I__13900 (
            .O(N__58332),
            .I(N__58252));
    InMux I__13899 (
            .O(N__58331),
            .I(N__58247));
    InMux I__13898 (
            .O(N__58330),
            .I(N__58247));
    InMux I__13897 (
            .O(N__58329),
            .I(N__58232));
    InMux I__13896 (
            .O(N__58328),
            .I(N__58232));
    InMux I__13895 (
            .O(N__58327),
            .I(N__58232));
    InMux I__13894 (
            .O(N__58326),
            .I(N__58232));
    InMux I__13893 (
            .O(N__58325),
            .I(N__58232));
    InMux I__13892 (
            .O(N__58324),
            .I(N__58232));
    InMux I__13891 (
            .O(N__58323),
            .I(N__58232));
    InMux I__13890 (
            .O(N__58322),
            .I(N__58229));
    InMux I__13889 (
            .O(N__58321),
            .I(N__58226));
    InMux I__13888 (
            .O(N__58320),
            .I(N__58223));
    InMux I__13887 (
            .O(N__58319),
            .I(N__58220));
    LocalMux I__13886 (
            .O(N__58314),
            .I(N__58176));
    LocalMux I__13885 (
            .O(N__58305),
            .I(N__58173));
    LocalMux I__13884 (
            .O(N__58300),
            .I(N__58170));
    LocalMux I__13883 (
            .O(N__58295),
            .I(N__58167));
    LocalMux I__13882 (
            .O(N__58286),
            .I(N__58164));
    LocalMux I__13881 (
            .O(N__58281),
            .I(N__58161));
    LocalMux I__13880 (
            .O(N__58276),
            .I(N__58158));
    LocalMux I__13879 (
            .O(N__58265),
            .I(N__58155));
    LocalMux I__13878 (
            .O(N__58262),
            .I(N__58152));
    LocalMux I__13877 (
            .O(N__58257),
            .I(N__58149));
    LocalMux I__13876 (
            .O(N__58252),
            .I(N__58146));
    LocalMux I__13875 (
            .O(N__58247),
            .I(N__58143));
    LocalMux I__13874 (
            .O(N__58232),
            .I(N__58140));
    LocalMux I__13873 (
            .O(N__58229),
            .I(N__58137));
    LocalMux I__13872 (
            .O(N__58226),
            .I(N__58134));
    LocalMux I__13871 (
            .O(N__58223),
            .I(N__58131));
    LocalMux I__13870 (
            .O(N__58220),
            .I(N__58128));
    SRMux I__13869 (
            .O(N__58219),
            .I(N__58011));
    SRMux I__13868 (
            .O(N__58218),
            .I(N__58011));
    SRMux I__13867 (
            .O(N__58217),
            .I(N__58011));
    SRMux I__13866 (
            .O(N__58216),
            .I(N__58011));
    SRMux I__13865 (
            .O(N__58215),
            .I(N__58011));
    SRMux I__13864 (
            .O(N__58214),
            .I(N__58011));
    SRMux I__13863 (
            .O(N__58213),
            .I(N__58011));
    SRMux I__13862 (
            .O(N__58212),
            .I(N__58011));
    SRMux I__13861 (
            .O(N__58211),
            .I(N__58011));
    SRMux I__13860 (
            .O(N__58210),
            .I(N__58011));
    SRMux I__13859 (
            .O(N__58209),
            .I(N__58011));
    SRMux I__13858 (
            .O(N__58208),
            .I(N__58011));
    SRMux I__13857 (
            .O(N__58207),
            .I(N__58011));
    SRMux I__13856 (
            .O(N__58206),
            .I(N__58011));
    SRMux I__13855 (
            .O(N__58205),
            .I(N__58011));
    SRMux I__13854 (
            .O(N__58204),
            .I(N__58011));
    SRMux I__13853 (
            .O(N__58203),
            .I(N__58011));
    SRMux I__13852 (
            .O(N__58202),
            .I(N__58011));
    SRMux I__13851 (
            .O(N__58201),
            .I(N__58011));
    SRMux I__13850 (
            .O(N__58200),
            .I(N__58011));
    SRMux I__13849 (
            .O(N__58199),
            .I(N__58011));
    SRMux I__13848 (
            .O(N__58198),
            .I(N__58011));
    SRMux I__13847 (
            .O(N__58197),
            .I(N__58011));
    SRMux I__13846 (
            .O(N__58196),
            .I(N__58011));
    SRMux I__13845 (
            .O(N__58195),
            .I(N__58011));
    SRMux I__13844 (
            .O(N__58194),
            .I(N__58011));
    SRMux I__13843 (
            .O(N__58193),
            .I(N__58011));
    SRMux I__13842 (
            .O(N__58192),
            .I(N__58011));
    SRMux I__13841 (
            .O(N__58191),
            .I(N__58011));
    SRMux I__13840 (
            .O(N__58190),
            .I(N__58011));
    SRMux I__13839 (
            .O(N__58189),
            .I(N__58011));
    SRMux I__13838 (
            .O(N__58188),
            .I(N__58011));
    SRMux I__13837 (
            .O(N__58187),
            .I(N__58011));
    SRMux I__13836 (
            .O(N__58186),
            .I(N__58011));
    SRMux I__13835 (
            .O(N__58185),
            .I(N__58011));
    SRMux I__13834 (
            .O(N__58184),
            .I(N__58011));
    SRMux I__13833 (
            .O(N__58183),
            .I(N__58011));
    SRMux I__13832 (
            .O(N__58182),
            .I(N__58011));
    SRMux I__13831 (
            .O(N__58181),
            .I(N__58011));
    SRMux I__13830 (
            .O(N__58180),
            .I(N__58011));
    SRMux I__13829 (
            .O(N__58179),
            .I(N__58011));
    Glb2LocalMux I__13828 (
            .O(N__58176),
            .I(N__58011));
    Glb2LocalMux I__13827 (
            .O(N__58173),
            .I(N__58011));
    Glb2LocalMux I__13826 (
            .O(N__58170),
            .I(N__58011));
    Glb2LocalMux I__13825 (
            .O(N__58167),
            .I(N__58011));
    Glb2LocalMux I__13824 (
            .O(N__58164),
            .I(N__58011));
    Glb2LocalMux I__13823 (
            .O(N__58161),
            .I(N__58011));
    Glb2LocalMux I__13822 (
            .O(N__58158),
            .I(N__58011));
    Glb2LocalMux I__13821 (
            .O(N__58155),
            .I(N__58011));
    Glb2LocalMux I__13820 (
            .O(N__58152),
            .I(N__58011));
    Glb2LocalMux I__13819 (
            .O(N__58149),
            .I(N__58011));
    Glb2LocalMux I__13818 (
            .O(N__58146),
            .I(N__58011));
    Glb2LocalMux I__13817 (
            .O(N__58143),
            .I(N__58011));
    Glb2LocalMux I__13816 (
            .O(N__58140),
            .I(N__58011));
    Glb2LocalMux I__13815 (
            .O(N__58137),
            .I(N__58011));
    Glb2LocalMux I__13814 (
            .O(N__58134),
            .I(N__58011));
    Glb2LocalMux I__13813 (
            .O(N__58131),
            .I(N__58011));
    Glb2LocalMux I__13812 (
            .O(N__58128),
            .I(N__58011));
    GlobalMux I__13811 (
            .O(N__58011),
            .I(N__58008));
    gio2CtrlBuf I__13810 (
            .O(N__58008),
            .I(N_665_g));
    InMux I__13809 (
            .O(N__58005),
            .I(N__58001));
    InMux I__13808 (
            .O(N__58004),
            .I(N__57998));
    LocalMux I__13807 (
            .O(N__58001),
            .I(N__57994));
    LocalMux I__13806 (
            .O(N__57998),
            .I(N__57991));
    InMux I__13805 (
            .O(N__57997),
            .I(N__57988));
    Odrv12 I__13804 (
            .O(N__57994),
            .I(\pid_side.error_d_regZ0Z_20 ));
    Odrv4 I__13803 (
            .O(N__57991),
            .I(\pid_side.error_d_regZ0Z_20 ));
    LocalMux I__13802 (
            .O(N__57988),
            .I(\pid_side.error_d_regZ0Z_20 ));
    InMux I__13801 (
            .O(N__57981),
            .I(N__57977));
    InMux I__13800 (
            .O(N__57980),
            .I(N__57974));
    LocalMux I__13799 (
            .O(N__57977),
            .I(N__57969));
    LocalMux I__13798 (
            .O(N__57974),
            .I(N__57969));
    Odrv4 I__13797 (
            .O(N__57969),
            .I(\pid_side.error_d_reg_prevZ0Z_20 ));
    CEMux I__13796 (
            .O(N__57966),
            .I(N__57909));
    CEMux I__13795 (
            .O(N__57965),
            .I(N__57909));
    CEMux I__13794 (
            .O(N__57964),
            .I(N__57909));
    CEMux I__13793 (
            .O(N__57963),
            .I(N__57909));
    CEMux I__13792 (
            .O(N__57962),
            .I(N__57909));
    CEMux I__13791 (
            .O(N__57961),
            .I(N__57909));
    CEMux I__13790 (
            .O(N__57960),
            .I(N__57909));
    CEMux I__13789 (
            .O(N__57959),
            .I(N__57909));
    CEMux I__13788 (
            .O(N__57958),
            .I(N__57909));
    CEMux I__13787 (
            .O(N__57957),
            .I(N__57909));
    CEMux I__13786 (
            .O(N__57956),
            .I(N__57909));
    CEMux I__13785 (
            .O(N__57955),
            .I(N__57909));
    CEMux I__13784 (
            .O(N__57954),
            .I(N__57909));
    CEMux I__13783 (
            .O(N__57953),
            .I(N__57909));
    CEMux I__13782 (
            .O(N__57952),
            .I(N__57909));
    CEMux I__13781 (
            .O(N__57951),
            .I(N__57909));
    CEMux I__13780 (
            .O(N__57950),
            .I(N__57909));
    CEMux I__13779 (
            .O(N__57949),
            .I(N__57909));
    CEMux I__13778 (
            .O(N__57948),
            .I(N__57909));
    GlobalMux I__13777 (
            .O(N__57909),
            .I(N__57906));
    gio2CtrlBuf I__13776 (
            .O(N__57906),
            .I(\pid_side.state_0_g_0 ));
    CascadeMux I__13775 (
            .O(N__57903),
            .I(N__57897));
    CascadeMux I__13774 (
            .O(N__57902),
            .I(N__57891));
    CascadeMux I__13773 (
            .O(N__57901),
            .I(N__57872));
    CascadeMux I__13772 (
            .O(N__57900),
            .I(N__57838));
    InMux I__13771 (
            .O(N__57897),
            .I(N__57824));
    InMux I__13770 (
            .O(N__57896),
            .I(N__57821));
    InMux I__13769 (
            .O(N__57895),
            .I(N__57818));
    InMux I__13768 (
            .O(N__57894),
            .I(N__57811));
    InMux I__13767 (
            .O(N__57891),
            .I(N__57811));
    InMux I__13766 (
            .O(N__57890),
            .I(N__57811));
    InMux I__13765 (
            .O(N__57889),
            .I(N__57808));
    InMux I__13764 (
            .O(N__57888),
            .I(N__57799));
    InMux I__13763 (
            .O(N__57887),
            .I(N__57799));
    InMux I__13762 (
            .O(N__57886),
            .I(N__57799));
    InMux I__13761 (
            .O(N__57885),
            .I(N__57799));
    InMux I__13760 (
            .O(N__57884),
            .I(N__57794));
    InMux I__13759 (
            .O(N__57883),
            .I(N__57794));
    InMux I__13758 (
            .O(N__57882),
            .I(N__57787));
    InMux I__13757 (
            .O(N__57881),
            .I(N__57787));
    InMux I__13756 (
            .O(N__57880),
            .I(N__57787));
    InMux I__13755 (
            .O(N__57879),
            .I(N__57782));
    InMux I__13754 (
            .O(N__57878),
            .I(N__57782));
    InMux I__13753 (
            .O(N__57877),
            .I(N__57775));
    InMux I__13752 (
            .O(N__57876),
            .I(N__57775));
    InMux I__13751 (
            .O(N__57875),
            .I(N__57775));
    InMux I__13750 (
            .O(N__57872),
            .I(N__57770));
    InMux I__13749 (
            .O(N__57871),
            .I(N__57770));
    InMux I__13748 (
            .O(N__57870),
            .I(N__57767));
    InMux I__13747 (
            .O(N__57869),
            .I(N__57760));
    InMux I__13746 (
            .O(N__57868),
            .I(N__57760));
    InMux I__13745 (
            .O(N__57867),
            .I(N__57760));
    InMux I__13744 (
            .O(N__57866),
            .I(N__57757));
    InMux I__13743 (
            .O(N__57865),
            .I(N__57754));
    InMux I__13742 (
            .O(N__57864),
            .I(N__57751));
    InMux I__13741 (
            .O(N__57863),
            .I(N__57746));
    InMux I__13740 (
            .O(N__57862),
            .I(N__57746));
    InMux I__13739 (
            .O(N__57861),
            .I(N__57743));
    InMux I__13738 (
            .O(N__57860),
            .I(N__57740));
    InMux I__13737 (
            .O(N__57859),
            .I(N__57737));
    InMux I__13736 (
            .O(N__57858),
            .I(N__57734));
    InMux I__13735 (
            .O(N__57857),
            .I(N__57727));
    InMux I__13734 (
            .O(N__57856),
            .I(N__57727));
    InMux I__13733 (
            .O(N__57855),
            .I(N__57727));
    InMux I__13732 (
            .O(N__57854),
            .I(N__57724));
    InMux I__13731 (
            .O(N__57853),
            .I(N__57719));
    InMux I__13730 (
            .O(N__57852),
            .I(N__57719));
    InMux I__13729 (
            .O(N__57851),
            .I(N__57716));
    InMux I__13728 (
            .O(N__57850),
            .I(N__57713));
    InMux I__13727 (
            .O(N__57849),
            .I(N__57710));
    InMux I__13726 (
            .O(N__57848),
            .I(N__57707));
    InMux I__13725 (
            .O(N__57847),
            .I(N__57704));
    InMux I__13724 (
            .O(N__57846),
            .I(N__57701));
    InMux I__13723 (
            .O(N__57845),
            .I(N__57698));
    InMux I__13722 (
            .O(N__57844),
            .I(N__57695));
    InMux I__13721 (
            .O(N__57843),
            .I(N__57690));
    InMux I__13720 (
            .O(N__57842),
            .I(N__57690));
    InMux I__13719 (
            .O(N__57841),
            .I(N__57687));
    InMux I__13718 (
            .O(N__57838),
            .I(N__57684));
    InMux I__13717 (
            .O(N__57837),
            .I(N__57681));
    InMux I__13716 (
            .O(N__57836),
            .I(N__57678));
    InMux I__13715 (
            .O(N__57835),
            .I(N__57675));
    InMux I__13714 (
            .O(N__57834),
            .I(N__57672));
    InMux I__13713 (
            .O(N__57833),
            .I(N__57669));
    InMux I__13712 (
            .O(N__57832),
            .I(N__57666));
    InMux I__13711 (
            .O(N__57831),
            .I(N__57663));
    InMux I__13710 (
            .O(N__57830),
            .I(N__57660));
    InMux I__13709 (
            .O(N__57829),
            .I(N__57657));
    InMux I__13708 (
            .O(N__57828),
            .I(N__57654));
    InMux I__13707 (
            .O(N__57827),
            .I(N__57651));
    LocalMux I__13706 (
            .O(N__57824),
            .I(N__57493));
    LocalMux I__13705 (
            .O(N__57821),
            .I(N__57490));
    LocalMux I__13704 (
            .O(N__57818),
            .I(N__57487));
    LocalMux I__13703 (
            .O(N__57811),
            .I(N__57484));
    LocalMux I__13702 (
            .O(N__57808),
            .I(N__57481));
    LocalMux I__13701 (
            .O(N__57799),
            .I(N__57478));
    LocalMux I__13700 (
            .O(N__57794),
            .I(N__57475));
    LocalMux I__13699 (
            .O(N__57787),
            .I(N__57472));
    LocalMux I__13698 (
            .O(N__57782),
            .I(N__57469));
    LocalMux I__13697 (
            .O(N__57775),
            .I(N__57466));
    LocalMux I__13696 (
            .O(N__57770),
            .I(N__57463));
    LocalMux I__13695 (
            .O(N__57767),
            .I(N__57460));
    LocalMux I__13694 (
            .O(N__57760),
            .I(N__57457));
    LocalMux I__13693 (
            .O(N__57757),
            .I(N__57454));
    LocalMux I__13692 (
            .O(N__57754),
            .I(N__57451));
    LocalMux I__13691 (
            .O(N__57751),
            .I(N__57448));
    LocalMux I__13690 (
            .O(N__57746),
            .I(N__57445));
    LocalMux I__13689 (
            .O(N__57743),
            .I(N__57442));
    LocalMux I__13688 (
            .O(N__57740),
            .I(N__57439));
    LocalMux I__13687 (
            .O(N__57737),
            .I(N__57436));
    LocalMux I__13686 (
            .O(N__57734),
            .I(N__57433));
    LocalMux I__13685 (
            .O(N__57727),
            .I(N__57430));
    LocalMux I__13684 (
            .O(N__57724),
            .I(N__57427));
    LocalMux I__13683 (
            .O(N__57719),
            .I(N__57424));
    LocalMux I__13682 (
            .O(N__57716),
            .I(N__57421));
    LocalMux I__13681 (
            .O(N__57713),
            .I(N__57418));
    LocalMux I__13680 (
            .O(N__57710),
            .I(N__57415));
    LocalMux I__13679 (
            .O(N__57707),
            .I(N__57412));
    LocalMux I__13678 (
            .O(N__57704),
            .I(N__57409));
    LocalMux I__13677 (
            .O(N__57701),
            .I(N__57406));
    LocalMux I__13676 (
            .O(N__57698),
            .I(N__57403));
    LocalMux I__13675 (
            .O(N__57695),
            .I(N__57400));
    LocalMux I__13674 (
            .O(N__57690),
            .I(N__57397));
    LocalMux I__13673 (
            .O(N__57687),
            .I(N__57394));
    LocalMux I__13672 (
            .O(N__57684),
            .I(N__57391));
    LocalMux I__13671 (
            .O(N__57681),
            .I(N__57388));
    LocalMux I__13670 (
            .O(N__57678),
            .I(N__57385));
    LocalMux I__13669 (
            .O(N__57675),
            .I(N__57382));
    LocalMux I__13668 (
            .O(N__57672),
            .I(N__57379));
    LocalMux I__13667 (
            .O(N__57669),
            .I(N__57376));
    LocalMux I__13666 (
            .O(N__57666),
            .I(N__57373));
    LocalMux I__13665 (
            .O(N__57663),
            .I(N__57370));
    LocalMux I__13664 (
            .O(N__57660),
            .I(N__57367));
    LocalMux I__13663 (
            .O(N__57657),
            .I(N__57364));
    LocalMux I__13662 (
            .O(N__57654),
            .I(N__57361));
    LocalMux I__13661 (
            .O(N__57651),
            .I(N__57358));
    SRMux I__13660 (
            .O(N__57650),
            .I(N__56955));
    SRMux I__13659 (
            .O(N__57649),
            .I(N__56955));
    SRMux I__13658 (
            .O(N__57648),
            .I(N__56955));
    SRMux I__13657 (
            .O(N__57647),
            .I(N__56955));
    SRMux I__13656 (
            .O(N__57646),
            .I(N__56955));
    SRMux I__13655 (
            .O(N__57645),
            .I(N__56955));
    SRMux I__13654 (
            .O(N__57644),
            .I(N__56955));
    SRMux I__13653 (
            .O(N__57643),
            .I(N__56955));
    SRMux I__13652 (
            .O(N__57642),
            .I(N__56955));
    SRMux I__13651 (
            .O(N__57641),
            .I(N__56955));
    SRMux I__13650 (
            .O(N__57640),
            .I(N__56955));
    SRMux I__13649 (
            .O(N__57639),
            .I(N__56955));
    SRMux I__13648 (
            .O(N__57638),
            .I(N__56955));
    SRMux I__13647 (
            .O(N__57637),
            .I(N__56955));
    SRMux I__13646 (
            .O(N__57636),
            .I(N__56955));
    SRMux I__13645 (
            .O(N__57635),
            .I(N__56955));
    SRMux I__13644 (
            .O(N__57634),
            .I(N__56955));
    SRMux I__13643 (
            .O(N__57633),
            .I(N__56955));
    SRMux I__13642 (
            .O(N__57632),
            .I(N__56955));
    SRMux I__13641 (
            .O(N__57631),
            .I(N__56955));
    SRMux I__13640 (
            .O(N__57630),
            .I(N__56955));
    SRMux I__13639 (
            .O(N__57629),
            .I(N__56955));
    SRMux I__13638 (
            .O(N__57628),
            .I(N__56955));
    SRMux I__13637 (
            .O(N__57627),
            .I(N__56955));
    SRMux I__13636 (
            .O(N__57626),
            .I(N__56955));
    SRMux I__13635 (
            .O(N__57625),
            .I(N__56955));
    SRMux I__13634 (
            .O(N__57624),
            .I(N__56955));
    SRMux I__13633 (
            .O(N__57623),
            .I(N__56955));
    SRMux I__13632 (
            .O(N__57622),
            .I(N__56955));
    SRMux I__13631 (
            .O(N__57621),
            .I(N__56955));
    SRMux I__13630 (
            .O(N__57620),
            .I(N__56955));
    SRMux I__13629 (
            .O(N__57619),
            .I(N__56955));
    SRMux I__13628 (
            .O(N__57618),
            .I(N__56955));
    SRMux I__13627 (
            .O(N__57617),
            .I(N__56955));
    SRMux I__13626 (
            .O(N__57616),
            .I(N__56955));
    SRMux I__13625 (
            .O(N__57615),
            .I(N__56955));
    SRMux I__13624 (
            .O(N__57614),
            .I(N__56955));
    SRMux I__13623 (
            .O(N__57613),
            .I(N__56955));
    SRMux I__13622 (
            .O(N__57612),
            .I(N__56955));
    SRMux I__13621 (
            .O(N__57611),
            .I(N__56955));
    SRMux I__13620 (
            .O(N__57610),
            .I(N__56955));
    SRMux I__13619 (
            .O(N__57609),
            .I(N__56955));
    SRMux I__13618 (
            .O(N__57608),
            .I(N__56955));
    SRMux I__13617 (
            .O(N__57607),
            .I(N__56955));
    SRMux I__13616 (
            .O(N__57606),
            .I(N__56955));
    SRMux I__13615 (
            .O(N__57605),
            .I(N__56955));
    SRMux I__13614 (
            .O(N__57604),
            .I(N__56955));
    SRMux I__13613 (
            .O(N__57603),
            .I(N__56955));
    SRMux I__13612 (
            .O(N__57602),
            .I(N__56955));
    SRMux I__13611 (
            .O(N__57601),
            .I(N__56955));
    SRMux I__13610 (
            .O(N__57600),
            .I(N__56955));
    SRMux I__13609 (
            .O(N__57599),
            .I(N__56955));
    SRMux I__13608 (
            .O(N__57598),
            .I(N__56955));
    SRMux I__13607 (
            .O(N__57597),
            .I(N__56955));
    SRMux I__13606 (
            .O(N__57596),
            .I(N__56955));
    SRMux I__13605 (
            .O(N__57595),
            .I(N__56955));
    SRMux I__13604 (
            .O(N__57594),
            .I(N__56955));
    SRMux I__13603 (
            .O(N__57593),
            .I(N__56955));
    SRMux I__13602 (
            .O(N__57592),
            .I(N__56955));
    SRMux I__13601 (
            .O(N__57591),
            .I(N__56955));
    SRMux I__13600 (
            .O(N__57590),
            .I(N__56955));
    SRMux I__13599 (
            .O(N__57589),
            .I(N__56955));
    SRMux I__13598 (
            .O(N__57588),
            .I(N__56955));
    SRMux I__13597 (
            .O(N__57587),
            .I(N__56955));
    SRMux I__13596 (
            .O(N__57586),
            .I(N__56955));
    SRMux I__13595 (
            .O(N__57585),
            .I(N__56955));
    SRMux I__13594 (
            .O(N__57584),
            .I(N__56955));
    SRMux I__13593 (
            .O(N__57583),
            .I(N__56955));
    SRMux I__13592 (
            .O(N__57582),
            .I(N__56955));
    SRMux I__13591 (
            .O(N__57581),
            .I(N__56955));
    SRMux I__13590 (
            .O(N__57580),
            .I(N__56955));
    SRMux I__13589 (
            .O(N__57579),
            .I(N__56955));
    SRMux I__13588 (
            .O(N__57578),
            .I(N__56955));
    SRMux I__13587 (
            .O(N__57577),
            .I(N__56955));
    SRMux I__13586 (
            .O(N__57576),
            .I(N__56955));
    SRMux I__13585 (
            .O(N__57575),
            .I(N__56955));
    SRMux I__13584 (
            .O(N__57574),
            .I(N__56955));
    SRMux I__13583 (
            .O(N__57573),
            .I(N__56955));
    SRMux I__13582 (
            .O(N__57572),
            .I(N__56955));
    SRMux I__13581 (
            .O(N__57571),
            .I(N__56955));
    SRMux I__13580 (
            .O(N__57570),
            .I(N__56955));
    SRMux I__13579 (
            .O(N__57569),
            .I(N__56955));
    SRMux I__13578 (
            .O(N__57568),
            .I(N__56955));
    SRMux I__13577 (
            .O(N__57567),
            .I(N__56955));
    SRMux I__13576 (
            .O(N__57566),
            .I(N__56955));
    SRMux I__13575 (
            .O(N__57565),
            .I(N__56955));
    SRMux I__13574 (
            .O(N__57564),
            .I(N__56955));
    SRMux I__13573 (
            .O(N__57563),
            .I(N__56955));
    SRMux I__13572 (
            .O(N__57562),
            .I(N__56955));
    SRMux I__13571 (
            .O(N__57561),
            .I(N__56955));
    SRMux I__13570 (
            .O(N__57560),
            .I(N__56955));
    SRMux I__13569 (
            .O(N__57559),
            .I(N__56955));
    SRMux I__13568 (
            .O(N__57558),
            .I(N__56955));
    SRMux I__13567 (
            .O(N__57557),
            .I(N__56955));
    SRMux I__13566 (
            .O(N__57556),
            .I(N__56955));
    SRMux I__13565 (
            .O(N__57555),
            .I(N__56955));
    SRMux I__13564 (
            .O(N__57554),
            .I(N__56955));
    SRMux I__13563 (
            .O(N__57553),
            .I(N__56955));
    SRMux I__13562 (
            .O(N__57552),
            .I(N__56955));
    SRMux I__13561 (
            .O(N__57551),
            .I(N__56955));
    SRMux I__13560 (
            .O(N__57550),
            .I(N__56955));
    SRMux I__13559 (
            .O(N__57549),
            .I(N__56955));
    SRMux I__13558 (
            .O(N__57548),
            .I(N__56955));
    SRMux I__13557 (
            .O(N__57547),
            .I(N__56955));
    SRMux I__13556 (
            .O(N__57546),
            .I(N__56955));
    SRMux I__13555 (
            .O(N__57545),
            .I(N__56955));
    SRMux I__13554 (
            .O(N__57544),
            .I(N__56955));
    SRMux I__13553 (
            .O(N__57543),
            .I(N__56955));
    SRMux I__13552 (
            .O(N__57542),
            .I(N__56955));
    SRMux I__13551 (
            .O(N__57541),
            .I(N__56955));
    SRMux I__13550 (
            .O(N__57540),
            .I(N__56955));
    SRMux I__13549 (
            .O(N__57539),
            .I(N__56955));
    SRMux I__13548 (
            .O(N__57538),
            .I(N__56955));
    SRMux I__13547 (
            .O(N__57537),
            .I(N__56955));
    SRMux I__13546 (
            .O(N__57536),
            .I(N__56955));
    SRMux I__13545 (
            .O(N__57535),
            .I(N__56955));
    SRMux I__13544 (
            .O(N__57534),
            .I(N__56955));
    SRMux I__13543 (
            .O(N__57533),
            .I(N__56955));
    SRMux I__13542 (
            .O(N__57532),
            .I(N__56955));
    SRMux I__13541 (
            .O(N__57531),
            .I(N__56955));
    SRMux I__13540 (
            .O(N__57530),
            .I(N__56955));
    SRMux I__13539 (
            .O(N__57529),
            .I(N__56955));
    SRMux I__13538 (
            .O(N__57528),
            .I(N__56955));
    SRMux I__13537 (
            .O(N__57527),
            .I(N__56955));
    SRMux I__13536 (
            .O(N__57526),
            .I(N__56955));
    SRMux I__13535 (
            .O(N__57525),
            .I(N__56955));
    SRMux I__13534 (
            .O(N__57524),
            .I(N__56955));
    SRMux I__13533 (
            .O(N__57523),
            .I(N__56955));
    SRMux I__13532 (
            .O(N__57522),
            .I(N__56955));
    SRMux I__13531 (
            .O(N__57521),
            .I(N__56955));
    SRMux I__13530 (
            .O(N__57520),
            .I(N__56955));
    SRMux I__13529 (
            .O(N__57519),
            .I(N__56955));
    SRMux I__13528 (
            .O(N__57518),
            .I(N__56955));
    SRMux I__13527 (
            .O(N__57517),
            .I(N__56955));
    SRMux I__13526 (
            .O(N__57516),
            .I(N__56955));
    SRMux I__13525 (
            .O(N__57515),
            .I(N__56955));
    SRMux I__13524 (
            .O(N__57514),
            .I(N__56955));
    SRMux I__13523 (
            .O(N__57513),
            .I(N__56955));
    SRMux I__13522 (
            .O(N__57512),
            .I(N__56955));
    SRMux I__13521 (
            .O(N__57511),
            .I(N__56955));
    SRMux I__13520 (
            .O(N__57510),
            .I(N__56955));
    SRMux I__13519 (
            .O(N__57509),
            .I(N__56955));
    SRMux I__13518 (
            .O(N__57508),
            .I(N__56955));
    SRMux I__13517 (
            .O(N__57507),
            .I(N__56955));
    SRMux I__13516 (
            .O(N__57506),
            .I(N__56955));
    SRMux I__13515 (
            .O(N__57505),
            .I(N__56955));
    SRMux I__13514 (
            .O(N__57504),
            .I(N__56955));
    SRMux I__13513 (
            .O(N__57503),
            .I(N__56955));
    SRMux I__13512 (
            .O(N__57502),
            .I(N__56955));
    SRMux I__13511 (
            .O(N__57501),
            .I(N__56955));
    SRMux I__13510 (
            .O(N__57500),
            .I(N__56955));
    SRMux I__13509 (
            .O(N__57499),
            .I(N__56955));
    SRMux I__13508 (
            .O(N__57498),
            .I(N__56955));
    SRMux I__13507 (
            .O(N__57497),
            .I(N__56955));
    SRMux I__13506 (
            .O(N__57496),
            .I(N__56955));
    Glb2LocalMux I__13505 (
            .O(N__57493),
            .I(N__56955));
    Glb2LocalMux I__13504 (
            .O(N__57490),
            .I(N__56955));
    Glb2LocalMux I__13503 (
            .O(N__57487),
            .I(N__56955));
    Glb2LocalMux I__13502 (
            .O(N__57484),
            .I(N__56955));
    Glb2LocalMux I__13501 (
            .O(N__57481),
            .I(N__56955));
    Glb2LocalMux I__13500 (
            .O(N__57478),
            .I(N__56955));
    Glb2LocalMux I__13499 (
            .O(N__57475),
            .I(N__56955));
    Glb2LocalMux I__13498 (
            .O(N__57472),
            .I(N__56955));
    Glb2LocalMux I__13497 (
            .O(N__57469),
            .I(N__56955));
    Glb2LocalMux I__13496 (
            .O(N__57466),
            .I(N__56955));
    Glb2LocalMux I__13495 (
            .O(N__57463),
            .I(N__56955));
    Glb2LocalMux I__13494 (
            .O(N__57460),
            .I(N__56955));
    Glb2LocalMux I__13493 (
            .O(N__57457),
            .I(N__56955));
    Glb2LocalMux I__13492 (
            .O(N__57454),
            .I(N__56955));
    Glb2LocalMux I__13491 (
            .O(N__57451),
            .I(N__56955));
    Glb2LocalMux I__13490 (
            .O(N__57448),
            .I(N__56955));
    Glb2LocalMux I__13489 (
            .O(N__57445),
            .I(N__56955));
    Glb2LocalMux I__13488 (
            .O(N__57442),
            .I(N__56955));
    Glb2LocalMux I__13487 (
            .O(N__57439),
            .I(N__56955));
    Glb2LocalMux I__13486 (
            .O(N__57436),
            .I(N__56955));
    Glb2LocalMux I__13485 (
            .O(N__57433),
            .I(N__56955));
    Glb2LocalMux I__13484 (
            .O(N__57430),
            .I(N__56955));
    Glb2LocalMux I__13483 (
            .O(N__57427),
            .I(N__56955));
    Glb2LocalMux I__13482 (
            .O(N__57424),
            .I(N__56955));
    Glb2LocalMux I__13481 (
            .O(N__57421),
            .I(N__56955));
    Glb2LocalMux I__13480 (
            .O(N__57418),
            .I(N__56955));
    Glb2LocalMux I__13479 (
            .O(N__57415),
            .I(N__56955));
    Glb2LocalMux I__13478 (
            .O(N__57412),
            .I(N__56955));
    Glb2LocalMux I__13477 (
            .O(N__57409),
            .I(N__56955));
    Glb2LocalMux I__13476 (
            .O(N__57406),
            .I(N__56955));
    Glb2LocalMux I__13475 (
            .O(N__57403),
            .I(N__56955));
    Glb2LocalMux I__13474 (
            .O(N__57400),
            .I(N__56955));
    Glb2LocalMux I__13473 (
            .O(N__57397),
            .I(N__56955));
    Glb2LocalMux I__13472 (
            .O(N__57394),
            .I(N__56955));
    Glb2LocalMux I__13471 (
            .O(N__57391),
            .I(N__56955));
    Glb2LocalMux I__13470 (
            .O(N__57388),
            .I(N__56955));
    Glb2LocalMux I__13469 (
            .O(N__57385),
            .I(N__56955));
    Glb2LocalMux I__13468 (
            .O(N__57382),
            .I(N__56955));
    Glb2LocalMux I__13467 (
            .O(N__57379),
            .I(N__56955));
    Glb2LocalMux I__13466 (
            .O(N__57376),
            .I(N__56955));
    Glb2LocalMux I__13465 (
            .O(N__57373),
            .I(N__56955));
    Glb2LocalMux I__13464 (
            .O(N__57370),
            .I(N__56955));
    Glb2LocalMux I__13463 (
            .O(N__57367),
            .I(N__56955));
    Glb2LocalMux I__13462 (
            .O(N__57364),
            .I(N__56955));
    Glb2LocalMux I__13461 (
            .O(N__57361),
            .I(N__56955));
    Glb2LocalMux I__13460 (
            .O(N__57358),
            .I(N__56955));
    GlobalMux I__13459 (
            .O(N__56955),
            .I(N__56952));
    gio2CtrlBuf I__13458 (
            .O(N__56952),
            .I(reset_system_g));
    InMux I__13457 (
            .O(N__56949),
            .I(N__56946));
    LocalMux I__13456 (
            .O(N__56946),
            .I(N__56943));
    Odrv4 I__13455 (
            .O(N__56943),
            .I(\pid_front.O_4 ));
    CascadeMux I__13454 (
            .O(N__56940),
            .I(N__56936));
    CascadeMux I__13453 (
            .O(N__56939),
            .I(N__56932));
    InMux I__13452 (
            .O(N__56936),
            .I(N__56929));
    InMux I__13451 (
            .O(N__56935),
            .I(N__56926));
    InMux I__13450 (
            .O(N__56932),
            .I(N__56923));
    LocalMux I__13449 (
            .O(N__56929),
            .I(N__56920));
    LocalMux I__13448 (
            .O(N__56926),
            .I(N__56915));
    LocalMux I__13447 (
            .O(N__56923),
            .I(N__56915));
    Span4Mux_v I__13446 (
            .O(N__56920),
            .I(N__56912));
    Sp12to4 I__13445 (
            .O(N__56915),
            .I(N__56909));
    Sp12to4 I__13444 (
            .O(N__56912),
            .I(N__56904));
    Span12Mux_h I__13443 (
            .O(N__56909),
            .I(N__56904));
    Odrv12 I__13442 (
            .O(N__56904),
            .I(\pid_front.error_d_regZ0Z_0 ));
    InMux I__13441 (
            .O(N__56901),
            .I(N__56898));
    LocalMux I__13440 (
            .O(N__56898),
            .I(\pid_front.O_5 ));
    InMux I__13439 (
            .O(N__56895),
            .I(N__56890));
    InMux I__13438 (
            .O(N__56894),
            .I(N__56887));
    CascadeMux I__13437 (
            .O(N__56893),
            .I(N__56884));
    LocalMux I__13436 (
            .O(N__56890),
            .I(N__56881));
    LocalMux I__13435 (
            .O(N__56887),
            .I(N__56878));
    InMux I__13434 (
            .O(N__56884),
            .I(N__56875));
    Span4Mux_v I__13433 (
            .O(N__56881),
            .I(N__56868));
    Span4Mux_v I__13432 (
            .O(N__56878),
            .I(N__56868));
    LocalMux I__13431 (
            .O(N__56875),
            .I(N__56868));
    Sp12to4 I__13430 (
            .O(N__56868),
            .I(N__56865));
    Span12Mux_h I__13429 (
            .O(N__56865),
            .I(N__56862));
    Odrv12 I__13428 (
            .O(N__56862),
            .I(\pid_front.error_d_regZ0Z_1 ));
    InMux I__13427 (
            .O(N__56859),
            .I(N__56856));
    LocalMux I__13426 (
            .O(N__56856),
            .I(N__56853));
    Odrv4 I__13425 (
            .O(N__56853),
            .I(\pid_front.O_17 ));
    InMux I__13424 (
            .O(N__56850),
            .I(N__56841));
    InMux I__13423 (
            .O(N__56849),
            .I(N__56841));
    InMux I__13422 (
            .O(N__56848),
            .I(N__56841));
    LocalMux I__13421 (
            .O(N__56841),
            .I(N__56838));
    Span12Mux_h I__13420 (
            .O(N__56838),
            .I(N__56835));
    Odrv12 I__13419 (
            .O(N__56835),
            .I(\pid_front.error_d_regZ0Z_13 ));
    InMux I__13418 (
            .O(N__56832),
            .I(N__56829));
    LocalMux I__13417 (
            .O(N__56829),
            .I(N__56826));
    Odrv4 I__13416 (
            .O(N__56826),
            .I(\pid_front.O_15 ));
    InMux I__13415 (
            .O(N__56823),
            .I(N__56819));
    InMux I__13414 (
            .O(N__56822),
            .I(N__56816));
    LocalMux I__13413 (
            .O(N__56819),
            .I(N__56812));
    LocalMux I__13412 (
            .O(N__56816),
            .I(N__56809));
    InMux I__13411 (
            .O(N__56815),
            .I(N__56806));
    Span4Mux_v I__13410 (
            .O(N__56812),
            .I(N__56803));
    Span4Mux_v I__13409 (
            .O(N__56809),
            .I(N__56800));
    LocalMux I__13408 (
            .O(N__56806),
            .I(N__56797));
    Span4Mux_h I__13407 (
            .O(N__56803),
            .I(N__56794));
    Sp12to4 I__13406 (
            .O(N__56800),
            .I(N__56787));
    Span12Mux_h I__13405 (
            .O(N__56797),
            .I(N__56787));
    Sp12to4 I__13404 (
            .O(N__56794),
            .I(N__56787));
    Odrv12 I__13403 (
            .O(N__56787),
            .I(\pid_front.error_d_regZ0Z_11 ));
    InMux I__13402 (
            .O(N__56784),
            .I(N__56781));
    LocalMux I__13401 (
            .O(N__56781),
            .I(N__56778));
    Odrv4 I__13400 (
            .O(N__56778),
            .I(\pid_front.O_13 ));
    CascadeMux I__13399 (
            .O(N__56775),
            .I(N__56770));
    InMux I__13398 (
            .O(N__56774),
            .I(N__56765));
    InMux I__13397 (
            .O(N__56773),
            .I(N__56765));
    InMux I__13396 (
            .O(N__56770),
            .I(N__56762));
    LocalMux I__13395 (
            .O(N__56765),
            .I(N__56759));
    LocalMux I__13394 (
            .O(N__56762),
            .I(N__56756));
    Span4Mux_v I__13393 (
            .O(N__56759),
            .I(N__56753));
    Span12Mux_h I__13392 (
            .O(N__56756),
            .I(N__56750));
    Span4Mux_h I__13391 (
            .O(N__56753),
            .I(N__56747));
    Span12Mux_h I__13390 (
            .O(N__56750),
            .I(N__56744));
    Sp12to4 I__13389 (
            .O(N__56747),
            .I(N__56741));
    Odrv12 I__13388 (
            .O(N__56744),
            .I(\pid_front.error_d_regZ0Z_9 ));
    Odrv12 I__13387 (
            .O(N__56741),
            .I(\pid_front.error_d_regZ0Z_9 ));
    InMux I__13386 (
            .O(N__56736),
            .I(N__56733));
    LocalMux I__13385 (
            .O(N__56733),
            .I(N__56730));
    Odrv4 I__13384 (
            .O(N__56730),
            .I(\pid_front.O_20 ));
    InMux I__13383 (
            .O(N__56727),
            .I(N__56724));
    LocalMux I__13382 (
            .O(N__56724),
            .I(N__56720));
    InMux I__13381 (
            .O(N__56723),
            .I(N__56717));
    Span4Mux_h I__13380 (
            .O(N__56720),
            .I(N__56714));
    LocalMux I__13379 (
            .O(N__56717),
            .I(N__56711));
    Span4Mux_v I__13378 (
            .O(N__56714),
            .I(N__56705));
    Span4Mux_h I__13377 (
            .O(N__56711),
            .I(N__56705));
    InMux I__13376 (
            .O(N__56710),
            .I(N__56702));
    Span4Mux_h I__13375 (
            .O(N__56705),
            .I(N__56699));
    LocalMux I__13374 (
            .O(N__56702),
            .I(N__56696));
    Span4Mux_h I__13373 (
            .O(N__56699),
            .I(N__56693));
    Span12Mux_h I__13372 (
            .O(N__56696),
            .I(N__56690));
    Span4Mux_h I__13371 (
            .O(N__56693),
            .I(N__56687));
    Odrv12 I__13370 (
            .O(N__56690),
            .I(\pid_front.error_d_regZ0Z_16 ));
    Odrv4 I__13369 (
            .O(N__56687),
            .I(\pid_front.error_d_regZ0Z_16 ));
    InMux I__13368 (
            .O(N__56682),
            .I(N__56679));
    LocalMux I__13367 (
            .O(N__56679),
            .I(N__56676));
    Odrv4 I__13366 (
            .O(N__56676),
            .I(\pid_front.O_21 ));
    InMux I__13365 (
            .O(N__56673),
            .I(N__56664));
    InMux I__13364 (
            .O(N__56672),
            .I(N__56664));
    InMux I__13363 (
            .O(N__56671),
            .I(N__56664));
    LocalMux I__13362 (
            .O(N__56664),
            .I(N__56661));
    Span4Mux_h I__13361 (
            .O(N__56661),
            .I(N__56658));
    Span4Mux_h I__13360 (
            .O(N__56658),
            .I(N__56655));
    Span4Mux_h I__13359 (
            .O(N__56655),
            .I(N__56652));
    Odrv4 I__13358 (
            .O(N__56652),
            .I(\pid_front.error_d_regZ0Z_17 ));
    InMux I__13357 (
            .O(N__56649),
            .I(N__56640));
    InMux I__13356 (
            .O(N__56648),
            .I(N__56640));
    InMux I__13355 (
            .O(N__56647),
            .I(N__56640));
    LocalMux I__13354 (
            .O(N__56640),
            .I(N__56637));
    Odrv12 I__13353 (
            .O(N__56637),
            .I(\pid_side.error_d_regZ0Z_7 ));
    InMux I__13352 (
            .O(N__56634),
            .I(N__56631));
    LocalMux I__13351 (
            .O(N__56631),
            .I(\pid_side.O_1_20 ));
    InMux I__13350 (
            .O(N__56628),
            .I(N__56619));
    InMux I__13349 (
            .O(N__56627),
            .I(N__56619));
    InMux I__13348 (
            .O(N__56626),
            .I(N__56619));
    LocalMux I__13347 (
            .O(N__56619),
            .I(N__56616));
    Span4Mux_v I__13346 (
            .O(N__56616),
            .I(N__56613));
    Odrv4 I__13345 (
            .O(N__56613),
            .I(\pid_side.error_d_regZ0Z_16 ));
    CEMux I__13344 (
            .O(N__56610),
            .I(N__56604));
    CEMux I__13343 (
            .O(N__56609),
            .I(N__56600));
    CEMux I__13342 (
            .O(N__56608),
            .I(N__56594));
    CEMux I__13341 (
            .O(N__56607),
            .I(N__56589));
    LocalMux I__13340 (
            .O(N__56604),
            .I(N__56586));
    CEMux I__13339 (
            .O(N__56603),
            .I(N__56583));
    LocalMux I__13338 (
            .O(N__56600),
            .I(N__56580));
    CEMux I__13337 (
            .O(N__56599),
            .I(N__56577));
    CEMux I__13336 (
            .O(N__56598),
            .I(N__56574));
    CEMux I__13335 (
            .O(N__56597),
            .I(N__56571));
    LocalMux I__13334 (
            .O(N__56594),
            .I(N__56568));
    CEMux I__13333 (
            .O(N__56593),
            .I(N__56565));
    CEMux I__13332 (
            .O(N__56592),
            .I(N__56561));
    LocalMux I__13331 (
            .O(N__56589),
            .I(N__56558));
    Span4Mux_v I__13330 (
            .O(N__56586),
            .I(N__56553));
    LocalMux I__13329 (
            .O(N__56583),
            .I(N__56553));
    Span4Mux_v I__13328 (
            .O(N__56580),
            .I(N__56544));
    LocalMux I__13327 (
            .O(N__56577),
            .I(N__56544));
    LocalMux I__13326 (
            .O(N__56574),
            .I(N__56544));
    LocalMux I__13325 (
            .O(N__56571),
            .I(N__56544));
    Span4Mux_v I__13324 (
            .O(N__56568),
            .I(N__56541));
    LocalMux I__13323 (
            .O(N__56565),
            .I(N__56538));
    CEMux I__13322 (
            .O(N__56564),
            .I(N__56535));
    LocalMux I__13321 (
            .O(N__56561),
            .I(N__56532));
    Span4Mux_v I__13320 (
            .O(N__56558),
            .I(N__56529));
    Span4Mux_v I__13319 (
            .O(N__56553),
            .I(N__56522));
    Span4Mux_v I__13318 (
            .O(N__56544),
            .I(N__56522));
    Span4Mux_s1_h I__13317 (
            .O(N__56541),
            .I(N__56522));
    Span4Mux_v I__13316 (
            .O(N__56538),
            .I(N__56515));
    LocalMux I__13315 (
            .O(N__56535),
            .I(N__56515));
    Span4Mux_v I__13314 (
            .O(N__56532),
            .I(N__56515));
    Odrv4 I__13313 (
            .O(N__56529),
            .I(\pid_side.N_599_0 ));
    Odrv4 I__13312 (
            .O(N__56522),
            .I(\pid_side.N_599_0 ));
    Odrv4 I__13311 (
            .O(N__56515),
            .I(\pid_side.N_599_0 ));
    InMux I__13310 (
            .O(N__56508),
            .I(N__56503));
    InMux I__13309 (
            .O(N__56507),
            .I(N__56500));
    InMux I__13308 (
            .O(N__56506),
            .I(N__56497));
    LocalMux I__13307 (
            .O(N__56503),
            .I(N__56494));
    LocalMux I__13306 (
            .O(N__56500),
            .I(N__56491));
    LocalMux I__13305 (
            .O(N__56497),
            .I(N__56488));
    Span4Mux_s3_h I__13304 (
            .O(N__56494),
            .I(N__56483));
    Span4Mux_v I__13303 (
            .O(N__56491),
            .I(N__56480));
    Span4Mux_v I__13302 (
            .O(N__56488),
            .I(N__56476));
    InMux I__13301 (
            .O(N__56487),
            .I(N__56473));
    InMux I__13300 (
            .O(N__56486),
            .I(N__56470));
    Span4Mux_h I__13299 (
            .O(N__56483),
            .I(N__56467));
    Span4Mux_h I__13298 (
            .O(N__56480),
            .I(N__56461));
    InMux I__13297 (
            .O(N__56479),
            .I(N__56458));
    Span4Mux_h I__13296 (
            .O(N__56476),
            .I(N__56455));
    LocalMux I__13295 (
            .O(N__56473),
            .I(N__56451));
    LocalMux I__13294 (
            .O(N__56470),
            .I(N__56448));
    Span4Mux_h I__13293 (
            .O(N__56467),
            .I(N__56445));
    InMux I__13292 (
            .O(N__56466),
            .I(N__56442));
    InMux I__13291 (
            .O(N__56465),
            .I(N__56437));
    InMux I__13290 (
            .O(N__56464),
            .I(N__56434));
    Span4Mux_v I__13289 (
            .O(N__56461),
            .I(N__56428));
    LocalMux I__13288 (
            .O(N__56458),
            .I(N__56428));
    Span4Mux_v I__13287 (
            .O(N__56455),
            .I(N__56425));
    InMux I__13286 (
            .O(N__56454),
            .I(N__56422));
    Span4Mux_v I__13285 (
            .O(N__56451),
            .I(N__56417));
    Span4Mux_s3_h I__13284 (
            .O(N__56448),
            .I(N__56417));
    Span4Mux_h I__13283 (
            .O(N__56445),
            .I(N__56412));
    LocalMux I__13282 (
            .O(N__56442),
            .I(N__56412));
    CascadeMux I__13281 (
            .O(N__56441),
            .I(N__56409));
    InMux I__13280 (
            .O(N__56440),
            .I(N__56406));
    LocalMux I__13279 (
            .O(N__56437),
            .I(N__56403));
    LocalMux I__13278 (
            .O(N__56434),
            .I(N__56400));
    InMux I__13277 (
            .O(N__56433),
            .I(N__56397));
    Span4Mux_h I__13276 (
            .O(N__56428),
            .I(N__56394));
    Span4Mux_v I__13275 (
            .O(N__56425),
            .I(N__56389));
    LocalMux I__13274 (
            .O(N__56422),
            .I(N__56389));
    Span4Mux_h I__13273 (
            .O(N__56417),
            .I(N__56385));
    Span4Mux_v I__13272 (
            .O(N__56412),
            .I(N__56381));
    InMux I__13271 (
            .O(N__56409),
            .I(N__56378));
    LocalMux I__13270 (
            .O(N__56406),
            .I(N__56375));
    Span4Mux_v I__13269 (
            .O(N__56403),
            .I(N__56368));
    Span4Mux_v I__13268 (
            .O(N__56400),
            .I(N__56368));
    LocalMux I__13267 (
            .O(N__56397),
            .I(N__56368));
    Span4Mux_h I__13266 (
            .O(N__56394),
            .I(N__56363));
    Span4Mux_v I__13265 (
            .O(N__56389),
            .I(N__56363));
    InMux I__13264 (
            .O(N__56388),
            .I(N__56360));
    Sp12to4 I__13263 (
            .O(N__56385),
            .I(N__56357));
    InMux I__13262 (
            .O(N__56384),
            .I(N__56354));
    Span4Mux_v I__13261 (
            .O(N__56381),
            .I(N__56345));
    LocalMux I__13260 (
            .O(N__56378),
            .I(N__56345));
    Span4Mux_v I__13259 (
            .O(N__56375),
            .I(N__56345));
    Span4Mux_h I__13258 (
            .O(N__56368),
            .I(N__56345));
    Odrv4 I__13257 (
            .O(N__56363),
            .I(uart_pc_data_0));
    LocalMux I__13256 (
            .O(N__56360),
            .I(uart_pc_data_0));
    Odrv12 I__13255 (
            .O(N__56357),
            .I(uart_pc_data_0));
    LocalMux I__13254 (
            .O(N__56354),
            .I(uart_pc_data_0));
    Odrv4 I__13253 (
            .O(N__56345),
            .I(uart_pc_data_0));
    InMux I__13252 (
            .O(N__56334),
            .I(N__56331));
    LocalMux I__13251 (
            .O(N__56331),
            .I(N__56328));
    Span4Mux_v I__13250 (
            .O(N__56328),
            .I(N__56325));
    Span4Mux_v I__13249 (
            .O(N__56325),
            .I(N__56321));
    InMux I__13248 (
            .O(N__56324),
            .I(N__56318));
    Odrv4 I__13247 (
            .O(N__56321),
            .I(xy_kd_0));
    LocalMux I__13246 (
            .O(N__56318),
            .I(xy_kd_0));
    InMux I__13245 (
            .O(N__56313),
            .I(N__56308));
    InMux I__13244 (
            .O(N__56312),
            .I(N__56305));
    InMux I__13243 (
            .O(N__56311),
            .I(N__56301));
    LocalMux I__13242 (
            .O(N__56308),
            .I(N__56298));
    LocalMux I__13241 (
            .O(N__56305),
            .I(N__56295));
    InMux I__13240 (
            .O(N__56304),
            .I(N__56292));
    LocalMux I__13239 (
            .O(N__56301),
            .I(N__56289));
    Span4Mux_h I__13238 (
            .O(N__56298),
            .I(N__56286));
    Span4Mux_h I__13237 (
            .O(N__56295),
            .I(N__56279));
    LocalMux I__13236 (
            .O(N__56292),
            .I(N__56279));
    Span4Mux_v I__13235 (
            .O(N__56289),
            .I(N__56275));
    Span4Mux_h I__13234 (
            .O(N__56286),
            .I(N__56272));
    InMux I__13233 (
            .O(N__56285),
            .I(N__56267));
    InMux I__13232 (
            .O(N__56284),
            .I(N__56263));
    Span4Mux_v I__13231 (
            .O(N__56279),
            .I(N__56260));
    InMux I__13230 (
            .O(N__56278),
            .I(N__56257));
    Span4Mux_v I__13229 (
            .O(N__56275),
            .I(N__56252));
    Span4Mux_h I__13228 (
            .O(N__56272),
            .I(N__56252));
    InMux I__13227 (
            .O(N__56271),
            .I(N__56249));
    InMux I__13226 (
            .O(N__56270),
            .I(N__56246));
    LocalMux I__13225 (
            .O(N__56267),
            .I(N__56243));
    InMux I__13224 (
            .O(N__56266),
            .I(N__56239));
    LocalMux I__13223 (
            .O(N__56263),
            .I(N__56236));
    Span4Mux_v I__13222 (
            .O(N__56260),
            .I(N__56233));
    LocalMux I__13221 (
            .O(N__56257),
            .I(N__56230));
    Span4Mux_h I__13220 (
            .O(N__56252),
            .I(N__56225));
    LocalMux I__13219 (
            .O(N__56249),
            .I(N__56225));
    LocalMux I__13218 (
            .O(N__56246),
            .I(N__56221));
    Span12Mux_v I__13217 (
            .O(N__56243),
            .I(N__56217));
    InMux I__13216 (
            .O(N__56242),
            .I(N__56214));
    LocalMux I__13215 (
            .O(N__56239),
            .I(N__56211));
    Span4Mux_v I__13214 (
            .O(N__56236),
            .I(N__56208));
    Span4Mux_v I__13213 (
            .O(N__56233),
            .I(N__56203));
    Span4Mux_v I__13212 (
            .O(N__56230),
            .I(N__56203));
    Span4Mux_v I__13211 (
            .O(N__56225),
            .I(N__56200));
    InMux I__13210 (
            .O(N__56224),
            .I(N__56197));
    Span4Mux_h I__13209 (
            .O(N__56221),
            .I(N__56194));
    InMux I__13208 (
            .O(N__56220),
            .I(N__56191));
    Span12Mux_h I__13207 (
            .O(N__56217),
            .I(N__56186));
    LocalMux I__13206 (
            .O(N__56214),
            .I(N__56186));
    Span4Mux_h I__13205 (
            .O(N__56211),
            .I(N__56183));
    Span4Mux_h I__13204 (
            .O(N__56208),
            .I(N__56174));
    Span4Mux_h I__13203 (
            .O(N__56203),
            .I(N__56174));
    Span4Mux_v I__13202 (
            .O(N__56200),
            .I(N__56174));
    LocalMux I__13201 (
            .O(N__56197),
            .I(N__56174));
    Odrv4 I__13200 (
            .O(N__56194),
            .I(uart_pc_data_1));
    LocalMux I__13199 (
            .O(N__56191),
            .I(uart_pc_data_1));
    Odrv12 I__13198 (
            .O(N__56186),
            .I(uart_pc_data_1));
    Odrv4 I__13197 (
            .O(N__56183),
            .I(uart_pc_data_1));
    Odrv4 I__13196 (
            .O(N__56174),
            .I(uart_pc_data_1));
    InMux I__13195 (
            .O(N__56163),
            .I(N__56160));
    LocalMux I__13194 (
            .O(N__56160),
            .I(N__56157));
    Span4Mux_v I__13193 (
            .O(N__56157),
            .I(N__56154));
    Span4Mux_v I__13192 (
            .O(N__56154),
            .I(N__56150));
    InMux I__13191 (
            .O(N__56153),
            .I(N__56147));
    Odrv4 I__13190 (
            .O(N__56150),
            .I(xy_kd_1));
    LocalMux I__13189 (
            .O(N__56147),
            .I(xy_kd_1));
    InMux I__13188 (
            .O(N__56142),
            .I(N__56136));
    InMux I__13187 (
            .O(N__56141),
            .I(N__56133));
    InMux I__13186 (
            .O(N__56140),
            .I(N__56129));
    InMux I__13185 (
            .O(N__56139),
            .I(N__56126));
    LocalMux I__13184 (
            .O(N__56136),
            .I(N__56121));
    LocalMux I__13183 (
            .O(N__56133),
            .I(N__56118));
    InMux I__13182 (
            .O(N__56132),
            .I(N__56115));
    LocalMux I__13181 (
            .O(N__56129),
            .I(N__56112));
    LocalMux I__13180 (
            .O(N__56126),
            .I(N__56107));
    InMux I__13179 (
            .O(N__56125),
            .I(N__56102));
    InMux I__13178 (
            .O(N__56124),
            .I(N__56099));
    Span4Mux_v I__13177 (
            .O(N__56121),
            .I(N__56096));
    Span4Mux_v I__13176 (
            .O(N__56118),
            .I(N__56093));
    LocalMux I__13175 (
            .O(N__56115),
            .I(N__56090));
    Span4Mux_v I__13174 (
            .O(N__56112),
            .I(N__56087));
    InMux I__13173 (
            .O(N__56111),
            .I(N__56084));
    InMux I__13172 (
            .O(N__56110),
            .I(N__56081));
    Span4Mux_v I__13171 (
            .O(N__56107),
            .I(N__56078));
    CascadeMux I__13170 (
            .O(N__56106),
            .I(N__56075));
    InMux I__13169 (
            .O(N__56105),
            .I(N__56070));
    LocalMux I__13168 (
            .O(N__56102),
            .I(N__56067));
    LocalMux I__13167 (
            .O(N__56099),
            .I(N__56064));
    Sp12to4 I__13166 (
            .O(N__56096),
            .I(N__56061));
    Sp12to4 I__13165 (
            .O(N__56093),
            .I(N__56058));
    Span4Mux_v I__13164 (
            .O(N__56090),
            .I(N__56053));
    Span4Mux_h I__13163 (
            .O(N__56087),
            .I(N__56053));
    LocalMux I__13162 (
            .O(N__56084),
            .I(N__56050));
    LocalMux I__13161 (
            .O(N__56081),
            .I(N__56047));
    Span4Mux_h I__13160 (
            .O(N__56078),
            .I(N__56043));
    InMux I__13159 (
            .O(N__56075),
            .I(N__56040));
    InMux I__13158 (
            .O(N__56074),
            .I(N__56037));
    CascadeMux I__13157 (
            .O(N__56073),
            .I(N__56034));
    LocalMux I__13156 (
            .O(N__56070),
            .I(N__56031));
    Span4Mux_v I__13155 (
            .O(N__56067),
            .I(N__56028));
    Span4Mux_v I__13154 (
            .O(N__56064),
            .I(N__56025));
    Span12Mux_h I__13153 (
            .O(N__56061),
            .I(N__56020));
    Span12Mux_s6_h I__13152 (
            .O(N__56058),
            .I(N__56020));
    Span4Mux_v I__13151 (
            .O(N__56053),
            .I(N__56017));
    Span4Mux_v I__13150 (
            .O(N__56050),
            .I(N__56013));
    Span4Mux_v I__13149 (
            .O(N__56047),
            .I(N__56010));
    InMux I__13148 (
            .O(N__56046),
            .I(N__56007));
    Span4Mux_v I__13147 (
            .O(N__56043),
            .I(N__56002));
    LocalMux I__13146 (
            .O(N__56040),
            .I(N__56002));
    LocalMux I__13145 (
            .O(N__56037),
            .I(N__55998));
    InMux I__13144 (
            .O(N__56034),
            .I(N__55995));
    Span4Mux_v I__13143 (
            .O(N__56031),
            .I(N__55990));
    Span4Mux_h I__13142 (
            .O(N__56028),
            .I(N__55990));
    Sp12to4 I__13141 (
            .O(N__56025),
            .I(N__55983));
    Span12Mux_v I__13140 (
            .O(N__56020),
            .I(N__55983));
    Sp12to4 I__13139 (
            .O(N__56017),
            .I(N__55983));
    InMux I__13138 (
            .O(N__56016),
            .I(N__55980));
    Span4Mux_h I__13137 (
            .O(N__56013),
            .I(N__55971));
    Span4Mux_v I__13136 (
            .O(N__56010),
            .I(N__55971));
    LocalMux I__13135 (
            .O(N__56007),
            .I(N__55971));
    Span4Mux_v I__13134 (
            .O(N__56002),
            .I(N__55971));
    InMux I__13133 (
            .O(N__56001),
            .I(N__55968));
    Span4Mux_v I__13132 (
            .O(N__55998),
            .I(N__55965));
    LocalMux I__13131 (
            .O(N__55995),
            .I(uart_pc_data_2));
    Odrv4 I__13130 (
            .O(N__55990),
            .I(uart_pc_data_2));
    Odrv12 I__13129 (
            .O(N__55983),
            .I(uart_pc_data_2));
    LocalMux I__13128 (
            .O(N__55980),
            .I(uart_pc_data_2));
    Odrv4 I__13127 (
            .O(N__55971),
            .I(uart_pc_data_2));
    LocalMux I__13126 (
            .O(N__55968),
            .I(uart_pc_data_2));
    Odrv4 I__13125 (
            .O(N__55965),
            .I(uart_pc_data_2));
    InMux I__13124 (
            .O(N__55950),
            .I(N__55947));
    LocalMux I__13123 (
            .O(N__55947),
            .I(N__55944));
    Span4Mux_v I__13122 (
            .O(N__55944),
            .I(N__55940));
    InMux I__13121 (
            .O(N__55943),
            .I(N__55937));
    Odrv4 I__13120 (
            .O(N__55940),
            .I(xy_kd_2));
    LocalMux I__13119 (
            .O(N__55937),
            .I(xy_kd_2));
    InMux I__13118 (
            .O(N__55932),
            .I(N__55928));
    InMux I__13117 (
            .O(N__55931),
            .I(N__55923));
    LocalMux I__13116 (
            .O(N__55928),
            .I(N__55919));
    InMux I__13115 (
            .O(N__55927),
            .I(N__55916));
    InMux I__13114 (
            .O(N__55926),
            .I(N__55913));
    LocalMux I__13113 (
            .O(N__55923),
            .I(N__55910));
    InMux I__13112 (
            .O(N__55922),
            .I(N__55907));
    Span4Mux_v I__13111 (
            .O(N__55919),
            .I(N__55904));
    LocalMux I__13110 (
            .O(N__55916),
            .I(N__55900));
    LocalMux I__13109 (
            .O(N__55913),
            .I(N__55895));
    Span4Mux_s1_h I__13108 (
            .O(N__55910),
            .I(N__55892));
    LocalMux I__13107 (
            .O(N__55907),
            .I(N__55889));
    Span4Mux_v I__13106 (
            .O(N__55904),
            .I(N__55886));
    InMux I__13105 (
            .O(N__55903),
            .I(N__55883));
    Span4Mux_v I__13104 (
            .O(N__55900),
            .I(N__55880));
    InMux I__13103 (
            .O(N__55899),
            .I(N__55877));
    InMux I__13102 (
            .O(N__55898),
            .I(N__55872));
    Span4Mux_v I__13101 (
            .O(N__55895),
            .I(N__55867));
    Span4Mux_h I__13100 (
            .O(N__55892),
            .I(N__55867));
    Span4Mux_h I__13099 (
            .O(N__55889),
            .I(N__55864));
    Span4Mux_v I__13098 (
            .O(N__55886),
            .I(N__55859));
    LocalMux I__13097 (
            .O(N__55883),
            .I(N__55859));
    Span4Mux_v I__13096 (
            .O(N__55880),
            .I(N__55856));
    LocalMux I__13095 (
            .O(N__55877),
            .I(N__55853));
    InMux I__13094 (
            .O(N__55876),
            .I(N__55850));
    InMux I__13093 (
            .O(N__55875),
            .I(N__55847));
    LocalMux I__13092 (
            .O(N__55872),
            .I(N__55842));
    Sp12to4 I__13091 (
            .O(N__55867),
            .I(N__55839));
    Sp12to4 I__13090 (
            .O(N__55864),
            .I(N__55836));
    Span4Mux_v I__13089 (
            .O(N__55859),
            .I(N__55832));
    Span4Mux_v I__13088 (
            .O(N__55856),
            .I(N__55825));
    Span4Mux_v I__13087 (
            .O(N__55853),
            .I(N__55825));
    LocalMux I__13086 (
            .O(N__55850),
            .I(N__55825));
    LocalMux I__13085 (
            .O(N__55847),
            .I(N__55822));
    InMux I__13084 (
            .O(N__55846),
            .I(N__55819));
    InMux I__13083 (
            .O(N__55845),
            .I(N__55814));
    Span4Mux_v I__13082 (
            .O(N__55842),
            .I(N__55811));
    Span12Mux_h I__13081 (
            .O(N__55839),
            .I(N__55806));
    Span12Mux_v I__13080 (
            .O(N__55836),
            .I(N__55806));
    InMux I__13079 (
            .O(N__55835),
            .I(N__55803));
    Span4Mux_h I__13078 (
            .O(N__55832),
            .I(N__55794));
    Span4Mux_h I__13077 (
            .O(N__55825),
            .I(N__55794));
    Span4Mux_v I__13076 (
            .O(N__55822),
            .I(N__55794));
    LocalMux I__13075 (
            .O(N__55819),
            .I(N__55794));
    InMux I__13074 (
            .O(N__55818),
            .I(N__55789));
    InMux I__13073 (
            .O(N__55817),
            .I(N__55789));
    LocalMux I__13072 (
            .O(N__55814),
            .I(N__55786));
    Odrv4 I__13071 (
            .O(N__55811),
            .I(uart_pc_data_5));
    Odrv12 I__13070 (
            .O(N__55806),
            .I(uart_pc_data_5));
    LocalMux I__13069 (
            .O(N__55803),
            .I(uart_pc_data_5));
    Odrv4 I__13068 (
            .O(N__55794),
            .I(uart_pc_data_5));
    LocalMux I__13067 (
            .O(N__55789),
            .I(uart_pc_data_5));
    Odrv4 I__13066 (
            .O(N__55786),
            .I(uart_pc_data_5));
    InMux I__13065 (
            .O(N__55773),
            .I(N__55770));
    LocalMux I__13064 (
            .O(N__55770),
            .I(N__55767));
    Span4Mux_v I__13063 (
            .O(N__55767),
            .I(N__55763));
    InMux I__13062 (
            .O(N__55766),
            .I(N__55760));
    Odrv4 I__13061 (
            .O(N__55763),
            .I(xy_kd_5));
    LocalMux I__13060 (
            .O(N__55760),
            .I(xy_kd_5));
    InMux I__13059 (
            .O(N__55755),
            .I(N__55751));
    InMux I__13058 (
            .O(N__55754),
            .I(N__55746));
    LocalMux I__13057 (
            .O(N__55751),
            .I(N__55743));
    InMux I__13056 (
            .O(N__55750),
            .I(N__55740));
    InMux I__13055 (
            .O(N__55749),
            .I(N__55737));
    LocalMux I__13054 (
            .O(N__55746),
            .I(N__55734));
    Span4Mux_v I__13053 (
            .O(N__55743),
            .I(N__55727));
    LocalMux I__13052 (
            .O(N__55740),
            .I(N__55724));
    LocalMux I__13051 (
            .O(N__55737),
            .I(N__55720));
    Span4Mux_v I__13050 (
            .O(N__55734),
            .I(N__55717));
    InMux I__13049 (
            .O(N__55733),
            .I(N__55713));
    InMux I__13048 (
            .O(N__55732),
            .I(N__55710));
    InMux I__13047 (
            .O(N__55731),
            .I(N__55706));
    InMux I__13046 (
            .O(N__55730),
            .I(N__55702));
    Sp12to4 I__13045 (
            .O(N__55727),
            .I(N__55699));
    Span4Mux_v I__13044 (
            .O(N__55724),
            .I(N__55696));
    InMux I__13043 (
            .O(N__55723),
            .I(N__55693));
    Span4Mux_v I__13042 (
            .O(N__55720),
            .I(N__55688));
    Span4Mux_h I__13041 (
            .O(N__55717),
            .I(N__55688));
    InMux I__13040 (
            .O(N__55716),
            .I(N__55685));
    LocalMux I__13039 (
            .O(N__55713),
            .I(N__55682));
    LocalMux I__13038 (
            .O(N__55710),
            .I(N__55679));
    InMux I__13037 (
            .O(N__55709),
            .I(N__55676));
    LocalMux I__13036 (
            .O(N__55706),
            .I(N__55673));
    InMux I__13035 (
            .O(N__55705),
            .I(N__55670));
    LocalMux I__13034 (
            .O(N__55702),
            .I(N__55667));
    Span12Mux_h I__13033 (
            .O(N__55699),
            .I(N__55659));
    Sp12to4 I__13032 (
            .O(N__55696),
            .I(N__55659));
    LocalMux I__13031 (
            .O(N__55693),
            .I(N__55659));
    Sp12to4 I__13030 (
            .O(N__55688),
            .I(N__55656));
    LocalMux I__13029 (
            .O(N__55685),
            .I(N__55653));
    Span4Mux_v I__13028 (
            .O(N__55682),
            .I(N__55650));
    Span4Mux_v I__13027 (
            .O(N__55679),
            .I(N__55647));
    LocalMux I__13026 (
            .O(N__55676),
            .I(N__55644));
    Span4Mux_h I__13025 (
            .O(N__55673),
            .I(N__55639));
    LocalMux I__13024 (
            .O(N__55670),
            .I(N__55639));
    Span4Mux_h I__13023 (
            .O(N__55667),
            .I(N__55636));
    InMux I__13022 (
            .O(N__55666),
            .I(N__55633));
    Span12Mux_v I__13021 (
            .O(N__55659),
            .I(N__55630));
    Span12Mux_h I__13020 (
            .O(N__55656),
            .I(N__55625));
    Span12Mux_s7_h I__13019 (
            .O(N__55653),
            .I(N__55625));
    Span4Mux_h I__13018 (
            .O(N__55650),
            .I(N__55616));
    Span4Mux_h I__13017 (
            .O(N__55647),
            .I(N__55616));
    Span4Mux_v I__13016 (
            .O(N__55644),
            .I(N__55616));
    Span4Mux_v I__13015 (
            .O(N__55639),
            .I(N__55616));
    Odrv4 I__13014 (
            .O(N__55636),
            .I(uart_pc_data_6));
    LocalMux I__13013 (
            .O(N__55633),
            .I(uart_pc_data_6));
    Odrv12 I__13012 (
            .O(N__55630),
            .I(uart_pc_data_6));
    Odrv12 I__13011 (
            .O(N__55625),
            .I(uart_pc_data_6));
    Odrv4 I__13010 (
            .O(N__55616),
            .I(uart_pc_data_6));
    InMux I__13009 (
            .O(N__55605),
            .I(N__55602));
    LocalMux I__13008 (
            .O(N__55602),
            .I(N__55599));
    Span4Mux_s0_h I__13007 (
            .O(N__55599),
            .I(N__55596));
    Span4Mux_v I__13006 (
            .O(N__55596),
            .I(N__55592));
    InMux I__13005 (
            .O(N__55595),
            .I(N__55589));
    Odrv4 I__13004 (
            .O(N__55592),
            .I(xy_kd_6));
    LocalMux I__13003 (
            .O(N__55589),
            .I(xy_kd_6));
    InMux I__13002 (
            .O(N__55584),
            .I(N__55578));
    InMux I__13001 (
            .O(N__55583),
            .I(N__55575));
    InMux I__13000 (
            .O(N__55582),
            .I(N__55571));
    InMux I__12999 (
            .O(N__55581),
            .I(N__55568));
    LocalMux I__12998 (
            .O(N__55578),
            .I(N__55562));
    LocalMux I__12997 (
            .O(N__55575),
            .I(N__55559));
    InMux I__12996 (
            .O(N__55574),
            .I(N__55556));
    LocalMux I__12995 (
            .O(N__55571),
            .I(N__55553));
    LocalMux I__12994 (
            .O(N__55568),
            .I(N__55550));
    InMux I__12993 (
            .O(N__55567),
            .I(N__55545));
    InMux I__12992 (
            .O(N__55566),
            .I(N__55542));
    InMux I__12991 (
            .O(N__55565),
            .I(N__55538));
    Span4Mux_v I__12990 (
            .O(N__55562),
            .I(N__55535));
    Span4Mux_s3_h I__12989 (
            .O(N__55559),
            .I(N__55531));
    LocalMux I__12988 (
            .O(N__55556),
            .I(N__55528));
    Span4Mux_v I__12987 (
            .O(N__55553),
            .I(N__55525));
    Span4Mux_v I__12986 (
            .O(N__55550),
            .I(N__55522));
    InMux I__12985 (
            .O(N__55549),
            .I(N__55518));
    InMux I__12984 (
            .O(N__55548),
            .I(N__55515));
    LocalMux I__12983 (
            .O(N__55545),
            .I(N__55512));
    LocalMux I__12982 (
            .O(N__55542),
            .I(N__55509));
    InMux I__12981 (
            .O(N__55541),
            .I(N__55506));
    LocalMux I__12980 (
            .O(N__55538),
            .I(N__55503));
    Span4Mux_h I__12979 (
            .O(N__55535),
            .I(N__55500));
    CascadeMux I__12978 (
            .O(N__55534),
            .I(N__55497));
    Span4Mux_h I__12977 (
            .O(N__55531),
            .I(N__55494));
    Span4Mux_v I__12976 (
            .O(N__55528),
            .I(N__55489));
    Span4Mux_h I__12975 (
            .O(N__55525),
            .I(N__55489));
    Span4Mux_h I__12974 (
            .O(N__55522),
            .I(N__55486));
    InMux I__12973 (
            .O(N__55521),
            .I(N__55483));
    LocalMux I__12972 (
            .O(N__55518),
            .I(N__55480));
    LocalMux I__12971 (
            .O(N__55515),
            .I(N__55477));
    Span4Mux_v I__12970 (
            .O(N__55512),
            .I(N__55474));
    Span4Mux_v I__12969 (
            .O(N__55509),
            .I(N__55471));
    LocalMux I__12968 (
            .O(N__55506),
            .I(N__55468));
    Span4Mux_s3_h I__12967 (
            .O(N__55503),
            .I(N__55465));
    Span4Mux_v I__12966 (
            .O(N__55500),
            .I(N__55462));
    InMux I__12965 (
            .O(N__55497),
            .I(N__55459));
    Sp12to4 I__12964 (
            .O(N__55494),
            .I(N__55456));
    Span4Mux_v I__12963 (
            .O(N__55489),
            .I(N__55453));
    Span4Mux_v I__12962 (
            .O(N__55486),
            .I(N__55450));
    LocalMux I__12961 (
            .O(N__55483),
            .I(N__55447));
    Span4Mux_v I__12960 (
            .O(N__55480),
            .I(N__55436));
    Span4Mux_v I__12959 (
            .O(N__55477),
            .I(N__55436));
    Span4Mux_h I__12958 (
            .O(N__55474),
            .I(N__55436));
    Span4Mux_h I__12957 (
            .O(N__55471),
            .I(N__55436));
    Span4Mux_h I__12956 (
            .O(N__55468),
            .I(N__55431));
    Span4Mux_h I__12955 (
            .O(N__55465),
            .I(N__55431));
    Span4Mux_v I__12954 (
            .O(N__55462),
            .I(N__55428));
    LocalMux I__12953 (
            .O(N__55459),
            .I(N__55421));
    Span12Mux_v I__12952 (
            .O(N__55456),
            .I(N__55421));
    Sp12to4 I__12951 (
            .O(N__55453),
            .I(N__55421));
    Span4Mux_v I__12950 (
            .O(N__55450),
            .I(N__55416));
    Span4Mux_h I__12949 (
            .O(N__55447),
            .I(N__55416));
    InMux I__12948 (
            .O(N__55446),
            .I(N__55413));
    InMux I__12947 (
            .O(N__55445),
            .I(N__55410));
    Odrv4 I__12946 (
            .O(N__55436),
            .I(uart_pc_data_7));
    Odrv4 I__12945 (
            .O(N__55431),
            .I(uart_pc_data_7));
    Odrv4 I__12944 (
            .O(N__55428),
            .I(uart_pc_data_7));
    Odrv12 I__12943 (
            .O(N__55421),
            .I(uart_pc_data_7));
    Odrv4 I__12942 (
            .O(N__55416),
            .I(uart_pc_data_7));
    LocalMux I__12941 (
            .O(N__55413),
            .I(uart_pc_data_7));
    LocalMux I__12940 (
            .O(N__55410),
            .I(uart_pc_data_7));
    InMux I__12939 (
            .O(N__55395),
            .I(N__55392));
    LocalMux I__12938 (
            .O(N__55392),
            .I(N__55389));
    Span4Mux_v I__12937 (
            .O(N__55389),
            .I(N__55385));
    InMux I__12936 (
            .O(N__55388),
            .I(N__55382));
    Odrv4 I__12935 (
            .O(N__55385),
            .I(xy_kd_7));
    LocalMux I__12934 (
            .O(N__55382),
            .I(xy_kd_7));
    InMux I__12933 (
            .O(N__55377),
            .I(N__55374));
    LocalMux I__12932 (
            .O(N__55374),
            .I(N__55369));
    InMux I__12931 (
            .O(N__55373),
            .I(N__55366));
    InMux I__12930 (
            .O(N__55372),
            .I(N__55363));
    Span4Mux_v I__12929 (
            .O(N__55369),
            .I(N__55357));
    LocalMux I__12928 (
            .O(N__55366),
            .I(N__55357));
    LocalMux I__12927 (
            .O(N__55363),
            .I(N__55350));
    InMux I__12926 (
            .O(N__55362),
            .I(N__55347));
    Span4Mux_v I__12925 (
            .O(N__55357),
            .I(N__55344));
    InMux I__12924 (
            .O(N__55356),
            .I(N__55339));
    InMux I__12923 (
            .O(N__55355),
            .I(N__55336));
    InMux I__12922 (
            .O(N__55354),
            .I(N__55333));
    InMux I__12921 (
            .O(N__55353),
            .I(N__55329));
    Span4Mux_v I__12920 (
            .O(N__55350),
            .I(N__55326));
    LocalMux I__12919 (
            .O(N__55347),
            .I(N__55323));
    Span4Mux_h I__12918 (
            .O(N__55344),
            .I(N__55320));
    InMux I__12917 (
            .O(N__55343),
            .I(N__55317));
    InMux I__12916 (
            .O(N__55342),
            .I(N__55314));
    LocalMux I__12915 (
            .O(N__55339),
            .I(N__55311));
    LocalMux I__12914 (
            .O(N__55336),
            .I(N__55308));
    LocalMux I__12913 (
            .O(N__55333),
            .I(N__55305));
    InMux I__12912 (
            .O(N__55332),
            .I(N__55302));
    LocalMux I__12911 (
            .O(N__55329),
            .I(N__55299));
    Span4Mux_v I__12910 (
            .O(N__55326),
            .I(N__55296));
    Sp12to4 I__12909 (
            .O(N__55323),
            .I(N__55293));
    Span4Mux_v I__12908 (
            .O(N__55320),
            .I(N__55290));
    LocalMux I__12907 (
            .O(N__55317),
            .I(N__55285));
    LocalMux I__12906 (
            .O(N__55314),
            .I(N__55285));
    Span12Mux_h I__12905 (
            .O(N__55311),
            .I(N__55281));
    Span4Mux_v I__12904 (
            .O(N__55308),
            .I(N__55273));
    Span4Mux_s3_h I__12903 (
            .O(N__55305),
            .I(N__55273));
    LocalMux I__12902 (
            .O(N__55302),
            .I(N__55273));
    Span4Mux_v I__12901 (
            .O(N__55299),
            .I(N__55270));
    Sp12to4 I__12900 (
            .O(N__55296),
            .I(N__55265));
    Span12Mux_v I__12899 (
            .O(N__55293),
            .I(N__55265));
    Span4Mux_v I__12898 (
            .O(N__55290),
            .I(N__55260));
    Span4Mux_v I__12897 (
            .O(N__55285),
            .I(N__55260));
    InMux I__12896 (
            .O(N__55284),
            .I(N__55257));
    Span12Mux_v I__12895 (
            .O(N__55281),
            .I(N__55254));
    InMux I__12894 (
            .O(N__55280),
            .I(N__55251));
    Span4Mux_h I__12893 (
            .O(N__55273),
            .I(N__55248));
    Sp12to4 I__12892 (
            .O(N__55270),
            .I(N__55239));
    Span12Mux_h I__12891 (
            .O(N__55265),
            .I(N__55239));
    Sp12to4 I__12890 (
            .O(N__55260),
            .I(N__55239));
    LocalMux I__12889 (
            .O(N__55257),
            .I(N__55239));
    Odrv12 I__12888 (
            .O(N__55254),
            .I(uart_pc_data_3));
    LocalMux I__12887 (
            .O(N__55251),
            .I(uart_pc_data_3));
    Odrv4 I__12886 (
            .O(N__55248),
            .I(uart_pc_data_3));
    Odrv12 I__12885 (
            .O(N__55239),
            .I(uart_pc_data_3));
    InMux I__12884 (
            .O(N__55230),
            .I(N__55227));
    LocalMux I__12883 (
            .O(N__55227),
            .I(N__55224));
    Span4Mux_v I__12882 (
            .O(N__55224),
            .I(N__55220));
    InMux I__12881 (
            .O(N__55223),
            .I(N__55217));
    Odrv4 I__12880 (
            .O(N__55220),
            .I(xy_kd_3));
    LocalMux I__12879 (
            .O(N__55217),
            .I(xy_kd_3));
    CEMux I__12878 (
            .O(N__55212),
            .I(N__55209));
    LocalMux I__12877 (
            .O(N__55209),
            .I(N__55206));
    Span4Mux_s3_h I__12876 (
            .O(N__55206),
            .I(N__55202));
    CEMux I__12875 (
            .O(N__55205),
            .I(N__55199));
    Span4Mux_h I__12874 (
            .O(N__55202),
            .I(N__55194));
    LocalMux I__12873 (
            .O(N__55199),
            .I(N__55194));
    Span4Mux_v I__12872 (
            .O(N__55194),
            .I(N__55191));
    Span4Mux_h I__12871 (
            .O(N__55191),
            .I(N__55188));
    Span4Mux_h I__12870 (
            .O(N__55188),
            .I(N__55185));
    Span4Mux_h I__12869 (
            .O(N__55185),
            .I(N__55182));
    Odrv4 I__12868 (
            .O(N__55182),
            .I(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ));
    InMux I__12867 (
            .O(N__55179),
            .I(N__55176));
    LocalMux I__12866 (
            .O(N__55176),
            .I(N__55173));
    Odrv4 I__12865 (
            .O(N__55173),
            .I(\pid_side.O_1_18 ));
    InMux I__12864 (
            .O(N__55170),
            .I(N__55165));
    InMux I__12863 (
            .O(N__55169),
            .I(N__55162));
    InMux I__12862 (
            .O(N__55168),
            .I(N__55159));
    LocalMux I__12861 (
            .O(N__55165),
            .I(N__55154));
    LocalMux I__12860 (
            .O(N__55162),
            .I(N__55154));
    LocalMux I__12859 (
            .O(N__55159),
            .I(N__55151));
    Span4Mux_h I__12858 (
            .O(N__55154),
            .I(N__55148));
    Span4Mux_h I__12857 (
            .O(N__55151),
            .I(N__55145));
    Odrv4 I__12856 (
            .O(N__55148),
            .I(\pid_side.error_d_regZ0Z_14 ));
    Odrv4 I__12855 (
            .O(N__55145),
            .I(\pid_side.error_d_regZ0Z_14 ));
    InMux I__12854 (
            .O(N__55140),
            .I(N__55137));
    LocalMux I__12853 (
            .O(N__55137),
            .I(\pid_side.O_1_7 ));
    InMux I__12852 (
            .O(N__55134),
            .I(N__55125));
    InMux I__12851 (
            .O(N__55133),
            .I(N__55125));
    InMux I__12850 (
            .O(N__55132),
            .I(N__55125));
    LocalMux I__12849 (
            .O(N__55125),
            .I(N__55122));
    Span4Mux_v I__12848 (
            .O(N__55122),
            .I(N__55119));
    Odrv4 I__12847 (
            .O(N__55119),
            .I(\pid_side.error_d_regZ0Z_3 ));
    InMux I__12846 (
            .O(N__55116),
            .I(N__55113));
    LocalMux I__12845 (
            .O(N__55113),
            .I(N__55110));
    Span4Mux_h I__12844 (
            .O(N__55110),
            .I(N__55107));
    Odrv4 I__12843 (
            .O(N__55107),
            .I(\pid_side.O_1_17 ));
    InMux I__12842 (
            .O(N__55104),
            .I(N__55095));
    InMux I__12841 (
            .O(N__55103),
            .I(N__55095));
    InMux I__12840 (
            .O(N__55102),
            .I(N__55095));
    LocalMux I__12839 (
            .O(N__55095),
            .I(N__55092));
    Span12Mux_v I__12838 (
            .O(N__55092),
            .I(N__55089));
    Odrv12 I__12837 (
            .O(N__55089),
            .I(\pid_side.error_d_regZ0Z_13 ));
    InMux I__12836 (
            .O(N__55086),
            .I(N__55083));
    LocalMux I__12835 (
            .O(N__55083),
            .I(\pid_side.O_1_14 ));
    InMux I__12834 (
            .O(N__55080),
            .I(N__55075));
    InMux I__12833 (
            .O(N__55079),
            .I(N__55070));
    InMux I__12832 (
            .O(N__55078),
            .I(N__55070));
    LocalMux I__12831 (
            .O(N__55075),
            .I(N__55067));
    LocalMux I__12830 (
            .O(N__55070),
            .I(N__55064));
    Span4Mux_v I__12829 (
            .O(N__55067),
            .I(N__55061));
    Span4Mux_h I__12828 (
            .O(N__55064),
            .I(N__55058));
    Odrv4 I__12827 (
            .O(N__55061),
            .I(\pid_side.error_d_regZ0Z_10 ));
    Odrv4 I__12826 (
            .O(N__55058),
            .I(\pid_side.error_d_regZ0Z_10 ));
    InMux I__12825 (
            .O(N__55053),
            .I(N__55050));
    LocalMux I__12824 (
            .O(N__55050),
            .I(N__55047));
    Odrv4 I__12823 (
            .O(N__55047),
            .I(\pid_side.O_1_23 ));
    InMux I__12822 (
            .O(N__55044),
            .I(N__55035));
    InMux I__12821 (
            .O(N__55043),
            .I(N__55035));
    InMux I__12820 (
            .O(N__55042),
            .I(N__55035));
    LocalMux I__12819 (
            .O(N__55035),
            .I(N__55032));
    Odrv12 I__12818 (
            .O(N__55032),
            .I(\pid_side.error_d_regZ0Z_19 ));
    InMux I__12817 (
            .O(N__55029),
            .I(N__55026));
    LocalMux I__12816 (
            .O(N__55026),
            .I(N__55023));
    Odrv4 I__12815 (
            .O(N__55023),
            .I(\pid_side.O_1_24 ));
    InMux I__12814 (
            .O(N__55020),
            .I(N__55017));
    LocalMux I__12813 (
            .O(N__55017),
            .I(\pid_side.O_1_10 ));
    InMux I__12812 (
            .O(N__55014),
            .I(N__55011));
    LocalMux I__12811 (
            .O(N__55011),
            .I(N__55006));
    InMux I__12810 (
            .O(N__55010),
            .I(N__55001));
    InMux I__12809 (
            .O(N__55009),
            .I(N__55001));
    Span4Mux_h I__12808 (
            .O(N__55006),
            .I(N__54996));
    LocalMux I__12807 (
            .O(N__55001),
            .I(N__54996));
    Odrv4 I__12806 (
            .O(N__54996),
            .I(\pid_side.error_d_regZ0Z_6 ));
    InMux I__12805 (
            .O(N__54993),
            .I(N__54990));
    LocalMux I__12804 (
            .O(N__54990),
            .I(N__54987));
    Odrv4 I__12803 (
            .O(N__54987),
            .I(\pid_side.O_1_22 ));
    InMux I__12802 (
            .O(N__54984),
            .I(N__54975));
    InMux I__12801 (
            .O(N__54983),
            .I(N__54975));
    InMux I__12800 (
            .O(N__54982),
            .I(N__54975));
    LocalMux I__12799 (
            .O(N__54975),
            .I(N__54972));
    Span4Mux_h I__12798 (
            .O(N__54972),
            .I(N__54969));
    Odrv4 I__12797 (
            .O(N__54969),
            .I(\pid_side.error_d_regZ0Z_18 ));
    InMux I__12796 (
            .O(N__54966),
            .I(N__54963));
    LocalMux I__12795 (
            .O(N__54963),
            .I(\pid_side.O_1_11 ));
    InMux I__12794 (
            .O(N__54960),
            .I(N__54954));
    InMux I__12793 (
            .O(N__54959),
            .I(N__54947));
    InMux I__12792 (
            .O(N__54958),
            .I(N__54947));
    InMux I__12791 (
            .O(N__54957),
            .I(N__54947));
    LocalMux I__12790 (
            .O(N__54954),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    LocalMux I__12789 (
            .O(N__54947),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    InMux I__12788 (
            .O(N__54942),
            .I(N__54939));
    LocalMux I__12787 (
            .O(N__54939),
            .I(N__54936));
    Span4Mux_h I__12786 (
            .O(N__54936),
            .I(N__54933));
    Odrv4 I__12785 (
            .O(N__54933),
            .I(\pid_side.error_p_reg_esr_RNIBNBR2Z0Z_7 ));
    InMux I__12784 (
            .O(N__54930),
            .I(N__54924));
    InMux I__12783 (
            .O(N__54929),
            .I(N__54917));
    InMux I__12782 (
            .O(N__54928),
            .I(N__54917));
    InMux I__12781 (
            .O(N__54927),
            .I(N__54917));
    LocalMux I__12780 (
            .O(N__54924),
            .I(\pid_side.error_p_regZ0Z_6 ));
    LocalMux I__12779 (
            .O(N__54917),
            .I(\pid_side.error_p_regZ0Z_6 ));
    InMux I__12778 (
            .O(N__54912),
            .I(N__54906));
    InMux I__12777 (
            .O(N__54911),
            .I(N__54899));
    InMux I__12776 (
            .O(N__54910),
            .I(N__54899));
    InMux I__12775 (
            .O(N__54909),
            .I(N__54899));
    LocalMux I__12774 (
            .O(N__54906),
            .I(\pid_side.error_d_reg_prevZ0Z_6 ));
    LocalMux I__12773 (
            .O(N__54899),
            .I(\pid_side.error_d_reg_prevZ0Z_6 ));
    InMux I__12772 (
            .O(N__54894),
            .I(N__54891));
    LocalMux I__12771 (
            .O(N__54891),
            .I(N__54888));
    Span12Mux_h I__12770 (
            .O(N__54888),
            .I(N__54885));
    Odrv12 I__12769 (
            .O(N__54885),
            .I(\pid_side.un1_pid_prereg_50_0 ));
    InMux I__12768 (
            .O(N__54882),
            .I(N__54879));
    LocalMux I__12767 (
            .O(N__54879),
            .I(N__54876));
    Span4Mux_h I__12766 (
            .O(N__54876),
            .I(N__54873));
    Odrv4 I__12765 (
            .O(N__54873),
            .I(\pid_side.O_1_15 ));
    InMux I__12764 (
            .O(N__54870),
            .I(N__54865));
    InMux I__12763 (
            .O(N__54869),
            .I(N__54860));
    InMux I__12762 (
            .O(N__54868),
            .I(N__54860));
    LocalMux I__12761 (
            .O(N__54865),
            .I(N__54857));
    LocalMux I__12760 (
            .O(N__54860),
            .I(N__54854));
    Span4Mux_h I__12759 (
            .O(N__54857),
            .I(N__54851));
    Odrv4 I__12758 (
            .O(N__54854),
            .I(\pid_side.error_d_regZ0Z_11 ));
    Odrv4 I__12757 (
            .O(N__54851),
            .I(\pid_side.error_d_regZ0Z_11 ));
    InMux I__12756 (
            .O(N__54846),
            .I(N__54843));
    LocalMux I__12755 (
            .O(N__54843),
            .I(N__54840));
    Odrv4 I__12754 (
            .O(N__54840),
            .I(\pid_side.O_1_21 ));
    InMux I__12753 (
            .O(N__54837),
            .I(N__54832));
    InMux I__12752 (
            .O(N__54836),
            .I(N__54827));
    InMux I__12751 (
            .O(N__54835),
            .I(N__54827));
    LocalMux I__12750 (
            .O(N__54832),
            .I(\pid_side.error_d_regZ0Z_17 ));
    LocalMux I__12749 (
            .O(N__54827),
            .I(\pid_side.error_d_regZ0Z_17 ));
    InMux I__12748 (
            .O(N__54822),
            .I(N__54819));
    LocalMux I__12747 (
            .O(N__54819),
            .I(N__54816));
    Odrv4 I__12746 (
            .O(N__54816),
            .I(\pid_side.O_1_19 ));
    InMux I__12745 (
            .O(N__54813),
            .I(N__54809));
    InMux I__12744 (
            .O(N__54812),
            .I(N__54805));
    LocalMux I__12743 (
            .O(N__54809),
            .I(N__54802));
    InMux I__12742 (
            .O(N__54808),
            .I(N__54799));
    LocalMux I__12741 (
            .O(N__54805),
            .I(N__54792));
    Span4Mux_h I__12740 (
            .O(N__54802),
            .I(N__54792));
    LocalMux I__12739 (
            .O(N__54799),
            .I(N__54792));
    Span4Mux_h I__12738 (
            .O(N__54792),
            .I(N__54789));
    Odrv4 I__12737 (
            .O(N__54789),
            .I(\pid_side.error_d_regZ0Z_15 ));
    InMux I__12736 (
            .O(N__54786),
            .I(N__54783));
    LocalMux I__12735 (
            .O(N__54783),
            .I(N__54780));
    Odrv4 I__12734 (
            .O(N__54780),
            .I(\pid_side.O_1_12 ));
    InMux I__12733 (
            .O(N__54777),
            .I(N__54768));
    InMux I__12732 (
            .O(N__54776),
            .I(N__54768));
    InMux I__12731 (
            .O(N__54775),
            .I(N__54768));
    LocalMux I__12730 (
            .O(N__54768),
            .I(N__54765));
    Odrv4 I__12729 (
            .O(N__54765),
            .I(\pid_side.error_d_regZ0Z_8 ));
    InMux I__12728 (
            .O(N__54762),
            .I(N__54759));
    LocalMux I__12727 (
            .O(N__54759),
            .I(N__54756));
    Odrv4 I__12726 (
            .O(N__54756),
            .I(\pid_side.O_1_9 ));
    InMux I__12725 (
            .O(N__54753),
            .I(N__54748));
    InMux I__12724 (
            .O(N__54752),
            .I(N__54743));
    InMux I__12723 (
            .O(N__54751),
            .I(N__54743));
    LocalMux I__12722 (
            .O(N__54748),
            .I(N__54740));
    LocalMux I__12721 (
            .O(N__54743),
            .I(N__54737));
    Span4Mux_h I__12720 (
            .O(N__54740),
            .I(N__54734));
    Span4Mux_h I__12719 (
            .O(N__54737),
            .I(N__54731));
    Span4Mux_v I__12718 (
            .O(N__54734),
            .I(N__54728));
    Span4Mux_v I__12717 (
            .O(N__54731),
            .I(N__54725));
    Odrv4 I__12716 (
            .O(N__54728),
            .I(\pid_side.error_d_regZ0Z_5 ));
    Odrv4 I__12715 (
            .O(N__54725),
            .I(\pid_side.error_d_regZ0Z_5 ));
    InMux I__12714 (
            .O(N__54720),
            .I(N__54717));
    LocalMux I__12713 (
            .O(N__54717),
            .I(N__54714));
    Odrv4 I__12712 (
            .O(N__54714),
            .I(\pid_side.O_1_16 ));
    InMux I__12711 (
            .O(N__54711),
            .I(N__54702));
    InMux I__12710 (
            .O(N__54710),
            .I(N__54702));
    InMux I__12709 (
            .O(N__54709),
            .I(N__54702));
    LocalMux I__12708 (
            .O(N__54702),
            .I(N__54699));
    Span4Mux_h I__12707 (
            .O(N__54699),
            .I(N__54696));
    Odrv4 I__12706 (
            .O(N__54696),
            .I(\pid_side.error_d_regZ0Z_12 ));
    InMux I__12705 (
            .O(N__54693),
            .I(N__54690));
    LocalMux I__12704 (
            .O(N__54690),
            .I(\pid_side.O_2_11 ));
    InMux I__12703 (
            .O(N__54687),
            .I(N__54684));
    LocalMux I__12702 (
            .O(N__54684),
            .I(\pid_side.O_2_23 ));
    InMux I__12701 (
            .O(N__54681),
            .I(N__54675));
    InMux I__12700 (
            .O(N__54680),
            .I(N__54675));
    LocalMux I__12699 (
            .O(N__54675),
            .I(N__54672));
    Span4Mux_h I__12698 (
            .O(N__54672),
            .I(N__54669));
    Span4Mux_v I__12697 (
            .O(N__54669),
            .I(N__54666));
    Odrv4 I__12696 (
            .O(N__54666),
            .I(\pid_side.error_p_regZ0Z_19 ));
    InMux I__12695 (
            .O(N__54663),
            .I(N__54660));
    LocalMux I__12694 (
            .O(N__54660),
            .I(\pid_side.O_2_16 ));
    CascadeMux I__12693 (
            .O(N__54657),
            .I(N__54653));
    CascadeMux I__12692 (
            .O(N__54656),
            .I(N__54650));
    InMux I__12691 (
            .O(N__54653),
            .I(N__54642));
    InMux I__12690 (
            .O(N__54650),
            .I(N__54642));
    InMux I__12689 (
            .O(N__54649),
            .I(N__54642));
    LocalMux I__12688 (
            .O(N__54642),
            .I(N__54639));
    Span4Mux_h I__12687 (
            .O(N__54639),
            .I(N__54636));
    Odrv4 I__12686 (
            .O(N__54636),
            .I(\pid_side.error_p_regZ0Z_12 ));
    InMux I__12685 (
            .O(N__54633),
            .I(N__54630));
    LocalMux I__12684 (
            .O(N__54630),
            .I(N__54626));
    InMux I__12683 (
            .O(N__54629),
            .I(N__54623));
    Span4Mux_v I__12682 (
            .O(N__54626),
            .I(N__54620));
    LocalMux I__12681 (
            .O(N__54623),
            .I(\pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6 ));
    Odrv4 I__12680 (
            .O(N__54620),
            .I(\pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6 ));
    CascadeMux I__12679 (
            .O(N__54615),
            .I(\pid_side.un1_pid_prereg_60_0_cascade_ ));
    CascadeMux I__12678 (
            .O(N__54612),
            .I(N__54609));
    InMux I__12677 (
            .O(N__54609),
            .I(N__54606));
    LocalMux I__12676 (
            .O(N__54606),
            .I(N__54603));
    Span4Mux_h I__12675 (
            .O(N__54603),
            .I(N__54600));
    Span4Mux_s1_h I__12674 (
            .O(N__54600),
            .I(N__54597));
    Odrv4 I__12673 (
            .O(N__54597),
            .I(\pid_side.error_p_reg_esr_RNI1DBR2Z0Z_6 ));
    CascadeMux I__12672 (
            .O(N__54594),
            .I(\pid_side.N_1570_i_cascade_ ));
    CascadeMux I__12671 (
            .O(N__54591),
            .I(N__54588));
    InMux I__12670 (
            .O(N__54588),
            .I(N__54585));
    LocalMux I__12669 (
            .O(N__54585),
            .I(N__54582));
    Span4Mux_h I__12668 (
            .O(N__54582),
            .I(N__54579));
    Odrv4 I__12667 (
            .O(N__54579),
            .I(\pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7 ));
    InMux I__12666 (
            .O(N__54576),
            .I(N__54573));
    LocalMux I__12665 (
            .O(N__54573),
            .I(\pid_side.un1_pid_prereg_70_0 ));
    InMux I__12664 (
            .O(N__54570),
            .I(N__54564));
    InMux I__12663 (
            .O(N__54569),
            .I(N__54557));
    InMux I__12662 (
            .O(N__54568),
            .I(N__54557));
    InMux I__12661 (
            .O(N__54567),
            .I(N__54557));
    LocalMux I__12660 (
            .O(N__54564),
            .I(\pid_side.error_p_regZ0Z_7 ));
    LocalMux I__12659 (
            .O(N__54557),
            .I(\pid_side.error_p_regZ0Z_7 ));
    CascadeMux I__12658 (
            .O(N__54552),
            .I(\pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7_cascade_ ));
    InMux I__12657 (
            .O(N__54549),
            .I(N__54546));
    LocalMux I__12656 (
            .O(N__54546),
            .I(N__54543));
    Span4Mux_v I__12655 (
            .O(N__54543),
            .I(N__54540));
    Odrv4 I__12654 (
            .O(N__54540),
            .I(\pid_side.O_1_6 ));
    InMux I__12653 (
            .O(N__54537),
            .I(N__54532));
    InMux I__12652 (
            .O(N__54536),
            .I(N__54527));
    InMux I__12651 (
            .O(N__54535),
            .I(N__54527));
    LocalMux I__12650 (
            .O(N__54532),
            .I(\pid_side.error_d_regZ0Z_2 ));
    LocalMux I__12649 (
            .O(N__54527),
            .I(\pid_side.error_d_regZ0Z_2 ));
    InMux I__12648 (
            .O(N__54522),
            .I(N__54519));
    LocalMux I__12647 (
            .O(N__54519),
            .I(N__54516));
    Odrv4 I__12646 (
            .O(N__54516),
            .I(\pid_side.O_2_17 ));
    InMux I__12645 (
            .O(N__54513),
            .I(N__54507));
    InMux I__12644 (
            .O(N__54512),
            .I(N__54507));
    LocalMux I__12643 (
            .O(N__54507),
            .I(N__54504));
    Odrv4 I__12642 (
            .O(N__54504),
            .I(\pid_side.error_p_regZ0Z_13 ));
    InMux I__12641 (
            .O(N__54501),
            .I(N__54498));
    LocalMux I__12640 (
            .O(N__54498),
            .I(\pid_side.O_2_12 ));
    CascadeMux I__12639 (
            .O(N__54495),
            .I(N__54490));
    InMux I__12638 (
            .O(N__54494),
            .I(N__54482));
    InMux I__12637 (
            .O(N__54493),
            .I(N__54482));
    InMux I__12636 (
            .O(N__54490),
            .I(N__54482));
    InMux I__12635 (
            .O(N__54489),
            .I(N__54479));
    LocalMux I__12634 (
            .O(N__54482),
            .I(N__54476));
    LocalMux I__12633 (
            .O(N__54479),
            .I(\pid_side.error_p_regZ0Z_8 ));
    Odrv4 I__12632 (
            .O(N__54476),
            .I(\pid_side.error_p_regZ0Z_8 ));
    InMux I__12631 (
            .O(N__54471),
            .I(N__54468));
    LocalMux I__12630 (
            .O(N__54468),
            .I(N__54465));
    Odrv4 I__12629 (
            .O(N__54465),
            .I(\pid_side.O_2_24 ));
    InMux I__12628 (
            .O(N__54462),
            .I(N__54459));
    LocalMux I__12627 (
            .O(N__54459),
            .I(N__54455));
    InMux I__12626 (
            .O(N__54458),
            .I(N__54452));
    Span4Mux_v I__12625 (
            .O(N__54455),
            .I(N__54447));
    LocalMux I__12624 (
            .O(N__54452),
            .I(N__54447));
    Sp12to4 I__12623 (
            .O(N__54447),
            .I(N__54444));
    Odrv12 I__12622 (
            .O(N__54444),
            .I(\pid_side.error_p_regZ0Z_20 ));
    InMux I__12621 (
            .O(N__54441),
            .I(N__54438));
    LocalMux I__12620 (
            .O(N__54438),
            .I(N__54435));
    Odrv4 I__12619 (
            .O(N__54435),
            .I(\pid_side.O_2_18 ));
    InMux I__12618 (
            .O(N__54432),
            .I(N__54428));
    InMux I__12617 (
            .O(N__54431),
            .I(N__54425));
    LocalMux I__12616 (
            .O(N__54428),
            .I(N__54422));
    LocalMux I__12615 (
            .O(N__54425),
            .I(N__54419));
    Span4Mux_h I__12614 (
            .O(N__54422),
            .I(N__54416));
    Odrv12 I__12613 (
            .O(N__54419),
            .I(\pid_side.error_p_regZ0Z_14 ));
    Odrv4 I__12612 (
            .O(N__54416),
            .I(\pid_side.error_p_regZ0Z_14 ));
    InMux I__12611 (
            .O(N__54411),
            .I(N__54408));
    LocalMux I__12610 (
            .O(N__54408),
            .I(\pid_side.O_2_14 ));
    InMux I__12609 (
            .O(N__54405),
            .I(N__54402));
    LocalMux I__12608 (
            .O(N__54402),
            .I(N__54398));
    InMux I__12607 (
            .O(N__54401),
            .I(N__54395));
    Span4Mux_h I__12606 (
            .O(N__54398),
            .I(N__54392));
    LocalMux I__12605 (
            .O(N__54395),
            .I(N__54389));
    Odrv4 I__12604 (
            .O(N__54392),
            .I(\pid_side.error_p_regZ0Z_10 ));
    Odrv12 I__12603 (
            .O(N__54389),
            .I(\pid_side.error_p_regZ0Z_10 ));
    InMux I__12602 (
            .O(N__54384),
            .I(N__54381));
    LocalMux I__12601 (
            .O(N__54381),
            .I(\pid_side.O_2_19 ));
    InMux I__12600 (
            .O(N__54378),
            .I(N__54374));
    InMux I__12599 (
            .O(N__54377),
            .I(N__54371));
    LocalMux I__12598 (
            .O(N__54374),
            .I(N__54366));
    LocalMux I__12597 (
            .O(N__54371),
            .I(N__54366));
    Span4Mux_h I__12596 (
            .O(N__54366),
            .I(N__54363));
    Odrv4 I__12595 (
            .O(N__54363),
            .I(\pid_side.error_p_regZ0Z_15 ));
    InMux I__12594 (
            .O(N__54360),
            .I(N__54357));
    LocalMux I__12593 (
            .O(N__54357),
            .I(\pid_side.O_2_10 ));
    InMux I__12592 (
            .O(N__54354),
            .I(N__54351));
    LocalMux I__12591 (
            .O(N__54351),
            .I(\pid_side.O_2_13 ));
    InMux I__12590 (
            .O(N__54348),
            .I(N__54343));
    InMux I__12589 (
            .O(N__54347),
            .I(N__54340));
    InMux I__12588 (
            .O(N__54346),
            .I(N__54337));
    LocalMux I__12587 (
            .O(N__54343),
            .I(N__54334));
    LocalMux I__12586 (
            .O(N__54340),
            .I(\pid_side.error_p_regZ0Z_9 ));
    LocalMux I__12585 (
            .O(N__54337),
            .I(\pid_side.error_p_regZ0Z_9 ));
    Odrv4 I__12584 (
            .O(N__54334),
            .I(\pid_side.error_p_regZ0Z_9 ));
    InMux I__12583 (
            .O(N__54327),
            .I(N__54324));
    LocalMux I__12582 (
            .O(N__54324),
            .I(N__54321));
    Span4Mux_h I__12581 (
            .O(N__54321),
            .I(N__54318));
    Odrv4 I__12580 (
            .O(N__54318),
            .I(\pid_front.O_14 ));
    InMux I__12579 (
            .O(N__54315),
            .I(N__54309));
    InMux I__12578 (
            .O(N__54314),
            .I(N__54309));
    LocalMux I__12577 (
            .O(N__54309),
            .I(N__54305));
    InMux I__12576 (
            .O(N__54308),
            .I(N__54302));
    Span4Mux_h I__12575 (
            .O(N__54305),
            .I(N__54297));
    LocalMux I__12574 (
            .O(N__54302),
            .I(N__54297));
    Sp12to4 I__12573 (
            .O(N__54297),
            .I(N__54294));
    Span12Mux_s7_v I__12572 (
            .O(N__54294),
            .I(N__54291));
    Odrv12 I__12571 (
            .O(N__54291),
            .I(\pid_front.error_d_regZ0Z_10 ));
    InMux I__12570 (
            .O(N__54288),
            .I(N__54285));
    LocalMux I__12569 (
            .O(N__54285),
            .I(N__54282));
    Odrv4 I__12568 (
            .O(N__54282),
            .I(\pid_side.O_2_8 ));
    InMux I__12567 (
            .O(N__54279),
            .I(N__54273));
    InMux I__12566 (
            .O(N__54278),
            .I(N__54273));
    LocalMux I__12565 (
            .O(N__54273),
            .I(N__54270));
    Odrv4 I__12564 (
            .O(N__54270),
            .I(\pid_side.error_p_regZ0Z_4 ));
    InMux I__12563 (
            .O(N__54267),
            .I(N__54264));
    LocalMux I__12562 (
            .O(N__54264),
            .I(\pid_side.O_2_5 ));
    CascadeMux I__12561 (
            .O(N__54261),
            .I(N__54258));
    InMux I__12560 (
            .O(N__54258),
            .I(N__54252));
    InMux I__12559 (
            .O(N__54257),
            .I(N__54252));
    LocalMux I__12558 (
            .O(N__54252),
            .I(N__54249));
    Odrv4 I__12557 (
            .O(N__54249),
            .I(\pid_side.error_p_regZ0Z_1 ));
    InMux I__12556 (
            .O(N__54246),
            .I(N__54243));
    LocalMux I__12555 (
            .O(N__54243),
            .I(\pid_side.O_2_7 ));
    InMux I__12554 (
            .O(N__54240),
            .I(N__54234));
    InMux I__12553 (
            .O(N__54239),
            .I(N__54234));
    LocalMux I__12552 (
            .O(N__54234),
            .I(\pid_side.error_p_regZ0Z_3 ));
    InMux I__12551 (
            .O(N__54231),
            .I(N__54228));
    LocalMux I__12550 (
            .O(N__54228),
            .I(N__54225));
    Span4Mux_h I__12549 (
            .O(N__54225),
            .I(N__54222));
    Odrv4 I__12548 (
            .O(N__54222),
            .I(\pid_side.O_2_22 ));
    InMux I__12547 (
            .O(N__54219),
            .I(N__54213));
    InMux I__12546 (
            .O(N__54218),
            .I(N__54213));
    LocalMux I__12545 (
            .O(N__54213),
            .I(N__54210));
    Span4Mux_v I__12544 (
            .O(N__54210),
            .I(N__54207));
    Odrv4 I__12543 (
            .O(N__54207),
            .I(\pid_side.error_p_regZ0Z_18 ));
    InMux I__12542 (
            .O(N__54204),
            .I(N__54201));
    LocalMux I__12541 (
            .O(N__54201),
            .I(\pid_side.O_2_6 ));
    InMux I__12540 (
            .O(N__54198),
            .I(N__54192));
    InMux I__12539 (
            .O(N__54197),
            .I(N__54192));
    LocalMux I__12538 (
            .O(N__54192),
            .I(\pid_side.error_p_regZ0Z_2 ));
    InMux I__12537 (
            .O(N__54189),
            .I(N__54186));
    LocalMux I__12536 (
            .O(N__54186),
            .I(N__54183));
    Odrv4 I__12535 (
            .O(N__54183),
            .I(\pid_side.O_2_20 ));
    InMux I__12534 (
            .O(N__54180),
            .I(N__54174));
    InMux I__12533 (
            .O(N__54179),
            .I(N__54174));
    LocalMux I__12532 (
            .O(N__54174),
            .I(N__54171));
    Span4Mux_v I__12531 (
            .O(N__54171),
            .I(N__54168));
    Span4Mux_h I__12530 (
            .O(N__54168),
            .I(N__54165));
    Odrv4 I__12529 (
            .O(N__54165),
            .I(\pid_side.error_p_regZ0Z_16 ));
    InMux I__12528 (
            .O(N__54162),
            .I(N__54159));
    LocalMux I__12527 (
            .O(N__54159),
            .I(N__54156));
    Odrv4 I__12526 (
            .O(N__54156),
            .I(\pid_side.O_2_21 ));
    InMux I__12525 (
            .O(N__54153),
            .I(N__54147));
    InMux I__12524 (
            .O(N__54152),
            .I(N__54147));
    LocalMux I__12523 (
            .O(N__54147),
            .I(N__54144));
    Odrv4 I__12522 (
            .O(N__54144),
            .I(\pid_side.error_p_regZ0Z_17 ));
    InMux I__12521 (
            .O(N__54141),
            .I(N__54136));
    InMux I__12520 (
            .O(N__54140),
            .I(N__54133));
    InMux I__12519 (
            .O(N__54139),
            .I(N__54130));
    LocalMux I__12518 (
            .O(N__54136),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    LocalMux I__12517 (
            .O(N__54133),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    LocalMux I__12516 (
            .O(N__54130),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    CascadeMux I__12515 (
            .O(N__54123),
            .I(N__54118));
    InMux I__12514 (
            .O(N__54122),
            .I(N__54113));
    InMux I__12513 (
            .O(N__54121),
            .I(N__54113));
    InMux I__12512 (
            .O(N__54118),
            .I(N__54110));
    LocalMux I__12511 (
            .O(N__54113),
            .I(N__54107));
    LocalMux I__12510 (
            .O(N__54110),
            .I(\pid_side.un1_pid_prereg_41 ));
    Odrv4 I__12509 (
            .O(N__54107),
            .I(\pid_side.un1_pid_prereg_41 ));
    InMux I__12508 (
            .O(N__54102),
            .I(N__54099));
    LocalMux I__12507 (
            .O(N__54099),
            .I(N__54096));
    Span4Mux_v I__12506 (
            .O(N__54096),
            .I(N__54091));
    InMux I__12505 (
            .O(N__54095),
            .I(N__54086));
    InMux I__12504 (
            .O(N__54094),
            .I(N__54086));
    Odrv4 I__12503 (
            .O(N__54091),
            .I(\pid_side.un1_pid_prereg_42 ));
    LocalMux I__12502 (
            .O(N__54086),
            .I(\pid_side.un1_pid_prereg_42 ));
    CascadeMux I__12501 (
            .O(N__54081),
            .I(N__54078));
    InMux I__12500 (
            .O(N__54078),
            .I(N__54072));
    InMux I__12499 (
            .O(N__54077),
            .I(N__54072));
    LocalMux I__12498 (
            .O(N__54072),
            .I(\pid_side.error_d_reg_prevZ0Z_17 ));
    InMux I__12497 (
            .O(N__54069),
            .I(N__54066));
    LocalMux I__12496 (
            .O(N__54066),
            .I(N__54063));
    Span4Mux_h I__12495 (
            .O(N__54063),
            .I(N__54060));
    Odrv4 I__12494 (
            .O(N__54060),
            .I(\pid_side.O_1_13 ));
    InMux I__12493 (
            .O(N__54057),
            .I(N__54054));
    LocalMux I__12492 (
            .O(N__54054),
            .I(N__54049));
    InMux I__12491 (
            .O(N__54053),
            .I(N__54044));
    InMux I__12490 (
            .O(N__54052),
            .I(N__54044));
    Sp12to4 I__12489 (
            .O(N__54049),
            .I(N__54039));
    LocalMux I__12488 (
            .O(N__54044),
            .I(N__54039));
    Odrv12 I__12487 (
            .O(N__54039),
            .I(\pid_side.error_d_regZ0Z_9 ));
    CascadeMux I__12486 (
            .O(N__54036),
            .I(N__54031));
    CascadeMux I__12485 (
            .O(N__54035),
            .I(N__54025));
    InMux I__12484 (
            .O(N__54034),
            .I(N__54022));
    InMux I__12483 (
            .O(N__54031),
            .I(N__54015));
    InMux I__12482 (
            .O(N__54030),
            .I(N__54015));
    InMux I__12481 (
            .O(N__54029),
            .I(N__54015));
    InMux I__12480 (
            .O(N__54028),
            .I(N__54010));
    InMux I__12479 (
            .O(N__54025),
            .I(N__54010));
    LocalMux I__12478 (
            .O(N__54022),
            .I(N__54007));
    LocalMux I__12477 (
            .O(N__54015),
            .I(N__54002));
    LocalMux I__12476 (
            .O(N__54010),
            .I(N__54002));
    Span4Mux_h I__12475 (
            .O(N__54007),
            .I(N__53999));
    Span4Mux_h I__12474 (
            .O(N__54002),
            .I(N__53996));
    Odrv4 I__12473 (
            .O(N__53999),
            .I(\pid_side.un1_pid_prereg_93 ));
    Odrv4 I__12472 (
            .O(N__53996),
            .I(\pid_side.un1_pid_prereg_93 ));
    CascadeMux I__12471 (
            .O(N__53991),
            .I(N__53987));
    InMux I__12470 (
            .O(N__53990),
            .I(N__53984));
    InMux I__12469 (
            .O(N__53987),
            .I(N__53975));
    LocalMux I__12468 (
            .O(N__53984),
            .I(N__53971));
    InMux I__12467 (
            .O(N__53983),
            .I(N__53962));
    InMux I__12466 (
            .O(N__53982),
            .I(N__53962));
    InMux I__12465 (
            .O(N__53981),
            .I(N__53962));
    InMux I__12464 (
            .O(N__53980),
            .I(N__53962));
    InMux I__12463 (
            .O(N__53979),
            .I(N__53957));
    InMux I__12462 (
            .O(N__53978),
            .I(N__53957));
    LocalMux I__12461 (
            .O(N__53975),
            .I(N__53954));
    InMux I__12460 (
            .O(N__53974),
            .I(N__53951));
    Span4Mux_h I__12459 (
            .O(N__53971),
            .I(N__53948));
    LocalMux I__12458 (
            .O(N__53962),
            .I(N__53939));
    LocalMux I__12457 (
            .O(N__53957),
            .I(N__53939));
    Span4Mux_v I__12456 (
            .O(N__53954),
            .I(N__53939));
    LocalMux I__12455 (
            .O(N__53951),
            .I(N__53939));
    Span4Mux_v I__12454 (
            .O(N__53948),
            .I(N__53936));
    Span4Mux_v I__12453 (
            .O(N__53939),
            .I(N__53933));
    Odrv4 I__12452 (
            .O(N__53936),
            .I(\pid_side.un1_pid_prereg_92 ));
    Odrv4 I__12451 (
            .O(N__53933),
            .I(\pid_side.un1_pid_prereg_92 ));
    InMux I__12450 (
            .O(N__53928),
            .I(N__53925));
    LocalMux I__12449 (
            .O(N__53925),
            .I(N__53922));
    Span4Mux_h I__12448 (
            .O(N__53922),
            .I(N__53919));
    Odrv4 I__12447 (
            .O(N__53919),
            .I(\pid_front.O_12 ));
    CascadeMux I__12446 (
            .O(N__53916),
            .I(N__53912));
    InMux I__12445 (
            .O(N__53915),
            .I(N__53908));
    InMux I__12444 (
            .O(N__53912),
            .I(N__53905));
    InMux I__12443 (
            .O(N__53911),
            .I(N__53902));
    LocalMux I__12442 (
            .O(N__53908),
            .I(N__53899));
    LocalMux I__12441 (
            .O(N__53905),
            .I(N__53894));
    LocalMux I__12440 (
            .O(N__53902),
            .I(N__53894));
    Span4Mux_v I__12439 (
            .O(N__53899),
            .I(N__53891));
    Span4Mux_h I__12438 (
            .O(N__53894),
            .I(N__53888));
    Span4Mux_h I__12437 (
            .O(N__53891),
            .I(N__53885));
    Span4Mux_h I__12436 (
            .O(N__53888),
            .I(N__53882));
    Sp12to4 I__12435 (
            .O(N__53885),
            .I(N__53879));
    Span4Mux_h I__12434 (
            .O(N__53882),
            .I(N__53876));
    Span12Mux_h I__12433 (
            .O(N__53879),
            .I(N__53873));
    Span4Mux_h I__12432 (
            .O(N__53876),
            .I(N__53870));
    Odrv12 I__12431 (
            .O(N__53873),
            .I(\pid_front.error_d_regZ0Z_8 ));
    Odrv4 I__12430 (
            .O(N__53870),
            .I(\pid_front.error_d_regZ0Z_8 ));
    InMux I__12429 (
            .O(N__53865),
            .I(N__53862));
    LocalMux I__12428 (
            .O(N__53862),
            .I(N__53859));
    Span4Mux_h I__12427 (
            .O(N__53859),
            .I(N__53856));
    Odrv4 I__12426 (
            .O(N__53856),
            .I(\pid_front.O_16 ));
    InMux I__12425 (
            .O(N__53853),
            .I(N__53850));
    LocalMux I__12424 (
            .O(N__53850),
            .I(N__53845));
    InMux I__12423 (
            .O(N__53849),
            .I(N__53840));
    InMux I__12422 (
            .O(N__53848),
            .I(N__53840));
    Span4Mux_h I__12421 (
            .O(N__53845),
            .I(N__53835));
    LocalMux I__12420 (
            .O(N__53840),
            .I(N__53835));
    Sp12to4 I__12419 (
            .O(N__53835),
            .I(N__53832));
    Span12Mux_s7_v I__12418 (
            .O(N__53832),
            .I(N__53829));
    Span12Mux_h I__12417 (
            .O(N__53829),
            .I(N__53826));
    Odrv12 I__12416 (
            .O(N__53826),
            .I(\pid_front.error_d_regZ0Z_12 ));
    CascadeMux I__12415 (
            .O(N__53823),
            .I(N__53820));
    InMux I__12414 (
            .O(N__53820),
            .I(N__53816));
    InMux I__12413 (
            .O(N__53819),
            .I(N__53811));
    LocalMux I__12412 (
            .O(N__53816),
            .I(N__53808));
    InMux I__12411 (
            .O(N__53815),
            .I(N__53803));
    InMux I__12410 (
            .O(N__53814),
            .I(N__53803));
    LocalMux I__12409 (
            .O(N__53811),
            .I(\pid_side.error_p_regZ0Z_5 ));
    Odrv4 I__12408 (
            .O(N__53808),
            .I(\pid_side.error_p_regZ0Z_5 ));
    LocalMux I__12407 (
            .O(N__53803),
            .I(\pid_side.error_p_regZ0Z_5 ));
    InMux I__12406 (
            .O(N__53796),
            .I(N__53792));
    CascadeMux I__12405 (
            .O(N__53795),
            .I(N__53789));
    LocalMux I__12404 (
            .O(N__53792),
            .I(N__53785));
    InMux I__12403 (
            .O(N__53789),
            .I(N__53779));
    InMux I__12402 (
            .O(N__53788),
            .I(N__53779));
    Span4Mux_v I__12401 (
            .O(N__53785),
            .I(N__53776));
    InMux I__12400 (
            .O(N__53784),
            .I(N__53773));
    LocalMux I__12399 (
            .O(N__53779),
            .I(N__53770));
    Odrv4 I__12398 (
            .O(N__53776),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    LocalMux I__12397 (
            .O(N__53773),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    Odrv4 I__12396 (
            .O(N__53770),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    CascadeMux I__12395 (
            .O(N__53763),
            .I(\pid_side.N_1566_i_cascade_ ));
    CascadeMux I__12394 (
            .O(N__53760),
            .I(\pid_side.N_1578_i_cascade_ ));
    CascadeMux I__12393 (
            .O(N__53757),
            .I(N__53753));
    CascadeMux I__12392 (
            .O(N__53756),
            .I(N__53750));
    InMux I__12391 (
            .O(N__53753),
            .I(N__53747));
    InMux I__12390 (
            .O(N__53750),
            .I(N__53744));
    LocalMux I__12389 (
            .O(N__53747),
            .I(N__53741));
    LocalMux I__12388 (
            .O(N__53744),
            .I(N__53738));
    Span4Mux_h I__12387 (
            .O(N__53741),
            .I(N__53735));
    Odrv4 I__12386 (
            .O(N__53738),
            .I(\pid_side.error_d_reg_esr_RNID3MD1Z0Z_9 ));
    Odrv4 I__12385 (
            .O(N__53735),
            .I(\pid_side.error_d_reg_esr_RNID3MD1Z0Z_9 ));
    CascadeMux I__12384 (
            .O(N__53730),
            .I(\pid_side.N_1574_i_cascade_ ));
    CascadeMux I__12383 (
            .O(N__53727),
            .I(N__53724));
    InMux I__12382 (
            .O(N__53724),
            .I(N__53721));
    LocalMux I__12381 (
            .O(N__53721),
            .I(N__53718));
    Span4Mux_v I__12380 (
            .O(N__53718),
            .I(N__53715));
    Odrv4 I__12379 (
            .O(N__53715),
            .I(\pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8 ));
    InMux I__12378 (
            .O(N__53712),
            .I(N__53709));
    LocalMux I__12377 (
            .O(N__53709),
            .I(\pid_side.un1_pid_prereg_80_0 ));
    CascadeMux I__12376 (
            .O(N__53706),
            .I(\pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8_cascade_ ));
    InMux I__12375 (
            .O(N__53703),
            .I(N__53700));
    LocalMux I__12374 (
            .O(N__53700),
            .I(N__53697));
    Span4Mux_h I__12373 (
            .O(N__53697),
            .I(N__53694));
    Odrv4 I__12372 (
            .O(N__53694),
            .I(\pid_side.error_p_reg_esr_RNIL1CR2Z0Z_8 ));
    InMux I__12371 (
            .O(N__53691),
            .I(N__53685));
    InMux I__12370 (
            .O(N__53690),
            .I(N__53678));
    InMux I__12369 (
            .O(N__53689),
            .I(N__53678));
    InMux I__12368 (
            .O(N__53688),
            .I(N__53678));
    LocalMux I__12367 (
            .O(N__53685),
            .I(\pid_side.error_d_reg_prevZ0Z_8 ));
    LocalMux I__12366 (
            .O(N__53678),
            .I(\pid_side.error_d_reg_prevZ0Z_8 ));
    CascadeMux I__12365 (
            .O(N__53673),
            .I(N__53669));
    InMux I__12364 (
            .O(N__53672),
            .I(N__53666));
    InMux I__12363 (
            .O(N__53669),
            .I(N__53663));
    LocalMux I__12362 (
            .O(N__53666),
            .I(\pid_side.un1_pid_prereg_2 ));
    LocalMux I__12361 (
            .O(N__53663),
            .I(\pid_side.un1_pid_prereg_2 ));
    CascadeMux I__12360 (
            .O(N__53658),
            .I(\pid_side.un1_pid_prereg_2_cascade_ ));
    InMux I__12359 (
            .O(N__53655),
            .I(N__53652));
    LocalMux I__12358 (
            .O(N__53652),
            .I(N__53649));
    Odrv4 I__12357 (
            .O(N__53649),
            .I(\pid_side.error_p_reg_esr_RNIRPSK1Z0Z_2 ));
    InMux I__12356 (
            .O(N__53646),
            .I(N__53639));
    InMux I__12355 (
            .O(N__53645),
            .I(N__53639));
    InMux I__12354 (
            .O(N__53644),
            .I(N__53636));
    LocalMux I__12353 (
            .O(N__53639),
            .I(N__53633));
    LocalMux I__12352 (
            .O(N__53636),
            .I(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ));
    Odrv4 I__12351 (
            .O(N__53633),
            .I(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ));
    CascadeMux I__12350 (
            .O(N__53628),
            .I(N__53625));
    InMux I__12349 (
            .O(N__53625),
            .I(N__53620));
    InMux I__12348 (
            .O(N__53624),
            .I(N__53615));
    InMux I__12347 (
            .O(N__53623),
            .I(N__53615));
    LocalMux I__12346 (
            .O(N__53620),
            .I(\pid_side.un1_pid_prereg_0 ));
    LocalMux I__12345 (
            .O(N__53615),
            .I(\pid_side.un1_pid_prereg_0 ));
    InMux I__12344 (
            .O(N__53610),
            .I(N__53604));
    InMux I__12343 (
            .O(N__53609),
            .I(N__53604));
    LocalMux I__12342 (
            .O(N__53604),
            .I(\pid_side.error_d_reg_prevZ0Z_3 ));
    InMux I__12341 (
            .O(N__53601),
            .I(N__53596));
    InMux I__12340 (
            .O(N__53600),
            .I(N__53591));
    InMux I__12339 (
            .O(N__53599),
            .I(N__53591));
    LocalMux I__12338 (
            .O(N__53596),
            .I(\pid_side.un1_pid_prereg_3 ));
    LocalMux I__12337 (
            .O(N__53591),
            .I(\pid_side.un1_pid_prereg_3 ));
    CascadeMux I__12336 (
            .O(N__53586),
            .I(N__53583));
    InMux I__12335 (
            .O(N__53583),
            .I(N__53577));
    InMux I__12334 (
            .O(N__53582),
            .I(N__53577));
    LocalMux I__12333 (
            .O(N__53577),
            .I(\pid_side.error_d_reg_prevZ0Z_2 ));
    InMux I__12332 (
            .O(N__53574),
            .I(N__53570));
    InMux I__12331 (
            .O(N__53573),
            .I(N__53567));
    LocalMux I__12330 (
            .O(N__53570),
            .I(N__53564));
    LocalMux I__12329 (
            .O(N__53567),
            .I(N__53561));
    Odrv4 I__12328 (
            .O(N__53564),
            .I(\pid_side.error_d_reg_prevZ0Z_14 ));
    Odrv4 I__12327 (
            .O(N__53561),
            .I(\pid_side.error_d_reg_prevZ0Z_14 ));
    CascadeMux I__12326 (
            .O(N__53556),
            .I(\pid_side.un1_pid_prereg_47_cascade_ ));
    CascadeMux I__12325 (
            .O(N__53553),
            .I(N__53550));
    InMux I__12324 (
            .O(N__53550),
            .I(N__53547));
    LocalMux I__12323 (
            .O(N__53547),
            .I(N__53544));
    Span4Mux_h I__12322 (
            .O(N__53544),
            .I(N__53541));
    Odrv4 I__12321 (
            .O(N__53541),
            .I(\pid_side.error_d_reg_prev_esr_RNIVB6H1Z0Z_17 ));
    InMux I__12320 (
            .O(N__53538),
            .I(N__53534));
    InMux I__12319 (
            .O(N__53537),
            .I(N__53531));
    LocalMux I__12318 (
            .O(N__53534),
            .I(N__53528));
    LocalMux I__12317 (
            .O(N__53531),
            .I(N__53523));
    Span4Mux_h I__12316 (
            .O(N__53528),
            .I(N__53523));
    Odrv4 I__12315 (
            .O(N__53523),
            .I(\pid_side.error_d_reg_prevZ0Z_10 ));
    InMux I__12314 (
            .O(N__53520),
            .I(N__53517));
    LocalMux I__12313 (
            .O(N__53517),
            .I(N__53514));
    Odrv4 I__12312 (
            .O(N__53514),
            .I(\pid_side.O_1_4 ));
    CascadeMux I__12311 (
            .O(N__53511),
            .I(N__53506));
    CascadeMux I__12310 (
            .O(N__53510),
            .I(N__53503));
    InMux I__12309 (
            .O(N__53509),
            .I(N__53500));
    InMux I__12308 (
            .O(N__53506),
            .I(N__53497));
    InMux I__12307 (
            .O(N__53503),
            .I(N__53494));
    LocalMux I__12306 (
            .O(N__53500),
            .I(N__53491));
    LocalMux I__12305 (
            .O(N__53497),
            .I(N__53486));
    LocalMux I__12304 (
            .O(N__53494),
            .I(N__53486));
    Span4Mux_h I__12303 (
            .O(N__53491),
            .I(N__53483));
    Span4Mux_h I__12302 (
            .O(N__53486),
            .I(N__53480));
    Span4Mux_v I__12301 (
            .O(N__53483),
            .I(N__53475));
    Span4Mux_v I__12300 (
            .O(N__53480),
            .I(N__53475));
    Odrv4 I__12299 (
            .O(N__53475),
            .I(\pid_side.error_d_regZ0Z_0 ));
    InMux I__12298 (
            .O(N__53472),
            .I(N__53469));
    LocalMux I__12297 (
            .O(N__53469),
            .I(N__53466));
    Span4Mux_v I__12296 (
            .O(N__53466),
            .I(N__53463));
    Odrv4 I__12295 (
            .O(N__53463),
            .I(\pid_side.O_1_8 ));
    InMux I__12294 (
            .O(N__53460),
            .I(N__53451));
    InMux I__12293 (
            .O(N__53459),
            .I(N__53451));
    InMux I__12292 (
            .O(N__53458),
            .I(N__53451));
    LocalMux I__12291 (
            .O(N__53451),
            .I(N__53448));
    Odrv12 I__12290 (
            .O(N__53448),
            .I(\pid_side.error_d_regZ0Z_4 ));
    InMux I__12289 (
            .O(N__53445),
            .I(N__53442));
    LocalMux I__12288 (
            .O(N__53442),
            .I(N__53439));
    Odrv4 I__12287 (
            .O(N__53439),
            .I(\pid_side.O_1_5 ));
    InMux I__12286 (
            .O(N__53436),
            .I(N__53432));
    CascadeMux I__12285 (
            .O(N__53435),
            .I(N__53428));
    LocalMux I__12284 (
            .O(N__53432),
            .I(N__53425));
    InMux I__12283 (
            .O(N__53431),
            .I(N__53420));
    InMux I__12282 (
            .O(N__53428),
            .I(N__53420));
    Span4Mux_h I__12281 (
            .O(N__53425),
            .I(N__53415));
    LocalMux I__12280 (
            .O(N__53420),
            .I(N__53415));
    Span4Mux_v I__12279 (
            .O(N__53415),
            .I(N__53412));
    Odrv4 I__12278 (
            .O(N__53412),
            .I(\pid_side.error_d_regZ0Z_1 ));
    InMux I__12277 (
            .O(N__53409),
            .I(N__53406));
    LocalMux I__12276 (
            .O(N__53406),
            .I(N__53402));
    CascadeMux I__12275 (
            .O(N__53405),
            .I(N__53398));
    Span4Mux_v I__12274 (
            .O(N__53402),
            .I(N__53393));
    InMux I__12273 (
            .O(N__53401),
            .I(N__53390));
    InMux I__12272 (
            .O(N__53398),
            .I(N__53387));
    InMux I__12271 (
            .O(N__53397),
            .I(N__53383));
    InMux I__12270 (
            .O(N__53396),
            .I(N__53380));
    Span4Mux_h I__12269 (
            .O(N__53393),
            .I(N__53376));
    LocalMux I__12268 (
            .O(N__53390),
            .I(N__53371));
    LocalMux I__12267 (
            .O(N__53387),
            .I(N__53371));
    InMux I__12266 (
            .O(N__53386),
            .I(N__53367));
    LocalMux I__12265 (
            .O(N__53383),
            .I(N__53364));
    LocalMux I__12264 (
            .O(N__53380),
            .I(N__53361));
    InMux I__12263 (
            .O(N__53379),
            .I(N__53357));
    Span4Mux_v I__12262 (
            .O(N__53376),
            .I(N__53354));
    Span4Mux_v I__12261 (
            .O(N__53371),
            .I(N__53351));
    InMux I__12260 (
            .O(N__53370),
            .I(N__53346));
    LocalMux I__12259 (
            .O(N__53367),
            .I(N__53343));
    Span4Mux_v I__12258 (
            .O(N__53364),
            .I(N__53340));
    Span4Mux_h I__12257 (
            .O(N__53361),
            .I(N__53337));
    InMux I__12256 (
            .O(N__53360),
            .I(N__53334));
    LocalMux I__12255 (
            .O(N__53357),
            .I(N__53331));
    Span4Mux_h I__12254 (
            .O(N__53354),
            .I(N__53326));
    Span4Mux_h I__12253 (
            .O(N__53351),
            .I(N__53326));
    InMux I__12252 (
            .O(N__53350),
            .I(N__53321));
    InMux I__12251 (
            .O(N__53349),
            .I(N__53318));
    LocalMux I__12250 (
            .O(N__53346),
            .I(N__53315));
    Span4Mux_v I__12249 (
            .O(N__53343),
            .I(N__53312));
    Span4Mux_v I__12248 (
            .O(N__53340),
            .I(N__53309));
    Sp12to4 I__12247 (
            .O(N__53337),
            .I(N__53306));
    LocalMux I__12246 (
            .O(N__53334),
            .I(N__53303));
    Span4Mux_v I__12245 (
            .O(N__53331),
            .I(N__53300));
    Span4Mux_v I__12244 (
            .O(N__53326),
            .I(N__53297));
    InMux I__12243 (
            .O(N__53325),
            .I(N__53294));
    InMux I__12242 (
            .O(N__53324),
            .I(N__53291));
    LocalMux I__12241 (
            .O(N__53321),
            .I(N__53288));
    LocalMux I__12240 (
            .O(N__53318),
            .I(N__53283));
    Span4Mux_h I__12239 (
            .O(N__53315),
            .I(N__53283));
    Span4Mux_h I__12238 (
            .O(N__53312),
            .I(N__53280));
    Sp12to4 I__12237 (
            .O(N__53309),
            .I(N__53275));
    Span12Mux_v I__12236 (
            .O(N__53306),
            .I(N__53275));
    Span4Mux_h I__12235 (
            .O(N__53303),
            .I(N__53266));
    Span4Mux_h I__12234 (
            .O(N__53300),
            .I(N__53266));
    Span4Mux_v I__12233 (
            .O(N__53297),
            .I(N__53266));
    LocalMux I__12232 (
            .O(N__53294),
            .I(N__53266));
    LocalMux I__12231 (
            .O(N__53291),
            .I(uart_pc_data_4));
    Odrv12 I__12230 (
            .O(N__53288),
            .I(uart_pc_data_4));
    Odrv4 I__12229 (
            .O(N__53283),
            .I(uart_pc_data_4));
    Odrv4 I__12228 (
            .O(N__53280),
            .I(uart_pc_data_4));
    Odrv12 I__12227 (
            .O(N__53275),
            .I(uart_pc_data_4));
    Odrv4 I__12226 (
            .O(N__53266),
            .I(uart_pc_data_4));
    InMux I__12225 (
            .O(N__53253),
            .I(N__53250));
    LocalMux I__12224 (
            .O(N__53250),
            .I(N__53246));
    InMux I__12223 (
            .O(N__53249),
            .I(N__53243));
    Span4Mux_s2_h I__12222 (
            .O(N__53246),
            .I(N__53240));
    LocalMux I__12221 (
            .O(N__53243),
            .I(N__53237));
    Span4Mux_v I__12220 (
            .O(N__53240),
            .I(N__53232));
    Span4Mux_s2_h I__12219 (
            .O(N__53237),
            .I(N__53232));
    Odrv4 I__12218 (
            .O(N__53232),
            .I(xy_kd_4));
    InMux I__12217 (
            .O(N__53229),
            .I(N__53225));
    InMux I__12216 (
            .O(N__53228),
            .I(N__53221));
    LocalMux I__12215 (
            .O(N__53225),
            .I(N__53218));
    InMux I__12214 (
            .O(N__53224),
            .I(N__53215));
    LocalMux I__12213 (
            .O(N__53221),
            .I(N__53212));
    Span4Mux_h I__12212 (
            .O(N__53218),
            .I(N__53206));
    LocalMux I__12211 (
            .O(N__53215),
            .I(N__53206));
    Span4Mux_h I__12210 (
            .O(N__53212),
            .I(N__53201));
    InMux I__12209 (
            .O(N__53211),
            .I(N__53198));
    Span4Mux_v I__12208 (
            .O(N__53206),
            .I(N__53195));
    InMux I__12207 (
            .O(N__53205),
            .I(N__53192));
    InMux I__12206 (
            .O(N__53204),
            .I(N__53189));
    Span4Mux_v I__12205 (
            .O(N__53201),
            .I(N__53186));
    LocalMux I__12204 (
            .O(N__53198),
            .I(N__53181));
    Span4Mux_v I__12203 (
            .O(N__53195),
            .I(N__53178));
    LocalMux I__12202 (
            .O(N__53192),
            .I(N__53173));
    LocalMux I__12201 (
            .O(N__53189),
            .I(N__53173));
    Span4Mux_v I__12200 (
            .O(N__53186),
            .I(N__53170));
    InMux I__12199 (
            .O(N__53185),
            .I(N__53167));
    InMux I__12198 (
            .O(N__53184),
            .I(N__53164));
    Span12Mux_v I__12197 (
            .O(N__53181),
            .I(N__53161));
    Sp12to4 I__12196 (
            .O(N__53178),
            .I(N__53156));
    Span12Mux_v I__12195 (
            .O(N__53173),
            .I(N__53156));
    Span4Mux_v I__12194 (
            .O(N__53170),
            .I(N__53149));
    LocalMux I__12193 (
            .O(N__53167),
            .I(N__53149));
    LocalMux I__12192 (
            .O(N__53164),
            .I(N__53149));
    Odrv12 I__12191 (
            .O(N__53161),
            .I(uart_drone_data_6));
    Odrv12 I__12190 (
            .O(N__53156),
            .I(uart_drone_data_6));
    Odrv4 I__12189 (
            .O(N__53149),
            .I(uart_drone_data_6));
    InMux I__12188 (
            .O(N__53142),
            .I(N__53136));
    InMux I__12187 (
            .O(N__53141),
            .I(N__53136));
    LocalMux I__12186 (
            .O(N__53136),
            .I(drone_H_disp_side_14));
    CEMux I__12185 (
            .O(N__53133),
            .I(N__53130));
    LocalMux I__12184 (
            .O(N__53130),
            .I(N__53126));
    CEMux I__12183 (
            .O(N__53129),
            .I(N__53123));
    Span4Mux_v I__12182 (
            .O(N__53126),
            .I(N__53118));
    LocalMux I__12181 (
            .O(N__53123),
            .I(N__53118));
    Span4Mux_h I__12180 (
            .O(N__53118),
            .I(N__53114));
    CEMux I__12179 (
            .O(N__53117),
            .I(N__53111));
    Span4Mux_h I__12178 (
            .O(N__53114),
            .I(N__53108));
    LocalMux I__12177 (
            .O(N__53111),
            .I(N__53105));
    Span4Mux_h I__12176 (
            .O(N__53108),
            .I(N__53102));
    Span4Mux_v I__12175 (
            .O(N__53105),
            .I(N__53099));
    Odrv4 I__12174 (
            .O(N__53102),
            .I(\dron_frame_decoder_1.N_497_0 ));
    Odrv4 I__12173 (
            .O(N__53099),
            .I(\dron_frame_decoder_1.N_497_0 ));
    InMux I__12172 (
            .O(N__53094),
            .I(N__53091));
    LocalMux I__12171 (
            .O(N__53091),
            .I(N__53088));
    Span4Mux_v I__12170 (
            .O(N__53088),
            .I(N__53085));
    Odrv4 I__12169 (
            .O(N__53085),
            .I(\pid_front.O_9 ));
    InMux I__12168 (
            .O(N__53082),
            .I(N__53073));
    InMux I__12167 (
            .O(N__53081),
            .I(N__53073));
    InMux I__12166 (
            .O(N__53080),
            .I(N__53073));
    LocalMux I__12165 (
            .O(N__53073),
            .I(N__53070));
    Span4Mux_h I__12164 (
            .O(N__53070),
            .I(N__53067));
    Span4Mux_h I__12163 (
            .O(N__53067),
            .I(N__53064));
    Span4Mux_h I__12162 (
            .O(N__53064),
            .I(N__53061));
    Odrv4 I__12161 (
            .O(N__53061),
            .I(\pid_front.error_d_regZ0Z_5 ));
    InMux I__12160 (
            .O(N__53058),
            .I(N__53055));
    LocalMux I__12159 (
            .O(N__53055),
            .I(N__53051));
    InMux I__12158 (
            .O(N__53054),
            .I(N__53048));
    Odrv12 I__12157 (
            .O(N__53051),
            .I(\pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1 ));
    LocalMux I__12156 (
            .O(N__53048),
            .I(\pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1 ));
    CascadeMux I__12155 (
            .O(N__53043),
            .I(N__53040));
    InMux I__12154 (
            .O(N__53040),
            .I(N__53037));
    LocalMux I__12153 (
            .O(N__53037),
            .I(N__53034));
    Odrv12 I__12152 (
            .O(N__53034),
            .I(\pid_side.error_p_reg_esr_RNI5PH23Z0Z_1 ));
    InMux I__12151 (
            .O(N__53031),
            .I(N__53028));
    LocalMux I__12150 (
            .O(N__53028),
            .I(N__53025));
    Odrv4 I__12149 (
            .O(N__53025),
            .I(\pid_side.O_2_4 ));
    InMux I__12148 (
            .O(N__53022),
            .I(N__53013));
    InMux I__12147 (
            .O(N__53021),
            .I(N__53013));
    InMux I__12146 (
            .O(N__53020),
            .I(N__53013));
    LocalMux I__12145 (
            .O(N__53013),
            .I(\pid_side.error_p_regZ0Z_0 ));
    InMux I__12144 (
            .O(N__53010),
            .I(N__53007));
    LocalMux I__12143 (
            .O(N__53007),
            .I(N__53004));
    Span4Mux_h I__12142 (
            .O(N__53004),
            .I(N__53001));
    Odrv4 I__12141 (
            .O(N__53001),
            .I(\pid_side.state_RNINK4UZ0Z_0 ));
    InMux I__12140 (
            .O(N__52998),
            .I(N__52992));
    InMux I__12139 (
            .O(N__52997),
            .I(N__52992));
    LocalMux I__12138 (
            .O(N__52992),
            .I(\pid_side.error_p_reg_esr_RNIE47JZ0Z_9 ));
    InMux I__12137 (
            .O(N__52989),
            .I(N__52986));
    LocalMux I__12136 (
            .O(N__52986),
            .I(N__52982));
    InMux I__12135 (
            .O(N__52985),
            .I(N__52979));
    Odrv4 I__12134 (
            .O(N__52982),
            .I(\pid_side.error_d_reg_prevZ0Z_15 ));
    LocalMux I__12133 (
            .O(N__52979),
            .I(\pid_side.error_d_reg_prevZ0Z_15 ));
    InMux I__12132 (
            .O(N__52974),
            .I(N__52971));
    LocalMux I__12131 (
            .O(N__52971),
            .I(N__52966));
    InMux I__12130 (
            .O(N__52970),
            .I(N__52961));
    InMux I__12129 (
            .O(N__52969),
            .I(N__52961));
    Odrv4 I__12128 (
            .O(N__52966),
            .I(\pid_side.un1_pid_prereg_24 ));
    LocalMux I__12127 (
            .O(N__52961),
            .I(\pid_side.un1_pid_prereg_24 ));
    InMux I__12126 (
            .O(N__52956),
            .I(N__52947));
    InMux I__12125 (
            .O(N__52955),
            .I(N__52947));
    InMux I__12124 (
            .O(N__52954),
            .I(N__52947));
    LocalMux I__12123 (
            .O(N__52947),
            .I(N__52944));
    Span4Mux_v I__12122 (
            .O(N__52944),
            .I(N__52941));
    Odrv4 I__12121 (
            .O(N__52941),
            .I(\pid_side.un1_pid_prereg_48 ));
    InMux I__12120 (
            .O(N__52938),
            .I(N__52935));
    LocalMux I__12119 (
            .O(N__52935),
            .I(N__52931));
    InMux I__12118 (
            .O(N__52934),
            .I(N__52928));
    Odrv12 I__12117 (
            .O(N__52931),
            .I(\pid_side.un1_pid_prereg_36 ));
    LocalMux I__12116 (
            .O(N__52928),
            .I(\pid_side.un1_pid_prereg_36 ));
    CascadeMux I__12115 (
            .O(N__52923),
            .I(N__52920));
    InMux I__12114 (
            .O(N__52920),
            .I(N__52917));
    LocalMux I__12113 (
            .O(N__52917),
            .I(N__52914));
    Span4Mux_h I__12112 (
            .O(N__52914),
            .I(N__52911));
    Odrv4 I__12111 (
            .O(N__52911),
            .I(\pid_side.error_d_reg_prev_esr_RNIOHC23Z0Z_16 ));
    CascadeMux I__12110 (
            .O(N__52908),
            .I(N__52905));
    InMux I__12109 (
            .O(N__52905),
            .I(N__52899));
    InMux I__12108 (
            .O(N__52904),
            .I(N__52899));
    LocalMux I__12107 (
            .O(N__52899),
            .I(\pid_side.error_d_reg_prevZ0Z_18 ));
    InMux I__12106 (
            .O(N__52896),
            .I(N__52893));
    LocalMux I__12105 (
            .O(N__52893),
            .I(N__52890));
    Span4Mux_v I__12104 (
            .O(N__52890),
            .I(N__52886));
    InMux I__12103 (
            .O(N__52889),
            .I(N__52883));
    Odrv4 I__12102 (
            .O(N__52886),
            .I(\pid_side.un1_pid_prereg_47 ));
    LocalMux I__12101 (
            .O(N__52883),
            .I(\pid_side.un1_pid_prereg_47 ));
    InMux I__12100 (
            .O(N__52878),
            .I(N__52874));
    InMux I__12099 (
            .O(N__52877),
            .I(N__52871));
    LocalMux I__12098 (
            .O(N__52874),
            .I(N__52868));
    LocalMux I__12097 (
            .O(N__52871),
            .I(N__52865));
    Odrv4 I__12096 (
            .O(N__52868),
            .I(\pid_side.error_d_reg_esr_RNI76TK1Z0Z_5 ));
    Odrv4 I__12095 (
            .O(N__52865),
            .I(\pid_side.error_d_reg_esr_RNI76TK1Z0Z_5 ));
    CascadeMux I__12094 (
            .O(N__52860),
            .I(\pid_side.un1_pid_prereg_40_0_cascade_ ));
    CascadeMux I__12093 (
            .O(N__52857),
            .I(N__52854));
    InMux I__12092 (
            .O(N__52854),
            .I(N__52851));
    LocalMux I__12091 (
            .O(N__52851),
            .I(N__52848));
    Odrv4 I__12090 (
            .O(N__52848),
            .I(\pid_side.error_d_reg_esr_RNI86Q93Z0Z_5 ));
    InMux I__12089 (
            .O(N__52845),
            .I(N__52839));
    InMux I__12088 (
            .O(N__52844),
            .I(N__52839));
    LocalMux I__12087 (
            .O(N__52839),
            .I(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ));
    CascadeMux I__12086 (
            .O(N__52836),
            .I(\pid_side.un1_pid_prereg_17_cascade_ ));
    InMux I__12085 (
            .O(N__52833),
            .I(N__52830));
    LocalMux I__12084 (
            .O(N__52830),
            .I(N__52827));
    Odrv4 I__12083 (
            .O(N__52827),
            .I(\pid_side.error_p_reg_esr_RNI10TK1Z0Z_3 ));
    CascadeMux I__12082 (
            .O(N__52824),
            .I(N__52821));
    InMux I__12081 (
            .O(N__52821),
            .I(N__52815));
    InMux I__12080 (
            .O(N__52820),
            .I(N__52815));
    LocalMux I__12079 (
            .O(N__52815),
            .I(\pid_side.error_d_reg_prevZ0Z_4 ));
    InMux I__12078 (
            .O(N__52812),
            .I(N__52806));
    InMux I__12077 (
            .O(N__52811),
            .I(N__52806));
    LocalMux I__12076 (
            .O(N__52806),
            .I(\pid_side.un1_pid_prereg_17 ));
    CascadeMux I__12075 (
            .O(N__52803),
            .I(N__52800));
    InMux I__12074 (
            .O(N__52800),
            .I(N__52797));
    LocalMux I__12073 (
            .O(N__52797),
            .I(N__52794));
    Odrv4 I__12072 (
            .O(N__52794),
            .I(\pid_side.error_p_reg_esr_RNISPP93Z0Z_2 ));
    InMux I__12071 (
            .O(N__52791),
            .I(N__52788));
    LocalMux I__12070 (
            .O(N__52788),
            .I(N__52785));
    Span4Mux_v I__12069 (
            .O(N__52785),
            .I(N__52782));
    Odrv4 I__12068 (
            .O(N__52782),
            .I(\pid_side.O_2_9 ));
    CascadeMux I__12067 (
            .O(N__52779),
            .I(N__52776));
    InMux I__12066 (
            .O(N__52776),
            .I(N__52773));
    LocalMux I__12065 (
            .O(N__52773),
            .I(drone_H_disp_side_i_13));
    InMux I__12064 (
            .O(N__52770),
            .I(N__52766));
    InMux I__12063 (
            .O(N__52769),
            .I(N__52763));
    LocalMux I__12062 (
            .O(N__52766),
            .I(N__52760));
    LocalMux I__12061 (
            .O(N__52763),
            .I(N__52757));
    Span12Mux_s4_h I__12060 (
            .O(N__52760),
            .I(N__52754));
    Span4Mux_s3_h I__12059 (
            .O(N__52757),
            .I(N__52751));
    Odrv12 I__12058 (
            .O(N__52754),
            .I(\pid_side.error_14 ));
    Odrv4 I__12057 (
            .O(N__52751),
            .I(\pid_side.error_14 ));
    InMux I__12056 (
            .O(N__52746),
            .I(\pid_side.error_cry_9 ));
    InMux I__12055 (
            .O(N__52743),
            .I(\pid_side.error_cry_10 ));
    InMux I__12054 (
            .O(N__52740),
            .I(N__52737));
    LocalMux I__12053 (
            .O(N__52737),
            .I(N__52733));
    InMux I__12052 (
            .O(N__52736),
            .I(N__52730));
    Span4Mux_s3_h I__12051 (
            .O(N__52733),
            .I(N__52727));
    LocalMux I__12050 (
            .O(N__52730),
            .I(N__52724));
    Span4Mux_v I__12049 (
            .O(N__52727),
            .I(N__52721));
    Span4Mux_s3_h I__12048 (
            .O(N__52724),
            .I(N__52718));
    Odrv4 I__12047 (
            .O(N__52721),
            .I(\pid_side.error_15 ));
    Odrv4 I__12046 (
            .O(N__52718),
            .I(\pid_side.error_15 ));
    InMux I__12045 (
            .O(N__52713),
            .I(N__52710));
    LocalMux I__12044 (
            .O(N__52710),
            .I(N__52705));
    InMux I__12043 (
            .O(N__52709),
            .I(N__52702));
    InMux I__12042 (
            .O(N__52708),
            .I(N__52699));
    Span4Mux_h I__12041 (
            .O(N__52705),
            .I(N__52694));
    LocalMux I__12040 (
            .O(N__52702),
            .I(N__52694));
    LocalMux I__12039 (
            .O(N__52699),
            .I(N__52690));
    Span4Mux_v I__12038 (
            .O(N__52694),
            .I(N__52687));
    InMux I__12037 (
            .O(N__52693),
            .I(N__52684));
    Span4Mux_v I__12036 (
            .O(N__52690),
            .I(N__52680));
    Span4Mux_h I__12035 (
            .O(N__52687),
            .I(N__52676));
    LocalMux I__12034 (
            .O(N__52684),
            .I(N__52673));
    InMux I__12033 (
            .O(N__52683),
            .I(N__52670));
    Span4Mux_h I__12032 (
            .O(N__52680),
            .I(N__52667));
    InMux I__12031 (
            .O(N__52679),
            .I(N__52664));
    Span4Mux_h I__12030 (
            .O(N__52676),
            .I(N__52656));
    Span4Mux_v I__12029 (
            .O(N__52673),
            .I(N__52656));
    LocalMux I__12028 (
            .O(N__52670),
            .I(N__52656));
    Span4Mux_v I__12027 (
            .O(N__52667),
            .I(N__52653));
    LocalMux I__12026 (
            .O(N__52664),
            .I(N__52650));
    CascadeMux I__12025 (
            .O(N__52663),
            .I(N__52646));
    Span4Mux_v I__12024 (
            .O(N__52656),
            .I(N__52643));
    Span4Mux_v I__12023 (
            .O(N__52653),
            .I(N__52638));
    Span4Mux_h I__12022 (
            .O(N__52650),
            .I(N__52638));
    InMux I__12021 (
            .O(N__52649),
            .I(N__52635));
    InMux I__12020 (
            .O(N__52646),
            .I(N__52632));
    Span4Mux_v I__12019 (
            .O(N__52643),
            .I(N__52629));
    Span4Mux_v I__12018 (
            .O(N__52638),
            .I(N__52626));
    LocalMux I__12017 (
            .O(N__52635),
            .I(N__52621));
    LocalMux I__12016 (
            .O(N__52632),
            .I(N__52621));
    Odrv4 I__12015 (
            .O(N__52629),
            .I(uart_drone_data_3));
    Odrv4 I__12014 (
            .O(N__52626),
            .I(uart_drone_data_3));
    Odrv4 I__12013 (
            .O(N__52621),
            .I(uart_drone_data_3));
    InMux I__12012 (
            .O(N__52614),
            .I(N__52608));
    InMux I__12011 (
            .O(N__52613),
            .I(N__52608));
    LocalMux I__12010 (
            .O(N__52608),
            .I(drone_H_disp_side_11));
    InMux I__12009 (
            .O(N__52605),
            .I(N__52602));
    LocalMux I__12008 (
            .O(N__52602),
            .I(N__52599));
    Span4Mux_v I__12007 (
            .O(N__52599),
            .I(N__52594));
    InMux I__12006 (
            .O(N__52598),
            .I(N__52591));
    InMux I__12005 (
            .O(N__52597),
            .I(N__52587));
    Span4Mux_h I__12004 (
            .O(N__52594),
            .I(N__52583));
    LocalMux I__12003 (
            .O(N__52591),
            .I(N__52580));
    InMux I__12002 (
            .O(N__52590),
            .I(N__52577));
    LocalMux I__12001 (
            .O(N__52587),
            .I(N__52573));
    InMux I__12000 (
            .O(N__52586),
            .I(N__52570));
    Span4Mux_h I__11999 (
            .O(N__52583),
            .I(N__52565));
    Span4Mux_v I__11998 (
            .O(N__52580),
            .I(N__52565));
    LocalMux I__11997 (
            .O(N__52577),
            .I(N__52562));
    InMux I__11996 (
            .O(N__52576),
            .I(N__52559));
    Span4Mux_h I__11995 (
            .O(N__52573),
            .I(N__52556));
    LocalMux I__11994 (
            .O(N__52570),
            .I(N__52553));
    Span4Mux_h I__11993 (
            .O(N__52565),
            .I(N__52546));
    Span4Mux_v I__11992 (
            .O(N__52562),
            .I(N__52546));
    LocalMux I__11991 (
            .O(N__52559),
            .I(N__52546));
    Span4Mux_v I__11990 (
            .O(N__52556),
            .I(N__52543));
    Sp12to4 I__11989 (
            .O(N__52553),
            .I(N__52538));
    Span4Mux_v I__11988 (
            .O(N__52546),
            .I(N__52535));
    Span4Mux_v I__11987 (
            .O(N__52543),
            .I(N__52532));
    InMux I__11986 (
            .O(N__52542),
            .I(N__52529));
    InMux I__11985 (
            .O(N__52541),
            .I(N__52526));
    Span12Mux_v I__11984 (
            .O(N__52538),
            .I(N__52523));
    Span4Mux_v I__11983 (
            .O(N__52535),
            .I(N__52520));
    Span4Mux_v I__11982 (
            .O(N__52532),
            .I(N__52513));
    LocalMux I__11981 (
            .O(N__52529),
            .I(N__52513));
    LocalMux I__11980 (
            .O(N__52526),
            .I(N__52513));
    Odrv12 I__11979 (
            .O(N__52523),
            .I(uart_drone_data_4));
    Odrv4 I__11978 (
            .O(N__52520),
            .I(uart_drone_data_4));
    Odrv4 I__11977 (
            .O(N__52513),
            .I(uart_drone_data_4));
    CascadeMux I__11976 (
            .O(N__52506),
            .I(N__52503));
    InMux I__11975 (
            .O(N__52503),
            .I(N__52498));
    InMux I__11974 (
            .O(N__52502),
            .I(N__52493));
    InMux I__11973 (
            .O(N__52501),
            .I(N__52493));
    LocalMux I__11972 (
            .O(N__52498),
            .I(drone_H_disp_side_12));
    LocalMux I__11971 (
            .O(N__52493),
            .I(drone_H_disp_side_12));
    InMux I__11970 (
            .O(N__52488),
            .I(N__52485));
    LocalMux I__11969 (
            .O(N__52485),
            .I(N__52481));
    InMux I__11968 (
            .O(N__52484),
            .I(N__52478));
    Span4Mux_v I__11967 (
            .O(N__52481),
            .I(N__52472));
    LocalMux I__11966 (
            .O(N__52478),
            .I(N__52472));
    InMux I__11965 (
            .O(N__52477),
            .I(N__52469));
    Span4Mux_h I__11964 (
            .O(N__52472),
            .I(N__52464));
    LocalMux I__11963 (
            .O(N__52469),
            .I(N__52461));
    InMux I__11962 (
            .O(N__52468),
            .I(N__52458));
    InMux I__11961 (
            .O(N__52467),
            .I(N__52454));
    Span4Mux_h I__11960 (
            .O(N__52464),
            .I(N__52449));
    Span4Mux_v I__11959 (
            .O(N__52461),
            .I(N__52449));
    LocalMux I__11958 (
            .O(N__52458),
            .I(N__52446));
    InMux I__11957 (
            .O(N__52457),
            .I(N__52443));
    LocalMux I__11956 (
            .O(N__52454),
            .I(N__52440));
    Span4Mux_h I__11955 (
            .O(N__52449),
            .I(N__52433));
    Span4Mux_v I__11954 (
            .O(N__52446),
            .I(N__52433));
    LocalMux I__11953 (
            .O(N__52443),
            .I(N__52433));
    Sp12to4 I__11952 (
            .O(N__52440),
            .I(N__52430));
    Span4Mux_v I__11951 (
            .O(N__52433),
            .I(N__52427));
    Span12Mux_v I__11950 (
            .O(N__52430),
            .I(N__52423));
    Span4Mux_v I__11949 (
            .O(N__52427),
            .I(N__52420));
    InMux I__11948 (
            .O(N__52426),
            .I(N__52417));
    Odrv12 I__11947 (
            .O(N__52423),
            .I(uart_drone_data_5));
    Odrv4 I__11946 (
            .O(N__52420),
            .I(uart_drone_data_5));
    LocalMux I__11945 (
            .O(N__52417),
            .I(uart_drone_data_5));
    CascadeMux I__11944 (
            .O(N__52410),
            .I(N__52407));
    InMux I__11943 (
            .O(N__52407),
            .I(N__52403));
    InMux I__11942 (
            .O(N__52406),
            .I(N__52400));
    LocalMux I__11941 (
            .O(N__52403),
            .I(drone_H_disp_side_13));
    LocalMux I__11940 (
            .O(N__52400),
            .I(drone_H_disp_side_13));
    InMux I__11939 (
            .O(N__52395),
            .I(N__52392));
    LocalMux I__11938 (
            .O(N__52392),
            .I(N__52388));
    InMux I__11937 (
            .O(N__52391),
            .I(N__52385));
    Span4Mux_v I__11936 (
            .O(N__52388),
            .I(N__52379));
    LocalMux I__11935 (
            .O(N__52385),
            .I(N__52379));
    InMux I__11934 (
            .O(N__52384),
            .I(N__52375));
    Span4Mux_v I__11933 (
            .O(N__52379),
            .I(N__52371));
    InMux I__11932 (
            .O(N__52378),
            .I(N__52368));
    LocalMux I__11931 (
            .O(N__52375),
            .I(N__52365));
    InMux I__11930 (
            .O(N__52374),
            .I(N__52362));
    Span4Mux_h I__11929 (
            .O(N__52371),
            .I(N__52356));
    LocalMux I__11928 (
            .O(N__52368),
            .I(N__52356));
    Span4Mux_h I__11927 (
            .O(N__52365),
            .I(N__52351));
    LocalMux I__11926 (
            .O(N__52362),
            .I(N__52351));
    InMux I__11925 (
            .O(N__52361),
            .I(N__52348));
    Span4Mux_v I__11924 (
            .O(N__52356),
            .I(N__52344));
    Sp12to4 I__11923 (
            .O(N__52351),
            .I(N__52341));
    LocalMux I__11922 (
            .O(N__52348),
            .I(N__52338));
    CascadeMux I__11921 (
            .O(N__52347),
            .I(N__52335));
    Span4Mux_v I__11920 (
            .O(N__52344),
            .I(N__52332));
    Span12Mux_v I__11919 (
            .O(N__52341),
            .I(N__52327));
    Span12Mux_v I__11918 (
            .O(N__52338),
            .I(N__52327));
    InMux I__11917 (
            .O(N__52335),
            .I(N__52324));
    Odrv4 I__11916 (
            .O(N__52332),
            .I(uart_drone_data_7));
    Odrv12 I__11915 (
            .O(N__52327),
            .I(uart_drone_data_7));
    LocalMux I__11914 (
            .O(N__52324),
            .I(uart_drone_data_7));
    InMux I__11913 (
            .O(N__52317),
            .I(N__52314));
    LocalMux I__11912 (
            .O(N__52314),
            .I(drone_H_disp_side_15));
    InMux I__11911 (
            .O(N__52311),
            .I(N__52308));
    LocalMux I__11910 (
            .O(N__52308),
            .I(N__52304));
    InMux I__11909 (
            .O(N__52307),
            .I(N__52301));
    Span4Mux_v I__11908 (
            .O(N__52304),
            .I(N__52295));
    LocalMux I__11907 (
            .O(N__52301),
            .I(N__52295));
    InMux I__11906 (
            .O(N__52300),
            .I(N__52292));
    Span4Mux_v I__11905 (
            .O(N__52295),
            .I(N__52288));
    LocalMux I__11904 (
            .O(N__52292),
            .I(N__52285));
    InMux I__11903 (
            .O(N__52291),
            .I(N__52282));
    Span4Mux_h I__11902 (
            .O(N__52288),
            .I(N__52279));
    Span4Mux_v I__11901 (
            .O(N__52285),
            .I(N__52274));
    LocalMux I__11900 (
            .O(N__52282),
            .I(N__52274));
    Span4Mux_h I__11899 (
            .O(N__52279),
            .I(N__52268));
    Span4Mux_v I__11898 (
            .O(N__52274),
            .I(N__52268));
    InMux I__11897 (
            .O(N__52273),
            .I(N__52265));
    Span4Mux_h I__11896 (
            .O(N__52268),
            .I(N__52260));
    LocalMux I__11895 (
            .O(N__52265),
            .I(N__52260));
    Span4Mux_v I__11894 (
            .O(N__52260),
            .I(N__52256));
    InMux I__11893 (
            .O(N__52259),
            .I(N__52253));
    Sp12to4 I__11892 (
            .O(N__52256),
            .I(N__52248));
    LocalMux I__11891 (
            .O(N__52253),
            .I(N__52248));
    Span12Mux_s10_h I__11890 (
            .O(N__52248),
            .I(N__52244));
    InMux I__11889 (
            .O(N__52247),
            .I(N__52241));
    Odrv12 I__11888 (
            .O(N__52244),
            .I(uart_drone_data_0));
    LocalMux I__11887 (
            .O(N__52241),
            .I(uart_drone_data_0));
    InMux I__11886 (
            .O(N__52236),
            .I(N__52233));
    LocalMux I__11885 (
            .O(N__52233),
            .I(\dron_frame_decoder_1.drone_H_disp_side_8 ));
    InMux I__11884 (
            .O(N__52230),
            .I(N__52227));
    LocalMux I__11883 (
            .O(N__52227),
            .I(N__52224));
    Span4Mux_h I__11882 (
            .O(N__52224),
            .I(N__52221));
    Odrv4 I__11881 (
            .O(N__52221),
            .I(\pid_front.O_10 ));
    InMux I__11880 (
            .O(N__52218),
            .I(N__52213));
    InMux I__11879 (
            .O(N__52217),
            .I(N__52208));
    InMux I__11878 (
            .O(N__52216),
            .I(N__52208));
    LocalMux I__11877 (
            .O(N__52213),
            .I(N__52203));
    LocalMux I__11876 (
            .O(N__52208),
            .I(N__52203));
    Span4Mux_h I__11875 (
            .O(N__52203),
            .I(N__52200));
    Span4Mux_h I__11874 (
            .O(N__52200),
            .I(N__52197));
    Span4Mux_h I__11873 (
            .O(N__52197),
            .I(N__52194));
    Odrv4 I__11872 (
            .O(N__52194),
            .I(\pid_front.error_d_regZ0Z_6 ));
    InMux I__11871 (
            .O(N__52191),
            .I(N__52188));
    LocalMux I__11870 (
            .O(N__52188),
            .I(drone_H_disp_side_i_6));
    CascadeMux I__11869 (
            .O(N__52185),
            .I(N__52182));
    InMux I__11868 (
            .O(N__52182),
            .I(N__52179));
    LocalMux I__11867 (
            .O(N__52179),
            .I(N__52176));
    Odrv4 I__11866 (
            .O(N__52176),
            .I(side_command_2));
    InMux I__11865 (
            .O(N__52173),
            .I(N__52170));
    LocalMux I__11864 (
            .O(N__52170),
            .I(N__52167));
    Span4Mux_s3_h I__11863 (
            .O(N__52167),
            .I(N__52163));
    InMux I__11862 (
            .O(N__52166),
            .I(N__52160));
    Span4Mux_v I__11861 (
            .O(N__52163),
            .I(N__52157));
    LocalMux I__11860 (
            .O(N__52160),
            .I(N__52154));
    Odrv4 I__11859 (
            .O(N__52157),
            .I(\pid_side.error_6 ));
    Odrv12 I__11858 (
            .O(N__52154),
            .I(\pid_side.error_6 ));
    InMux I__11857 (
            .O(N__52149),
            .I(\pid_side.error_cry_1_0 ));
    InMux I__11856 (
            .O(N__52146),
            .I(N__52143));
    LocalMux I__11855 (
            .O(N__52143),
            .I(drone_H_disp_side_i_7));
    CascadeMux I__11854 (
            .O(N__52140),
            .I(N__52137));
    InMux I__11853 (
            .O(N__52137),
            .I(N__52134));
    LocalMux I__11852 (
            .O(N__52134),
            .I(side_command_3));
    InMux I__11851 (
            .O(N__52131),
            .I(N__52128));
    LocalMux I__11850 (
            .O(N__52128),
            .I(N__52124));
    InMux I__11849 (
            .O(N__52127),
            .I(N__52121));
    Span12Mux_s4_h I__11848 (
            .O(N__52124),
            .I(N__52118));
    LocalMux I__11847 (
            .O(N__52121),
            .I(N__52115));
    Odrv12 I__11846 (
            .O(N__52118),
            .I(\pid_side.error_7 ));
    Odrv12 I__11845 (
            .O(N__52115),
            .I(\pid_side.error_7 ));
    InMux I__11844 (
            .O(N__52110),
            .I(\pid_side.error_cry_2_0 ));
    InMux I__11843 (
            .O(N__52107),
            .I(N__52104));
    LocalMux I__11842 (
            .O(N__52104),
            .I(drone_H_disp_side_i_8));
    CascadeMux I__11841 (
            .O(N__52101),
            .I(N__52098));
    InMux I__11840 (
            .O(N__52098),
            .I(N__52095));
    LocalMux I__11839 (
            .O(N__52095),
            .I(N__52092));
    Span4Mux_h I__11838 (
            .O(N__52092),
            .I(N__52089));
    Odrv4 I__11837 (
            .O(N__52089),
            .I(side_command_4));
    InMux I__11836 (
            .O(N__52086),
            .I(N__52083));
    LocalMux I__11835 (
            .O(N__52083),
            .I(N__52079));
    InMux I__11834 (
            .O(N__52082),
            .I(N__52076));
    Span4Mux_v I__11833 (
            .O(N__52079),
            .I(N__52071));
    LocalMux I__11832 (
            .O(N__52076),
            .I(N__52071));
    Span4Mux_v I__11831 (
            .O(N__52071),
            .I(N__52068));
    Odrv4 I__11830 (
            .O(N__52068),
            .I(\pid_side.error_8 ));
    InMux I__11829 (
            .O(N__52065),
            .I(bfn_21_18_0_));
    InMux I__11828 (
            .O(N__52062),
            .I(N__52059));
    LocalMux I__11827 (
            .O(N__52059),
            .I(N__52056));
    Span4Mux_v I__11826 (
            .O(N__52056),
            .I(N__52053));
    Span4Mux_h I__11825 (
            .O(N__52053),
            .I(N__52050));
    Span4Mux_h I__11824 (
            .O(N__52050),
            .I(N__52047));
    Odrv4 I__11823 (
            .O(N__52047),
            .I(drone_H_disp_side_i_9));
    CascadeMux I__11822 (
            .O(N__52044),
            .I(N__52041));
    InMux I__11821 (
            .O(N__52041),
            .I(N__52038));
    LocalMux I__11820 (
            .O(N__52038),
            .I(N__52035));
    Odrv4 I__11819 (
            .O(N__52035),
            .I(side_command_5));
    InMux I__11818 (
            .O(N__52032),
            .I(N__52029));
    LocalMux I__11817 (
            .O(N__52029),
            .I(N__52025));
    InMux I__11816 (
            .O(N__52028),
            .I(N__52022));
    Span4Mux_v I__11815 (
            .O(N__52025),
            .I(N__52017));
    LocalMux I__11814 (
            .O(N__52022),
            .I(N__52017));
    Span4Mux_v I__11813 (
            .O(N__52017),
            .I(N__52014));
    Odrv4 I__11812 (
            .O(N__52014),
            .I(\pid_side.error_9 ));
    InMux I__11811 (
            .O(N__52011),
            .I(\pid_side.error_cry_4 ));
    InMux I__11810 (
            .O(N__52008),
            .I(N__52005));
    LocalMux I__11809 (
            .O(N__52005),
            .I(N__52002));
    Span12Mux_s6_h I__11808 (
            .O(N__52002),
            .I(N__51999));
    Odrv12 I__11807 (
            .O(N__51999),
            .I(drone_H_disp_side_i_10));
    CascadeMux I__11806 (
            .O(N__51996),
            .I(N__51993));
    InMux I__11805 (
            .O(N__51993),
            .I(N__51990));
    LocalMux I__11804 (
            .O(N__51990),
            .I(N__51987));
    Span4Mux_h I__11803 (
            .O(N__51987),
            .I(N__51984));
    Odrv4 I__11802 (
            .O(N__51984),
            .I(side_command_6));
    InMux I__11801 (
            .O(N__51981),
            .I(N__51978));
    LocalMux I__11800 (
            .O(N__51978),
            .I(N__51974));
    InMux I__11799 (
            .O(N__51977),
            .I(N__51971));
    Span4Mux_v I__11798 (
            .O(N__51974),
            .I(N__51968));
    LocalMux I__11797 (
            .O(N__51971),
            .I(N__51965));
    Span4Mux_h I__11796 (
            .O(N__51968),
            .I(N__51962));
    Span4Mux_s3_h I__11795 (
            .O(N__51965),
            .I(N__51959));
    Odrv4 I__11794 (
            .O(N__51962),
            .I(\pid_side.error_10 ));
    Odrv4 I__11793 (
            .O(N__51959),
            .I(\pid_side.error_10 ));
    InMux I__11792 (
            .O(N__51954),
            .I(\pid_side.error_cry_5 ));
    InMux I__11791 (
            .O(N__51951),
            .I(N__51948));
    LocalMux I__11790 (
            .O(N__51948),
            .I(\pid_side.error_axbZ0Z_7 ));
    InMux I__11789 (
            .O(N__51945),
            .I(N__51942));
    LocalMux I__11788 (
            .O(N__51942),
            .I(N__51938));
    InMux I__11787 (
            .O(N__51941),
            .I(N__51935));
    Span4Mux_v I__11786 (
            .O(N__51938),
            .I(N__51932));
    LocalMux I__11785 (
            .O(N__51935),
            .I(N__51929));
    Span4Mux_h I__11784 (
            .O(N__51932),
            .I(N__51926));
    Span4Mux_s3_h I__11783 (
            .O(N__51929),
            .I(N__51923));
    Odrv4 I__11782 (
            .O(N__51926),
            .I(\pid_side.error_11 ));
    Odrv4 I__11781 (
            .O(N__51923),
            .I(\pid_side.error_11 ));
    InMux I__11780 (
            .O(N__51918),
            .I(\pid_side.error_cry_6 ));
    InMux I__11779 (
            .O(N__51915),
            .I(N__51912));
    LocalMux I__11778 (
            .O(N__51912),
            .I(\pid_side.error_axb_8_l_ofxZ0 ));
    InMux I__11777 (
            .O(N__51909),
            .I(N__51906));
    LocalMux I__11776 (
            .O(N__51906),
            .I(N__51902));
    InMux I__11775 (
            .O(N__51905),
            .I(N__51899));
    Span4Mux_s3_h I__11774 (
            .O(N__51902),
            .I(N__51896));
    LocalMux I__11773 (
            .O(N__51899),
            .I(N__51893));
    Span4Mux_v I__11772 (
            .O(N__51896),
            .I(N__51890));
    Span4Mux_s3_h I__11771 (
            .O(N__51893),
            .I(N__51887));
    Odrv4 I__11770 (
            .O(N__51890),
            .I(\pid_side.error_12 ));
    Odrv4 I__11769 (
            .O(N__51887),
            .I(\pid_side.error_12 ));
    InMux I__11768 (
            .O(N__51882),
            .I(\pid_side.error_cry_7 ));
    InMux I__11767 (
            .O(N__51879),
            .I(N__51876));
    LocalMux I__11766 (
            .O(N__51876),
            .I(drone_H_disp_side_i_12));
    InMux I__11765 (
            .O(N__51873),
            .I(N__51870));
    LocalMux I__11764 (
            .O(N__51870),
            .I(N__51866));
    InMux I__11763 (
            .O(N__51869),
            .I(N__51863));
    Span4Mux_s3_h I__11762 (
            .O(N__51866),
            .I(N__51860));
    LocalMux I__11761 (
            .O(N__51863),
            .I(N__51857));
    Span4Mux_v I__11760 (
            .O(N__51860),
            .I(N__51854));
    Span4Mux_s3_h I__11759 (
            .O(N__51857),
            .I(N__51851));
    Odrv4 I__11758 (
            .O(N__51854),
            .I(\pid_side.error_13 ));
    Odrv4 I__11757 (
            .O(N__51851),
            .I(\pid_side.error_13 ));
    InMux I__11756 (
            .O(N__51846),
            .I(\pid_side.error_cry_8 ));
    InMux I__11755 (
            .O(N__51843),
            .I(N__51837));
    InMux I__11754 (
            .O(N__51842),
            .I(N__51837));
    LocalMux I__11753 (
            .O(N__51837),
            .I(\pid_side.error_d_reg_prevZ0Z_19 ));
    CascadeMux I__11752 (
            .O(N__51834),
            .I(N__51830));
    InMux I__11751 (
            .O(N__51833),
            .I(N__51827));
    InMux I__11750 (
            .O(N__51830),
            .I(N__51823));
    LocalMux I__11749 (
            .O(N__51827),
            .I(N__51820));
    InMux I__11748 (
            .O(N__51826),
            .I(N__51817));
    LocalMux I__11747 (
            .O(N__51823),
            .I(\pid_side.un1_pid_prereg_57 ));
    Odrv4 I__11746 (
            .O(N__51820),
            .I(\pid_side.un1_pid_prereg_57 ));
    LocalMux I__11745 (
            .O(N__51817),
            .I(\pid_side.un1_pid_prereg_57 ));
    CEMux I__11744 (
            .O(N__51810),
            .I(N__51806));
    CEMux I__11743 (
            .O(N__51809),
            .I(N__51803));
    LocalMux I__11742 (
            .O(N__51806),
            .I(N__51800));
    LocalMux I__11741 (
            .O(N__51803),
            .I(N__51797));
    Span4Mux_h I__11740 (
            .O(N__51800),
            .I(N__51794));
    Span4Mux_h I__11739 (
            .O(N__51797),
            .I(N__51789));
    Span4Mux_h I__11738 (
            .O(N__51794),
            .I(N__51789));
    Odrv4 I__11737 (
            .O(N__51789),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    InMux I__11736 (
            .O(N__51786),
            .I(N__51783));
    LocalMux I__11735 (
            .O(N__51783),
            .I(N__51780));
    Span4Mux_v I__11734 (
            .O(N__51780),
            .I(N__51776));
    InMux I__11733 (
            .O(N__51779),
            .I(N__51773));
    Span4Mux_h I__11732 (
            .O(N__51776),
            .I(N__51769));
    LocalMux I__11731 (
            .O(N__51773),
            .I(N__51766));
    InMux I__11730 (
            .O(N__51772),
            .I(N__51763));
    Odrv4 I__11729 (
            .O(N__51769),
            .I(drone_H_disp_side_0));
    Odrv12 I__11728 (
            .O(N__51766),
            .I(drone_H_disp_side_0));
    LocalMux I__11727 (
            .O(N__51763),
            .I(drone_H_disp_side_0));
    InMux I__11726 (
            .O(N__51756),
            .I(N__51753));
    LocalMux I__11725 (
            .O(N__51753),
            .I(\pid_side.error_axb_0 ));
    InMux I__11724 (
            .O(N__51750),
            .I(N__51747));
    LocalMux I__11723 (
            .O(N__51747),
            .I(\pid_side.error_axbZ0Z_1 ));
    InMux I__11722 (
            .O(N__51744),
            .I(N__51741));
    LocalMux I__11721 (
            .O(N__51741),
            .I(N__51737));
    InMux I__11720 (
            .O(N__51740),
            .I(N__51734));
    Span4Mux_v I__11719 (
            .O(N__51737),
            .I(N__51731));
    LocalMux I__11718 (
            .O(N__51734),
            .I(N__51728));
    Span4Mux_h I__11717 (
            .O(N__51731),
            .I(N__51725));
    Span4Mux_s1_h I__11716 (
            .O(N__51728),
            .I(N__51722));
    Odrv4 I__11715 (
            .O(N__51725),
            .I(\pid_side.error_1 ));
    Odrv4 I__11714 (
            .O(N__51722),
            .I(\pid_side.error_1 ));
    InMux I__11713 (
            .O(N__51717),
            .I(\pid_side.error_cry_0 ));
    InMux I__11712 (
            .O(N__51714),
            .I(N__51711));
    LocalMux I__11711 (
            .O(N__51711),
            .I(\pid_side.error_axbZ0Z_2 ));
    InMux I__11710 (
            .O(N__51708),
            .I(N__51705));
    LocalMux I__11709 (
            .O(N__51705),
            .I(N__51701));
    InMux I__11708 (
            .O(N__51704),
            .I(N__51698));
    Span4Mux_v I__11707 (
            .O(N__51701),
            .I(N__51695));
    LocalMux I__11706 (
            .O(N__51698),
            .I(N__51692));
    Span4Mux_h I__11705 (
            .O(N__51695),
            .I(N__51689));
    Span4Mux_s1_h I__11704 (
            .O(N__51692),
            .I(N__51686));
    Odrv4 I__11703 (
            .O(N__51689),
            .I(\pid_side.error_2 ));
    Odrv4 I__11702 (
            .O(N__51686),
            .I(\pid_side.error_2 ));
    InMux I__11701 (
            .O(N__51681),
            .I(\pid_side.error_cry_1 ));
    InMux I__11700 (
            .O(N__51678),
            .I(N__51675));
    LocalMux I__11699 (
            .O(N__51675),
            .I(\pid_side.error_axbZ0Z_3 ));
    InMux I__11698 (
            .O(N__51672),
            .I(N__51669));
    LocalMux I__11697 (
            .O(N__51669),
            .I(N__51666));
    Span4Mux_v I__11696 (
            .O(N__51666),
            .I(N__51662));
    InMux I__11695 (
            .O(N__51665),
            .I(N__51659));
    Span4Mux_v I__11694 (
            .O(N__51662),
            .I(N__51654));
    LocalMux I__11693 (
            .O(N__51659),
            .I(N__51654));
    Span4Mux_s0_h I__11692 (
            .O(N__51654),
            .I(N__51651));
    Odrv4 I__11691 (
            .O(N__51651),
            .I(\pid_side.error_3 ));
    InMux I__11690 (
            .O(N__51648),
            .I(\pid_side.error_cry_2 ));
    InMux I__11689 (
            .O(N__51645),
            .I(N__51642));
    LocalMux I__11688 (
            .O(N__51642),
            .I(drone_H_disp_side_i_4));
    CascadeMux I__11687 (
            .O(N__51639),
            .I(N__51636));
    InMux I__11686 (
            .O(N__51636),
            .I(N__51633));
    LocalMux I__11685 (
            .O(N__51633),
            .I(N__51630));
    Odrv4 I__11684 (
            .O(N__51630),
            .I(side_command_0));
    InMux I__11683 (
            .O(N__51627),
            .I(N__51624));
    LocalMux I__11682 (
            .O(N__51624),
            .I(N__51621));
    Span4Mux_s3_h I__11681 (
            .O(N__51621),
            .I(N__51617));
    InMux I__11680 (
            .O(N__51620),
            .I(N__51614));
    Span4Mux_v I__11679 (
            .O(N__51617),
            .I(N__51611));
    LocalMux I__11678 (
            .O(N__51614),
            .I(N__51608));
    Odrv4 I__11677 (
            .O(N__51611),
            .I(\pid_side.error_4 ));
    Odrv12 I__11676 (
            .O(N__51608),
            .I(\pid_side.error_4 ));
    InMux I__11675 (
            .O(N__51603),
            .I(\pid_side.error_cry_3 ));
    InMux I__11674 (
            .O(N__51600),
            .I(N__51597));
    LocalMux I__11673 (
            .O(N__51597),
            .I(N__51594));
    Odrv4 I__11672 (
            .O(N__51594),
            .I(drone_H_disp_side_i_5));
    CascadeMux I__11671 (
            .O(N__51591),
            .I(N__51588));
    InMux I__11670 (
            .O(N__51588),
            .I(N__51585));
    LocalMux I__11669 (
            .O(N__51585),
            .I(side_command_1));
    InMux I__11668 (
            .O(N__51582),
            .I(N__51579));
    LocalMux I__11667 (
            .O(N__51579),
            .I(N__51576));
    Span4Mux_s3_h I__11666 (
            .O(N__51576),
            .I(N__51572));
    InMux I__11665 (
            .O(N__51575),
            .I(N__51569));
    Span4Mux_v I__11664 (
            .O(N__51572),
            .I(N__51566));
    LocalMux I__11663 (
            .O(N__51569),
            .I(N__51563));
    Odrv4 I__11662 (
            .O(N__51566),
            .I(\pid_side.error_5 ));
    Odrv12 I__11661 (
            .O(N__51563),
            .I(\pid_side.error_5 ));
    InMux I__11660 (
            .O(N__51558),
            .I(\pid_side.error_cry_0_0 ));
    InMux I__11659 (
            .O(N__51555),
            .I(N__51552));
    LocalMux I__11658 (
            .O(N__51552),
            .I(\pid_side.un1_pid_prereg_107_0 ));
    InMux I__11657 (
            .O(N__51549),
            .I(N__51545));
    InMux I__11656 (
            .O(N__51548),
            .I(N__51542));
    LocalMux I__11655 (
            .O(N__51545),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11 ));
    LocalMux I__11654 (
            .O(N__51542),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11 ));
    InMux I__11653 (
            .O(N__51537),
            .I(N__51528));
    InMux I__11652 (
            .O(N__51536),
            .I(N__51528));
    InMux I__11651 (
            .O(N__51535),
            .I(N__51528));
    LocalMux I__11650 (
            .O(N__51528),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    InMux I__11649 (
            .O(N__51525),
            .I(N__51520));
    InMux I__11648 (
            .O(N__51524),
            .I(N__51515));
    InMux I__11647 (
            .O(N__51523),
            .I(N__51515));
    LocalMux I__11646 (
            .O(N__51520),
            .I(N__51510));
    LocalMux I__11645 (
            .O(N__51515),
            .I(N__51510));
    Odrv12 I__11644 (
            .O(N__51510),
            .I(\pid_side.error_d_reg_prev_esr_RNI2VN9Z0Z_12 ));
    InMux I__11643 (
            .O(N__51507),
            .I(N__51503));
    InMux I__11642 (
            .O(N__51506),
            .I(N__51500));
    LocalMux I__11641 (
            .O(N__51503),
            .I(\pid_side.error_d_reg_prevZ0Z_11 ));
    LocalMux I__11640 (
            .O(N__51500),
            .I(\pid_side.error_d_reg_prevZ0Z_11 ));
    InMux I__11639 (
            .O(N__51495),
            .I(N__51492));
    LocalMux I__11638 (
            .O(N__51492),
            .I(N__51489));
    Span4Mux_h I__11637 (
            .O(N__51489),
            .I(N__51486));
    Odrv4 I__11636 (
            .O(N__51486),
            .I(\pid_side.O_2_15 ));
    InMux I__11635 (
            .O(N__51483),
            .I(N__51479));
    InMux I__11634 (
            .O(N__51482),
            .I(N__51476));
    LocalMux I__11633 (
            .O(N__51479),
            .I(N__51473));
    LocalMux I__11632 (
            .O(N__51476),
            .I(\pid_side.error_p_regZ0Z_11 ));
    Odrv4 I__11631 (
            .O(N__51473),
            .I(\pid_side.error_p_regZ0Z_11 ));
    InMux I__11630 (
            .O(N__51468),
            .I(N__51465));
    LocalMux I__11629 (
            .O(N__51465),
            .I(N__51462));
    Span12Mux_s9_h I__11628 (
            .O(N__51462),
            .I(N__51459));
    Odrv12 I__11627 (
            .O(N__51459),
            .I(\ppm_encoder_1.N_291 ));
    InMux I__11626 (
            .O(N__51456),
            .I(N__51453));
    LocalMux I__11625 (
            .O(N__51453),
            .I(N__51445));
    InMux I__11624 (
            .O(N__51452),
            .I(N__51442));
    InMux I__11623 (
            .O(N__51451),
            .I(N__51437));
    InMux I__11622 (
            .O(N__51450),
            .I(N__51437));
    CascadeMux I__11621 (
            .O(N__51449),
            .I(N__51433));
    CascadeMux I__11620 (
            .O(N__51448),
            .I(N__51428));
    Span4Mux_v I__11619 (
            .O(N__51445),
            .I(N__51419));
    LocalMux I__11618 (
            .O(N__51442),
            .I(N__51419));
    LocalMux I__11617 (
            .O(N__51437),
            .I(N__51419));
    InMux I__11616 (
            .O(N__51436),
            .I(N__51416));
    InMux I__11615 (
            .O(N__51433),
            .I(N__51412));
    CascadeMux I__11614 (
            .O(N__51432),
            .I(N__51406));
    InMux I__11613 (
            .O(N__51431),
            .I(N__51401));
    InMux I__11612 (
            .O(N__51428),
            .I(N__51397));
    InMux I__11611 (
            .O(N__51427),
            .I(N__51394));
    InMux I__11610 (
            .O(N__51426),
            .I(N__51391));
    Span4Mux_v I__11609 (
            .O(N__51419),
            .I(N__51386));
    LocalMux I__11608 (
            .O(N__51416),
            .I(N__51386));
    InMux I__11607 (
            .O(N__51415),
            .I(N__51383));
    LocalMux I__11606 (
            .O(N__51412),
            .I(N__51378));
    InMux I__11605 (
            .O(N__51411),
            .I(N__51375));
    InMux I__11604 (
            .O(N__51410),
            .I(N__51372));
    InMux I__11603 (
            .O(N__51409),
            .I(N__51369));
    InMux I__11602 (
            .O(N__51406),
            .I(N__51366));
    InMux I__11601 (
            .O(N__51405),
            .I(N__51362));
    InMux I__11600 (
            .O(N__51404),
            .I(N__51359));
    LocalMux I__11599 (
            .O(N__51401),
            .I(N__51356));
    CascadeMux I__11598 (
            .O(N__51400),
            .I(N__51353));
    LocalMux I__11597 (
            .O(N__51397),
            .I(N__51350));
    LocalMux I__11596 (
            .O(N__51394),
            .I(N__51347));
    LocalMux I__11595 (
            .O(N__51391),
            .I(N__51342));
    Span4Mux_v I__11594 (
            .O(N__51386),
            .I(N__51342));
    LocalMux I__11593 (
            .O(N__51383),
            .I(N__51339));
    InMux I__11592 (
            .O(N__51382),
            .I(N__51334));
    InMux I__11591 (
            .O(N__51381),
            .I(N__51334));
    Span4Mux_v I__11590 (
            .O(N__51378),
            .I(N__51329));
    LocalMux I__11589 (
            .O(N__51375),
            .I(N__51329));
    LocalMux I__11588 (
            .O(N__51372),
            .I(N__51324));
    LocalMux I__11587 (
            .O(N__51369),
            .I(N__51324));
    LocalMux I__11586 (
            .O(N__51366),
            .I(N__51321));
    InMux I__11585 (
            .O(N__51365),
            .I(N__51318));
    LocalMux I__11584 (
            .O(N__51362),
            .I(N__51315));
    LocalMux I__11583 (
            .O(N__51359),
            .I(N__51310));
    Span4Mux_h I__11582 (
            .O(N__51356),
            .I(N__51310));
    InMux I__11581 (
            .O(N__51353),
            .I(N__51307));
    Span4Mux_h I__11580 (
            .O(N__51350),
            .I(N__51298));
    Span4Mux_v I__11579 (
            .O(N__51347),
            .I(N__51298));
    Span4Mux_h I__11578 (
            .O(N__51342),
            .I(N__51298));
    Span4Mux_h I__11577 (
            .O(N__51339),
            .I(N__51298));
    LocalMux I__11576 (
            .O(N__51334),
            .I(N__51291));
    Span4Mux_v I__11575 (
            .O(N__51329),
            .I(N__51291));
    Span4Mux_v I__11574 (
            .O(N__51324),
            .I(N__51291));
    Span4Mux_v I__11573 (
            .O(N__51321),
            .I(N__51282));
    LocalMux I__11572 (
            .O(N__51318),
            .I(N__51282));
    Span4Mux_h I__11571 (
            .O(N__51315),
            .I(N__51282));
    Span4Mux_v I__11570 (
            .O(N__51310),
            .I(N__51282));
    LocalMux I__11569 (
            .O(N__51307),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__11568 (
            .O(N__51298),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__11567 (
            .O(N__51291),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__11566 (
            .O(N__51282),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    InMux I__11565 (
            .O(N__51273),
            .I(N__51270));
    LocalMux I__11564 (
            .O(N__51270),
            .I(N__51266));
    InMux I__11563 (
            .O(N__51269),
            .I(N__51262));
    Span4Mux_v I__11562 (
            .O(N__51266),
            .I(N__51259));
    InMux I__11561 (
            .O(N__51265),
            .I(N__51256));
    LocalMux I__11560 (
            .O(N__51262),
            .I(N__51249));
    Sp12to4 I__11559 (
            .O(N__51259),
            .I(N__51249));
    LocalMux I__11558 (
            .O(N__51256),
            .I(N__51249));
    Odrv12 I__11557 (
            .O(N__51249),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__11556 (
            .O(N__51246),
            .I(N__51243));
    LocalMux I__11555 (
            .O(N__51243),
            .I(N__51240));
    Span4Mux_h I__11554 (
            .O(N__51240),
            .I(N__51237));
    Span4Mux_h I__11553 (
            .O(N__51237),
            .I(N__51234));
    Span4Mux_v I__11552 (
            .O(N__51234),
            .I(N__51231));
    Odrv4 I__11551 (
            .O(N__51231),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ));
    CascadeMux I__11550 (
            .O(N__51228),
            .I(N__51223));
    InMux I__11549 (
            .O(N__51227),
            .I(N__51220));
    InMux I__11548 (
            .O(N__51226),
            .I(N__51215));
    InMux I__11547 (
            .O(N__51223),
            .I(N__51215));
    LocalMux I__11546 (
            .O(N__51220),
            .I(N__51210));
    LocalMux I__11545 (
            .O(N__51215),
            .I(N__51210));
    Span4Mux_v I__11544 (
            .O(N__51210),
            .I(N__51207));
    Odrv4 I__11543 (
            .O(N__51207),
            .I(\pid_side.un1_pid_prereg_56 ));
    CascadeMux I__11542 (
            .O(N__51204),
            .I(N__51201));
    InMux I__11541 (
            .O(N__51201),
            .I(N__51198));
    LocalMux I__11540 (
            .O(N__51198),
            .I(\pid_side.error_d_reg_prev_esr_RNIO9BH1Z0Z_20 ));
    InMux I__11539 (
            .O(N__51195),
            .I(N__51192));
    LocalMux I__11538 (
            .O(N__51192),
            .I(N__51189));
    Odrv4 I__11537 (
            .O(N__51189),
            .I(\pid_side.error_d_reg_prev_esr_RNILJFJ2Z0Z_12 ));
    CascadeMux I__11536 (
            .O(N__51186),
            .I(\pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10_cascade_ ));
    CascadeMux I__11535 (
            .O(N__51183),
            .I(N__51180));
    InMux I__11534 (
            .O(N__51180),
            .I(N__51176));
    InMux I__11533 (
            .O(N__51179),
            .I(N__51173));
    LocalMux I__11532 (
            .O(N__51176),
            .I(N__51170));
    LocalMux I__11531 (
            .O(N__51173),
            .I(\pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10 ));
    Odrv4 I__11530 (
            .O(N__51170),
            .I(\pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10 ));
    CascadeMux I__11529 (
            .O(N__51165),
            .I(N__51162));
    InMux I__11528 (
            .O(N__51162),
            .I(N__51159));
    LocalMux I__11527 (
            .O(N__51159),
            .I(N__51155));
    InMux I__11526 (
            .O(N__51158),
            .I(N__51152));
    Odrv4 I__11525 (
            .O(N__51155),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11 ));
    LocalMux I__11524 (
            .O(N__51152),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11 ));
    CascadeMux I__11523 (
            .O(N__51147),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11_cascade_ ));
    InMux I__11522 (
            .O(N__51144),
            .I(N__51138));
    InMux I__11521 (
            .O(N__51143),
            .I(N__51138));
    LocalMux I__11520 (
            .O(N__51138),
            .I(\pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10 ));
    CascadeMux I__11519 (
            .O(N__51135),
            .I(N__51132));
    InMux I__11518 (
            .O(N__51132),
            .I(N__51129));
    LocalMux I__11517 (
            .O(N__51129),
            .I(N__51126));
    Odrv4 I__11516 (
            .O(N__51126),
            .I(\pid_side.error_d_reg_prev_esr_RNIQCA21Z0Z_10 ));
    InMux I__11515 (
            .O(N__51123),
            .I(N__51119));
    CascadeMux I__11514 (
            .O(N__51122),
            .I(N__51116));
    LocalMux I__11513 (
            .O(N__51119),
            .I(N__51113));
    InMux I__11512 (
            .O(N__51116),
            .I(N__51110));
    Odrv12 I__11511 (
            .O(N__51113),
            .I(\pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12 ));
    LocalMux I__11510 (
            .O(N__51110),
            .I(\pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12 ));
    CascadeMux I__11509 (
            .O(N__51105),
            .I(\pid_side.N_1590_i_cascade_ ));
    InMux I__11508 (
            .O(N__51102),
            .I(N__51099));
    LocalMux I__11507 (
            .O(N__51099),
            .I(N__51096));
    Odrv4 I__11506 (
            .O(N__51096),
            .I(\pid_side.error_d_reg_esr_RNIVTFJ2Z0Z_12 ));
    InMux I__11505 (
            .O(N__51093),
            .I(N__51090));
    LocalMux I__11504 (
            .O(N__51090),
            .I(N__51087));
    Odrv4 I__11503 (
            .O(N__51087),
            .I(\pid_side.error_d_reg_prev_esr_RNI4NA21Z0Z_12 ));
    InMux I__11502 (
            .O(N__51084),
            .I(N__51081));
    LocalMux I__11501 (
            .O(N__51081),
            .I(\pid_side.error_d_reg_prev_esr_RNIDP5H1Z0Z_14 ));
    InMux I__11500 (
            .O(N__51078),
            .I(N__51075));
    LocalMux I__11499 (
            .O(N__51075),
            .I(\pid_side.error_d_reg_esr_RNIKMFP2Z0Z_10 ));
    InMux I__11498 (
            .O(N__51072),
            .I(N__51069));
    LocalMux I__11497 (
            .O(N__51069),
            .I(\pid_side.N_1582_i ));
    CascadeMux I__11496 (
            .O(N__51066),
            .I(\pid_side.N_1582_i_cascade_ ));
    InMux I__11495 (
            .O(N__51063),
            .I(N__51060));
    LocalMux I__11494 (
            .O(N__51060),
            .I(\pid_side.error_d_reg_esr_RNI104E2Z0Z_10 ));
    InMux I__11493 (
            .O(N__51057),
            .I(N__51054));
    LocalMux I__11492 (
            .O(N__51054),
            .I(N__51051));
    Odrv4 I__11491 (
            .O(N__51051),
            .I(\pid_side.error_d_reg_prev_esr_RNIKCB23Z0Z_13 ));
    InMux I__11490 (
            .O(N__51048),
            .I(N__51043));
    InMux I__11489 (
            .O(N__51047),
            .I(N__51038));
    InMux I__11488 (
            .O(N__51046),
            .I(N__51038));
    LocalMux I__11487 (
            .O(N__51043),
            .I(\pid_side.un1_pid_prereg_23 ));
    LocalMux I__11486 (
            .O(N__51038),
            .I(\pid_side.un1_pid_prereg_23 ));
    CascadeMux I__11485 (
            .O(N__51033),
            .I(N__51030));
    InMux I__11484 (
            .O(N__51030),
            .I(N__51027));
    LocalMux I__11483 (
            .O(N__51027),
            .I(N__51023));
    InMux I__11482 (
            .O(N__51026),
            .I(N__51020));
    Odrv12 I__11481 (
            .O(N__51023),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ));
    LocalMux I__11480 (
            .O(N__51020),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ));
    CascadeMux I__11479 (
            .O(N__51015),
            .I(N__51012));
    InMux I__11478 (
            .O(N__51012),
            .I(N__51006));
    InMux I__11477 (
            .O(N__51011),
            .I(N__51006));
    LocalMux I__11476 (
            .O(N__51006),
            .I(\pid_side.un1_pid_prereg_18 ));
    CascadeMux I__11475 (
            .O(N__51003),
            .I(N__51000));
    InMux I__11474 (
            .O(N__51000),
            .I(N__50997));
    LocalMux I__11473 (
            .O(N__50997),
            .I(\pid_side.error_d_reg_prev_esr_RNIBAGJ2Z0Z_12 ));
    InMux I__11472 (
            .O(N__50994),
            .I(N__50989));
    InMux I__11471 (
            .O(N__50993),
            .I(N__50984));
    InMux I__11470 (
            .O(N__50992),
            .I(N__50984));
    LocalMux I__11469 (
            .O(N__50989),
            .I(\pid_side.un1_pid_prereg_29 ));
    LocalMux I__11468 (
            .O(N__50984),
            .I(\pid_side.un1_pid_prereg_29 ));
    InMux I__11467 (
            .O(N__50979),
            .I(N__50973));
    InMux I__11466 (
            .O(N__50978),
            .I(N__50973));
    LocalMux I__11465 (
            .O(N__50973),
            .I(\pid_side.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__11464 (
            .O(N__50970),
            .I(\pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1_cascade_ ));
    CascadeMux I__11463 (
            .O(N__50967),
            .I(N__50963));
    InMux I__11462 (
            .O(N__50966),
            .I(N__50960));
    InMux I__11461 (
            .O(N__50963),
            .I(N__50957));
    LocalMux I__11460 (
            .O(N__50960),
            .I(\pid_side.un1_pid_prereg ));
    LocalMux I__11459 (
            .O(N__50957),
            .I(\pid_side.un1_pid_prereg ));
    InMux I__11458 (
            .O(N__50952),
            .I(N__50943));
    InMux I__11457 (
            .O(N__50951),
            .I(N__50943));
    InMux I__11456 (
            .O(N__50950),
            .I(N__50943));
    LocalMux I__11455 (
            .O(N__50943),
            .I(\pid_side.error_d_reg_prevZ0Z_0 ));
    InMux I__11454 (
            .O(N__50940),
            .I(N__50937));
    LocalMux I__11453 (
            .O(N__50937),
            .I(N__50933));
    InMux I__11452 (
            .O(N__50936),
            .I(N__50930));
    Odrv12 I__11451 (
            .O(N__50933),
            .I(\pid_side.un1_pid_prereg_axb_0 ));
    LocalMux I__11450 (
            .O(N__50930),
            .I(\pid_side.un1_pid_prereg_axb_0 ));
    InMux I__11449 (
            .O(N__50925),
            .I(N__50922));
    LocalMux I__11448 (
            .O(N__50922),
            .I(\pid_side.error_p_reg_esr_RNIAVKD1Z0Z_1 ));
    CascadeMux I__11447 (
            .O(N__50919),
            .I(\pid_side.un1_pid_prereg_18_cascade_ ));
    CascadeMux I__11446 (
            .O(N__50916),
            .I(N__50913));
    InMux I__11445 (
            .O(N__50913),
            .I(N__50910));
    LocalMux I__11444 (
            .O(N__50910),
            .I(N__50907));
    Odrv4 I__11443 (
            .O(N__50907),
            .I(\pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13 ));
    CascadeMux I__11442 (
            .O(N__50904),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13_cascade_ ));
    InMux I__11441 (
            .O(N__50901),
            .I(N__50895));
    InMux I__11440 (
            .O(N__50900),
            .I(N__50895));
    LocalMux I__11439 (
            .O(N__50895),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    CascadeMux I__11438 (
            .O(N__50892),
            .I(N__50889));
    InMux I__11437 (
            .O(N__50889),
            .I(N__50883));
    InMux I__11436 (
            .O(N__50888),
            .I(N__50883));
    LocalMux I__11435 (
            .O(N__50883),
            .I(N__50880));
    Odrv4 I__11434 (
            .O(N__50880),
            .I(side_command_7));
    InMux I__11433 (
            .O(N__50877),
            .I(N__50874));
    LocalMux I__11432 (
            .O(N__50874),
            .I(N__50871));
    Odrv12 I__11431 (
            .O(N__50871),
            .I(\pid_front.O_7 ));
    InMux I__11430 (
            .O(N__50868),
            .I(N__50859));
    InMux I__11429 (
            .O(N__50867),
            .I(N__50859));
    InMux I__11428 (
            .O(N__50866),
            .I(N__50859));
    LocalMux I__11427 (
            .O(N__50859),
            .I(N__50856));
    Span4Mux_h I__11426 (
            .O(N__50856),
            .I(N__50853));
    Span4Mux_h I__11425 (
            .O(N__50853),
            .I(N__50850));
    Odrv4 I__11424 (
            .O(N__50850),
            .I(\pid_front.error_d_regZ0Z_3 ));
    CascadeMux I__11423 (
            .O(N__50847),
            .I(N__50844));
    InMux I__11422 (
            .O(N__50844),
            .I(N__50841));
    LocalMux I__11421 (
            .O(N__50841),
            .I(N__50838));
    Span4Mux_h I__11420 (
            .O(N__50838),
            .I(N__50835));
    Odrv4 I__11419 (
            .O(N__50835),
            .I(\pid_side.error_p_reg_esr_RNI5QI23Z0Z_5 ));
    InMux I__11418 (
            .O(N__50832),
            .I(N__50829));
    LocalMux I__11417 (
            .O(N__50829),
            .I(N__50825));
    InMux I__11416 (
            .O(N__50828),
            .I(N__50822));
    Odrv12 I__11415 (
            .O(N__50825),
            .I(\pid_side.un1_pid_prereg_axb_1 ));
    LocalMux I__11414 (
            .O(N__50822),
            .I(\pid_side.un1_pid_prereg_axb_1 ));
    CascadeMux I__11413 (
            .O(N__50817),
            .I(\pid_side.error_p_reg_esr_RNISH6JZ0Z_0_cascade_ ));
    InMux I__11412 (
            .O(N__50814),
            .I(N__50811));
    LocalMux I__11411 (
            .O(N__50811),
            .I(\pid_side.error_d_reg_esr_RNIFP9R2Z0Z_1 ));
    InMux I__11410 (
            .O(N__50808),
            .I(N__50802));
    InMux I__11409 (
            .O(N__50807),
            .I(N__50802));
    LocalMux I__11408 (
            .O(N__50802),
            .I(\pid_side.N_1546_i ));
    InMux I__11407 (
            .O(N__50799),
            .I(N__50796));
    LocalMux I__11406 (
            .O(N__50796),
            .I(N__50793));
    Span4Mux_h I__11405 (
            .O(N__50793),
            .I(N__50790));
    Span4Mux_h I__11404 (
            .O(N__50790),
            .I(N__50787));
    Span4Mux_v I__11403 (
            .O(N__50787),
            .I(N__50784));
    Odrv4 I__11402 (
            .O(N__50784),
            .I(drone_H_disp_front_i_9));
    InMux I__11401 (
            .O(N__50781),
            .I(N__50776));
    InMux I__11400 (
            .O(N__50780),
            .I(N__50773));
    InMux I__11399 (
            .O(N__50779),
            .I(N__50769));
    LocalMux I__11398 (
            .O(N__50776),
            .I(N__50762));
    LocalMux I__11397 (
            .O(N__50773),
            .I(N__50762));
    InMux I__11396 (
            .O(N__50772),
            .I(N__50759));
    LocalMux I__11395 (
            .O(N__50769),
            .I(N__50756));
    InMux I__11394 (
            .O(N__50768),
            .I(N__50753));
    InMux I__11393 (
            .O(N__50767),
            .I(N__50750));
    Span4Mux_v I__11392 (
            .O(N__50762),
            .I(N__50746));
    LocalMux I__11391 (
            .O(N__50759),
            .I(N__50743));
    Span4Mux_h I__11390 (
            .O(N__50756),
            .I(N__50738));
    LocalMux I__11389 (
            .O(N__50753),
            .I(N__50738));
    LocalMux I__11388 (
            .O(N__50750),
            .I(N__50735));
    InMux I__11387 (
            .O(N__50749),
            .I(N__50732));
    Sp12to4 I__11386 (
            .O(N__50746),
            .I(N__50728));
    Span4Mux_h I__11385 (
            .O(N__50743),
            .I(N__50725));
    Span4Mux_v I__11384 (
            .O(N__50738),
            .I(N__50718));
    Span4Mux_h I__11383 (
            .O(N__50735),
            .I(N__50718));
    LocalMux I__11382 (
            .O(N__50732),
            .I(N__50718));
    InMux I__11381 (
            .O(N__50731),
            .I(N__50715));
    Span12Mux_h I__11380 (
            .O(N__50728),
            .I(N__50706));
    Sp12to4 I__11379 (
            .O(N__50725),
            .I(N__50706));
    Sp12to4 I__11378 (
            .O(N__50718),
            .I(N__50706));
    LocalMux I__11377 (
            .O(N__50715),
            .I(N__50706));
    Odrv12 I__11376 (
            .O(N__50706),
            .I(uart_drone_data_1));
    InMux I__11375 (
            .O(N__50703),
            .I(N__50700));
    LocalMux I__11374 (
            .O(N__50700),
            .I(\dron_frame_decoder_1.drone_H_disp_front_9 ));
    CEMux I__11373 (
            .O(N__50697),
            .I(N__50693));
    CEMux I__11372 (
            .O(N__50696),
            .I(N__50689));
    LocalMux I__11371 (
            .O(N__50693),
            .I(N__50686));
    CEMux I__11370 (
            .O(N__50692),
            .I(N__50683));
    LocalMux I__11369 (
            .O(N__50689),
            .I(N__50680));
    Span4Mux_h I__11368 (
            .O(N__50686),
            .I(N__50677));
    LocalMux I__11367 (
            .O(N__50683),
            .I(N__50674));
    Sp12to4 I__11366 (
            .O(N__50680),
            .I(N__50671));
    Sp12to4 I__11365 (
            .O(N__50677),
            .I(N__50668));
    Span4Mux_h I__11364 (
            .O(N__50674),
            .I(N__50665));
    Span12Mux_v I__11363 (
            .O(N__50671),
            .I(N__50662));
    Span12Mux_v I__11362 (
            .O(N__50668),
            .I(N__50659));
    Sp12to4 I__11361 (
            .O(N__50665),
            .I(N__50656));
    Odrv12 I__11360 (
            .O(N__50662),
            .I(\dron_frame_decoder_1.N_481_0 ));
    Odrv12 I__11359 (
            .O(N__50659),
            .I(\dron_frame_decoder_1.N_481_0 ));
    Odrv12 I__11358 (
            .O(N__50656),
            .I(\dron_frame_decoder_1.N_481_0 ));
    InMux I__11357 (
            .O(N__50649),
            .I(N__50646));
    LocalMux I__11356 (
            .O(N__50646),
            .I(\dron_frame_decoder_1.drone_H_disp_side_4 ));
    InMux I__11355 (
            .O(N__50643),
            .I(N__50640));
    LocalMux I__11354 (
            .O(N__50640),
            .I(N__50637));
    Odrv4 I__11353 (
            .O(N__50637),
            .I(\dron_frame_decoder_1.drone_H_disp_side_6 ));
    InMux I__11352 (
            .O(N__50634),
            .I(N__50631));
    LocalMux I__11351 (
            .O(N__50631),
            .I(N__50628));
    Odrv4 I__11350 (
            .O(N__50628),
            .I(\dron_frame_decoder_1.drone_H_disp_side_7 ));
    InMux I__11349 (
            .O(N__50625),
            .I(N__50619));
    InMux I__11348 (
            .O(N__50624),
            .I(N__50612));
    InMux I__11347 (
            .O(N__50623),
            .I(N__50612));
    InMux I__11346 (
            .O(N__50622),
            .I(N__50612));
    LocalMux I__11345 (
            .O(N__50619),
            .I(N__50602));
    LocalMux I__11344 (
            .O(N__50612),
            .I(N__50599));
    InMux I__11343 (
            .O(N__50611),
            .I(N__50596));
    InMux I__11342 (
            .O(N__50610),
            .I(N__50583));
    InMux I__11341 (
            .O(N__50609),
            .I(N__50583));
    InMux I__11340 (
            .O(N__50608),
            .I(N__50583));
    InMux I__11339 (
            .O(N__50607),
            .I(N__50583));
    InMux I__11338 (
            .O(N__50606),
            .I(N__50583));
    InMux I__11337 (
            .O(N__50605),
            .I(N__50583));
    Span4Mux_h I__11336 (
            .O(N__50602),
            .I(N__50580));
    Span4Mux_h I__11335 (
            .O(N__50599),
            .I(N__50577));
    LocalMux I__11334 (
            .O(N__50596),
            .I(N__50574));
    LocalMux I__11333 (
            .O(N__50583),
            .I(N__50571));
    Span4Mux_h I__11332 (
            .O(N__50580),
            .I(N__50568));
    Span4Mux_h I__11331 (
            .O(N__50577),
            .I(N__50565));
    Span12Mux_h I__11330 (
            .O(N__50574),
            .I(N__50562));
    Span12Mux_h I__11329 (
            .O(N__50571),
            .I(N__50559));
    Span4Mux_v I__11328 (
            .O(N__50568),
            .I(N__50556));
    Span4Mux_h I__11327 (
            .O(N__50565),
            .I(N__50553));
    Odrv12 I__11326 (
            .O(N__50562),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv12 I__11325 (
            .O(N__50559),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__11324 (
            .O(N__50556),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__11323 (
            .O(N__50553),
            .I(\pid_front.stateZ0Z_1 ));
    InMux I__11322 (
            .O(N__50544),
            .I(N__50541));
    LocalMux I__11321 (
            .O(N__50541),
            .I(N__50538));
    Span4Mux_h I__11320 (
            .O(N__50538),
            .I(N__50535));
    Span4Mux_h I__11319 (
            .O(N__50535),
            .I(N__50532));
    Odrv4 I__11318 (
            .O(N__50532),
            .I(\pid_front.un1_pid_prereg_cry_0_THRU_CO ));
    InMux I__11317 (
            .O(N__50529),
            .I(N__50526));
    LocalMux I__11316 (
            .O(N__50526),
            .I(N__50523));
    Span4Mux_v I__11315 (
            .O(N__50523),
            .I(N__50520));
    Span4Mux_h I__11314 (
            .O(N__50520),
            .I(N__50516));
    InMux I__11313 (
            .O(N__50519),
            .I(N__50513));
    Odrv4 I__11312 (
            .O(N__50516),
            .I(\pid_front.un1_pid_prereg_axb_1 ));
    LocalMux I__11311 (
            .O(N__50513),
            .I(\pid_front.un1_pid_prereg_axb_1 ));
    InMux I__11310 (
            .O(N__50508),
            .I(N__50502));
    CascadeMux I__11309 (
            .O(N__50507),
            .I(N__50499));
    InMux I__11308 (
            .O(N__50506),
            .I(N__50494));
    InMux I__11307 (
            .O(N__50505),
            .I(N__50494));
    LocalMux I__11306 (
            .O(N__50502),
            .I(N__50490));
    InMux I__11305 (
            .O(N__50499),
            .I(N__50487));
    LocalMux I__11304 (
            .O(N__50494),
            .I(N__50484));
    InMux I__11303 (
            .O(N__50493),
            .I(N__50481));
    Span4Mux_v I__11302 (
            .O(N__50490),
            .I(N__50477));
    LocalMux I__11301 (
            .O(N__50487),
            .I(N__50474));
    Span12Mux_v I__11300 (
            .O(N__50484),
            .I(N__50471));
    LocalMux I__11299 (
            .O(N__50481),
            .I(N__50468));
    InMux I__11298 (
            .O(N__50480),
            .I(N__50465));
    Span4Mux_h I__11297 (
            .O(N__50477),
            .I(N__50462));
    Span4Mux_v I__11296 (
            .O(N__50474),
            .I(N__50459));
    Span12Mux_h I__11295 (
            .O(N__50471),
            .I(N__50454));
    Span12Mux_s4_v I__11294 (
            .O(N__50468),
            .I(N__50454));
    LocalMux I__11293 (
            .O(N__50465),
            .I(N__50447));
    Span4Mux_h I__11292 (
            .O(N__50462),
            .I(N__50447));
    Span4Mux_v I__11291 (
            .O(N__50459),
            .I(N__50447));
    Odrv12 I__11290 (
            .O(N__50454),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv4 I__11289 (
            .O(N__50447),
            .I(\pid_front.stateZ0Z_0 ));
    InMux I__11288 (
            .O(N__50442),
            .I(N__50438));
    InMux I__11287 (
            .O(N__50441),
            .I(N__50435));
    LocalMux I__11286 (
            .O(N__50438),
            .I(N__50431));
    LocalMux I__11285 (
            .O(N__50435),
            .I(N__50428));
    CascadeMux I__11284 (
            .O(N__50434),
            .I(N__50425));
    Span4Mux_v I__11283 (
            .O(N__50431),
            .I(N__50420));
    Span4Mux_v I__11282 (
            .O(N__50428),
            .I(N__50420));
    InMux I__11281 (
            .O(N__50425),
            .I(N__50417));
    Sp12to4 I__11280 (
            .O(N__50420),
            .I(N__50414));
    LocalMux I__11279 (
            .O(N__50417),
            .I(\pid_front.pid_preregZ0Z_1 ));
    Odrv12 I__11278 (
            .O(N__50414),
            .I(\pid_front.pid_preregZ0Z_1 ));
    InMux I__11277 (
            .O(N__50409),
            .I(N__50406));
    LocalMux I__11276 (
            .O(N__50406),
            .I(drone_H_disp_side_1));
    InMux I__11275 (
            .O(N__50403),
            .I(N__50399));
    InMux I__11274 (
            .O(N__50402),
            .I(N__50395));
    LocalMux I__11273 (
            .O(N__50399),
            .I(N__50391));
    InMux I__11272 (
            .O(N__50398),
            .I(N__50388));
    LocalMux I__11271 (
            .O(N__50395),
            .I(N__50385));
    InMux I__11270 (
            .O(N__50394),
            .I(N__50380));
    Span4Mux_v I__11269 (
            .O(N__50391),
            .I(N__50375));
    LocalMux I__11268 (
            .O(N__50388),
            .I(N__50375));
    Span4Mux_h I__11267 (
            .O(N__50385),
            .I(N__50372));
    InMux I__11266 (
            .O(N__50384),
            .I(N__50369));
    InMux I__11265 (
            .O(N__50383),
            .I(N__50366));
    LocalMux I__11264 (
            .O(N__50380),
            .I(N__50363));
    Span4Mux_v I__11263 (
            .O(N__50375),
            .I(N__50360));
    Span4Mux_h I__11262 (
            .O(N__50372),
            .I(N__50357));
    LocalMux I__11261 (
            .O(N__50369),
            .I(N__50354));
    LocalMux I__11260 (
            .O(N__50366),
            .I(N__50351));
    Span12Mux_s4_h I__11259 (
            .O(N__50363),
            .I(N__50348));
    Span4Mux_v I__11258 (
            .O(N__50360),
            .I(N__50345));
    Span4Mux_h I__11257 (
            .O(N__50357),
            .I(N__50340));
    Span4Mux_v I__11256 (
            .O(N__50354),
            .I(N__50340));
    Span4Mux_v I__11255 (
            .O(N__50351),
            .I(N__50337));
    Span12Mux_v I__11254 (
            .O(N__50348),
            .I(N__50333));
    Span4Mux_v I__11253 (
            .O(N__50345),
            .I(N__50330));
    Span4Mux_v I__11252 (
            .O(N__50340),
            .I(N__50327));
    Span4Mux_v I__11251 (
            .O(N__50337),
            .I(N__50324));
    InMux I__11250 (
            .O(N__50336),
            .I(N__50321));
    Odrv12 I__11249 (
            .O(N__50333),
            .I(uart_drone_data_2));
    Odrv4 I__11248 (
            .O(N__50330),
            .I(uart_drone_data_2));
    Odrv4 I__11247 (
            .O(N__50327),
            .I(uart_drone_data_2));
    Odrv4 I__11246 (
            .O(N__50324),
            .I(uart_drone_data_2));
    LocalMux I__11245 (
            .O(N__50321),
            .I(uart_drone_data_2));
    InMux I__11244 (
            .O(N__50310),
            .I(N__50307));
    LocalMux I__11243 (
            .O(N__50307),
            .I(drone_H_disp_side_2));
    InMux I__11242 (
            .O(N__50304),
            .I(N__50301));
    LocalMux I__11241 (
            .O(N__50301),
            .I(drone_H_disp_side_3));
    CEMux I__11240 (
            .O(N__50298),
            .I(N__50294));
    CEMux I__11239 (
            .O(N__50297),
            .I(N__50291));
    LocalMux I__11238 (
            .O(N__50294),
            .I(N__50288));
    LocalMux I__11237 (
            .O(N__50291),
            .I(N__50285));
    Span4Mux_h I__11236 (
            .O(N__50288),
            .I(N__50280));
    Span4Mux_v I__11235 (
            .O(N__50285),
            .I(N__50280));
    Sp12to4 I__11234 (
            .O(N__50280),
            .I(N__50277));
    Odrv12 I__11233 (
            .O(N__50277),
            .I(\dron_frame_decoder_1.N_505_0 ));
    InMux I__11232 (
            .O(N__50274),
            .I(N__50271));
    LocalMux I__11231 (
            .O(N__50271),
            .I(N__50268));
    Odrv12 I__11230 (
            .O(N__50268),
            .I(\pid_side.error_d_reg_prev_esr_RNIGJM23Z0Z_20 ));
    InMux I__11229 (
            .O(N__50265),
            .I(N__50262));
    LocalMux I__11228 (
            .O(N__50262),
            .I(N__50259));
    Odrv12 I__11227 (
            .O(N__50259),
            .I(\pid_side.un1_pid_prereg_axb_21 ));
    InMux I__11226 (
            .O(N__50256),
            .I(N__50253));
    LocalMux I__11225 (
            .O(N__50253),
            .I(N__50250));
    Span4Mux_v I__11224 (
            .O(N__50250),
            .I(N__50247));
    Odrv4 I__11223 (
            .O(N__50247),
            .I(\ppm_encoder_1.N_286 ));
    InMux I__11222 (
            .O(N__50244),
            .I(N__50241));
    LocalMux I__11221 (
            .O(N__50241),
            .I(N__50237));
    InMux I__11220 (
            .O(N__50240),
            .I(N__50234));
    Span4Mux_v I__11219 (
            .O(N__50237),
            .I(N__50230));
    LocalMux I__11218 (
            .O(N__50234),
            .I(N__50227));
    InMux I__11217 (
            .O(N__50233),
            .I(N__50224));
    Span4Mux_h I__11216 (
            .O(N__50230),
            .I(N__50219));
    Span4Mux_v I__11215 (
            .O(N__50227),
            .I(N__50219));
    LocalMux I__11214 (
            .O(N__50224),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    Odrv4 I__11213 (
            .O(N__50219),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    InMux I__11212 (
            .O(N__50214),
            .I(N__50211));
    LocalMux I__11211 (
            .O(N__50211),
            .I(N__50208));
    Span4Mux_h I__11210 (
            .O(N__50208),
            .I(N__50205));
    Span4Mux_v I__11209 (
            .O(N__50205),
            .I(N__50202));
    Span4Mux_v I__11208 (
            .O(N__50202),
            .I(N__50199));
    Odrv4 I__11207 (
            .O(N__50199),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ));
    CascadeMux I__11206 (
            .O(N__50196),
            .I(N__50193));
    InMux I__11205 (
            .O(N__50193),
            .I(N__50190));
    LocalMux I__11204 (
            .O(N__50190),
            .I(N__50187));
    Odrv12 I__11203 (
            .O(N__50187),
            .I(\pid_side.error_d_reg_prev_esr_RNIGV8H1Z0Z_19 ));
    CascadeMux I__11202 (
            .O(N__50184),
            .I(\pid_side.un1_pid_prereg_30_cascade_ ));
    CascadeMux I__11201 (
            .O(N__50181),
            .I(N__50178));
    InMux I__11200 (
            .O(N__50178),
            .I(N__50175));
    LocalMux I__11199 (
            .O(N__50175),
            .I(\pid_side.error_d_reg_prev_esr_RNI0PB23Z0Z_14 ));
    InMux I__11198 (
            .O(N__50172),
            .I(N__50169));
    LocalMux I__11197 (
            .O(N__50169),
            .I(\pid_side.error_d_reg_prev_esr_RNI4UC23Z0Z_17 ));
    CascadeMux I__11196 (
            .O(N__50166),
            .I(N__50163));
    InMux I__11195 (
            .O(N__50163),
            .I(N__50160));
    LocalMux I__11194 (
            .O(N__50160),
            .I(\pid_side.error_d_reg_prev_esr_RNI5I6H1Z0Z_18 ));
    InMux I__11193 (
            .O(N__50157),
            .I(N__50154));
    LocalMux I__11192 (
            .O(N__50154),
            .I(N__50151));
    Odrv4 I__11191 (
            .O(N__50151),
            .I(\pid_side.error_d_reg_prev_esr_RNIP56H1Z0Z_16 ));
    CascadeMux I__11190 (
            .O(N__50148),
            .I(N__50145));
    InMux I__11189 (
            .O(N__50145),
            .I(N__50139));
    InMux I__11188 (
            .O(N__50144),
            .I(N__50139));
    LocalMux I__11187 (
            .O(N__50139),
            .I(\pid_side.error_d_reg_prevZ0Z_16 ));
    InMux I__11186 (
            .O(N__50136),
            .I(N__50131));
    InMux I__11185 (
            .O(N__50135),
            .I(N__50126));
    InMux I__11184 (
            .O(N__50134),
            .I(N__50126));
    LocalMux I__11183 (
            .O(N__50131),
            .I(\pid_side.un1_pid_prereg_35 ));
    LocalMux I__11182 (
            .O(N__50126),
            .I(\pid_side.un1_pid_prereg_35 ));
    CascadeMux I__11181 (
            .O(N__50121),
            .I(\pid_side.un1_pid_prereg_36_cascade_ ));
    InMux I__11180 (
            .O(N__50118),
            .I(N__50114));
    InMux I__11179 (
            .O(N__50117),
            .I(N__50111));
    LocalMux I__11178 (
            .O(N__50114),
            .I(\pid_side.un1_pid_prereg_30 ));
    LocalMux I__11177 (
            .O(N__50111),
            .I(\pid_side.un1_pid_prereg_30 ));
    CascadeMux I__11176 (
            .O(N__50106),
            .I(N__50103));
    InMux I__11175 (
            .O(N__50103),
            .I(N__50100));
    LocalMux I__11174 (
            .O(N__50100),
            .I(N__50097));
    Odrv4 I__11173 (
            .O(N__50097),
            .I(\pid_side.error_d_reg_prev_esr_RNIC5C23Z0Z_15 ));
    InMux I__11172 (
            .O(N__50094),
            .I(N__50091));
    LocalMux I__11171 (
            .O(N__50091),
            .I(N__50088));
    Odrv4 I__11170 (
            .O(N__50088),
            .I(\pid_side.error_d_reg_prev_esr_RNI89K23Z0Z_19 ));
    InMux I__11169 (
            .O(N__50085),
            .I(N__50082));
    LocalMux I__11168 (
            .O(N__50082),
            .I(N__50079));
    Span4Mux_h I__11167 (
            .O(N__50079),
            .I(N__50076));
    Odrv4 I__11166 (
            .O(N__50076),
            .I(\pid_side.pid_preregZ0Z_19 ));
    InMux I__11165 (
            .O(N__50073),
            .I(\pid_side.un1_pid_prereg_cry_16 ));
    InMux I__11164 (
            .O(N__50070),
            .I(N__50067));
    LocalMux I__11163 (
            .O(N__50067),
            .I(N__50064));
    Odrv4 I__11162 (
            .O(N__50064),
            .I(\pid_side.pid_preregZ0Z_20 ));
    InMux I__11161 (
            .O(N__50061),
            .I(\pid_side.un1_pid_prereg_cry_17 ));
    InMux I__11160 (
            .O(N__50058),
            .I(N__50055));
    LocalMux I__11159 (
            .O(N__50055),
            .I(N__50052));
    Odrv4 I__11158 (
            .O(N__50052),
            .I(\pid_side.pid_preregZ0Z_21 ));
    InMux I__11157 (
            .O(N__50049),
            .I(\pid_side.un1_pid_prereg_cry_18 ));
    InMux I__11156 (
            .O(N__50046),
            .I(N__50043));
    LocalMux I__11155 (
            .O(N__50043),
            .I(N__50040));
    Span4Mux_h I__11154 (
            .O(N__50040),
            .I(N__50037));
    Odrv4 I__11153 (
            .O(N__50037),
            .I(\pid_side.pid_preregZ0Z_22 ));
    InMux I__11152 (
            .O(N__50034),
            .I(\pid_side.un1_pid_prereg_cry_19 ));
    InMux I__11151 (
            .O(N__50031),
            .I(\pid_side.un1_pid_prereg_cry_20 ));
    CascadeMux I__11150 (
            .O(N__50028),
            .I(N__50025));
    InMux I__11149 (
            .O(N__50025),
            .I(N__50021));
    InMux I__11148 (
            .O(N__50024),
            .I(N__50017));
    LocalMux I__11147 (
            .O(N__50021),
            .I(N__50011));
    InMux I__11146 (
            .O(N__50020),
            .I(N__50008));
    LocalMux I__11145 (
            .O(N__50017),
            .I(N__50005));
    InMux I__11144 (
            .O(N__50016),
            .I(N__49998));
    InMux I__11143 (
            .O(N__50015),
            .I(N__49998));
    InMux I__11142 (
            .O(N__50014),
            .I(N__49998));
    Span4Mux_v I__11141 (
            .O(N__50011),
            .I(N__49993));
    LocalMux I__11140 (
            .O(N__50008),
            .I(N__49993));
    Span4Mux_h I__11139 (
            .O(N__50005),
            .I(N__49990));
    LocalMux I__11138 (
            .O(N__49998),
            .I(N__49987));
    Odrv4 I__11137 (
            .O(N__49993),
            .I(\pid_side.pid_preregZ0Z_23 ));
    Odrv4 I__11136 (
            .O(N__49990),
            .I(\pid_side.pid_preregZ0Z_23 ));
    Odrv12 I__11135 (
            .O(N__49987),
            .I(\pid_side.pid_preregZ0Z_23 ));
    InMux I__11134 (
            .O(N__49980),
            .I(N__49977));
    LocalMux I__11133 (
            .O(N__49977),
            .I(\pid_side.error_d_reg_prev_esr_RNILHF23Z0Z_18 ));
    InMux I__11132 (
            .O(N__49974),
            .I(N__49971));
    LocalMux I__11131 (
            .O(N__49971),
            .I(\pid_side.error_d_reg_prev_esr_RNIJV5H1Z0Z_15 ));
    InMux I__11130 (
            .O(N__49968),
            .I(N__49962));
    InMux I__11129 (
            .O(N__49967),
            .I(N__49959));
    InMux I__11128 (
            .O(N__49966),
            .I(N__49956));
    InMux I__11127 (
            .O(N__49965),
            .I(N__49953));
    LocalMux I__11126 (
            .O(N__49962),
            .I(N__49950));
    LocalMux I__11125 (
            .O(N__49959),
            .I(N__49947));
    LocalMux I__11124 (
            .O(N__49956),
            .I(N__49942));
    LocalMux I__11123 (
            .O(N__49953),
            .I(N__49942));
    Span4Mux_h I__11122 (
            .O(N__49950),
            .I(N__49939));
    Odrv12 I__11121 (
            .O(N__49947),
            .I(\pid_side.pid_preregZ0Z_10 ));
    Odrv4 I__11120 (
            .O(N__49942),
            .I(\pid_side.pid_preregZ0Z_10 ));
    Odrv4 I__11119 (
            .O(N__49939),
            .I(\pid_side.pid_preregZ0Z_10 ));
    InMux I__11118 (
            .O(N__49932),
            .I(\pid_side.un1_pid_prereg_cry_7 ));
    InMux I__11117 (
            .O(N__49929),
            .I(N__49923));
    InMux I__11116 (
            .O(N__49928),
            .I(N__49920));
    InMux I__11115 (
            .O(N__49927),
            .I(N__49917));
    InMux I__11114 (
            .O(N__49926),
            .I(N__49914));
    LocalMux I__11113 (
            .O(N__49923),
            .I(N__49911));
    LocalMux I__11112 (
            .O(N__49920),
            .I(N__49904));
    LocalMux I__11111 (
            .O(N__49917),
            .I(N__49904));
    LocalMux I__11110 (
            .O(N__49914),
            .I(N__49904));
    Span4Mux_h I__11109 (
            .O(N__49911),
            .I(N__49901));
    Odrv12 I__11108 (
            .O(N__49904),
            .I(\pid_side.pid_preregZ0Z_11 ));
    Odrv4 I__11107 (
            .O(N__49901),
            .I(\pid_side.pid_preregZ0Z_11 ));
    InMux I__11106 (
            .O(N__49896),
            .I(\pid_side.un1_pid_prereg_cry_8 ));
    CascadeMux I__11105 (
            .O(N__49893),
            .I(N__49889));
    InMux I__11104 (
            .O(N__49892),
            .I(N__49886));
    InMux I__11103 (
            .O(N__49889),
            .I(N__49883));
    LocalMux I__11102 (
            .O(N__49886),
            .I(N__49876));
    LocalMux I__11101 (
            .O(N__49883),
            .I(N__49876));
    InMux I__11100 (
            .O(N__49882),
            .I(N__49871));
    InMux I__11099 (
            .O(N__49881),
            .I(N__49871));
    Span4Mux_v I__11098 (
            .O(N__49876),
            .I(N__49868));
    LocalMux I__11097 (
            .O(N__49871),
            .I(N__49865));
    Odrv4 I__11096 (
            .O(N__49868),
            .I(\pid_side.pid_preregZ0Z_12 ));
    Odrv4 I__11095 (
            .O(N__49865),
            .I(\pid_side.pid_preregZ0Z_12 ));
    InMux I__11094 (
            .O(N__49860),
            .I(\pid_side.un1_pid_prereg_cry_9 ));
    InMux I__11093 (
            .O(N__49857),
            .I(N__49851));
    InMux I__11092 (
            .O(N__49856),
            .I(N__49848));
    InMux I__11091 (
            .O(N__49855),
            .I(N__49843));
    InMux I__11090 (
            .O(N__49854),
            .I(N__49843));
    LocalMux I__11089 (
            .O(N__49851),
            .I(N__49835));
    LocalMux I__11088 (
            .O(N__49848),
            .I(N__49835));
    LocalMux I__11087 (
            .O(N__49843),
            .I(N__49835));
    InMux I__11086 (
            .O(N__49842),
            .I(N__49832));
    Span4Mux_v I__11085 (
            .O(N__49835),
            .I(N__49827));
    LocalMux I__11084 (
            .O(N__49832),
            .I(N__49827));
    Odrv4 I__11083 (
            .O(N__49827),
            .I(\pid_side.pid_preregZ0Z_13 ));
    InMux I__11082 (
            .O(N__49824),
            .I(\pid_side.un1_pid_prereg_cry_10 ));
    InMux I__11081 (
            .O(N__49821),
            .I(N__49818));
    LocalMux I__11080 (
            .O(N__49818),
            .I(N__49815));
    Span4Mux_h I__11079 (
            .O(N__49815),
            .I(N__49812));
    Odrv4 I__11078 (
            .O(N__49812),
            .I(\pid_side.pid_preregZ0Z_14 ));
    InMux I__11077 (
            .O(N__49809),
            .I(\pid_side.un1_pid_prereg_cry_11 ));
    InMux I__11076 (
            .O(N__49806),
            .I(N__49803));
    LocalMux I__11075 (
            .O(N__49803),
            .I(N__49800));
    Odrv4 I__11074 (
            .O(N__49800),
            .I(\pid_side.pid_preregZ0Z_15 ));
    InMux I__11073 (
            .O(N__49797),
            .I(\pid_side.un1_pid_prereg_cry_12 ));
    InMux I__11072 (
            .O(N__49794),
            .I(N__49791));
    LocalMux I__11071 (
            .O(N__49791),
            .I(N__49788));
    Odrv4 I__11070 (
            .O(N__49788),
            .I(\pid_side.pid_preregZ0Z_16 ));
    InMux I__11069 (
            .O(N__49785),
            .I(bfn_20_11_0_));
    InMux I__11068 (
            .O(N__49782),
            .I(N__49779));
    LocalMux I__11067 (
            .O(N__49779),
            .I(N__49776));
    Odrv4 I__11066 (
            .O(N__49776),
            .I(\pid_side.pid_preregZ0Z_17 ));
    InMux I__11065 (
            .O(N__49773),
            .I(\pid_side.un1_pid_prereg_cry_14 ));
    CascadeMux I__11064 (
            .O(N__49770),
            .I(N__49767));
    InMux I__11063 (
            .O(N__49767),
            .I(N__49764));
    LocalMux I__11062 (
            .O(N__49764),
            .I(N__49761));
    Odrv4 I__11061 (
            .O(N__49761),
            .I(\pid_side.pid_preregZ0Z_18 ));
    InMux I__11060 (
            .O(N__49758),
            .I(\pid_side.un1_pid_prereg_cry_15 ));
    InMux I__11059 (
            .O(N__49755),
            .I(N__49752));
    LocalMux I__11058 (
            .O(N__49752),
            .I(N__49749));
    Span4Mux_v I__11057 (
            .O(N__49749),
            .I(N__49745));
    InMux I__11056 (
            .O(N__49748),
            .I(N__49742));
    Span4Mux_h I__11055 (
            .O(N__49745),
            .I(N__49739));
    LocalMux I__11054 (
            .O(N__49742),
            .I(N__49736));
    Odrv4 I__11053 (
            .O(N__49739),
            .I(\pid_side.pid_preregZ0Z_2 ));
    Odrv4 I__11052 (
            .O(N__49736),
            .I(\pid_side.pid_preregZ0Z_2 ));
    InMux I__11051 (
            .O(N__49731),
            .I(\pid_side.un1_pid_prereg_cry_1 ));
    InMux I__11050 (
            .O(N__49728),
            .I(N__49725));
    LocalMux I__11049 (
            .O(N__49725),
            .I(N__49721));
    CascadeMux I__11048 (
            .O(N__49724),
            .I(N__49718));
    Span4Mux_v I__11047 (
            .O(N__49721),
            .I(N__49715));
    InMux I__11046 (
            .O(N__49718),
            .I(N__49712));
    Span4Mux_h I__11045 (
            .O(N__49715),
            .I(N__49709));
    LocalMux I__11044 (
            .O(N__49712),
            .I(N__49706));
    Odrv4 I__11043 (
            .O(N__49709),
            .I(\pid_side.pid_preregZ0Z_3 ));
    Odrv4 I__11042 (
            .O(N__49706),
            .I(\pid_side.pid_preregZ0Z_3 ));
    InMux I__11041 (
            .O(N__49701),
            .I(\pid_side.un1_pid_prereg_cry_0_0 ));
    InMux I__11040 (
            .O(N__49698),
            .I(N__49691));
    CascadeMux I__11039 (
            .O(N__49697),
            .I(N__49688));
    CascadeMux I__11038 (
            .O(N__49696),
            .I(N__49685));
    CascadeMux I__11037 (
            .O(N__49695),
            .I(N__49682));
    CascadeMux I__11036 (
            .O(N__49694),
            .I(N__49678));
    LocalMux I__11035 (
            .O(N__49691),
            .I(N__49675));
    InMux I__11034 (
            .O(N__49688),
            .I(N__49672));
    InMux I__11033 (
            .O(N__49685),
            .I(N__49665));
    InMux I__11032 (
            .O(N__49682),
            .I(N__49665));
    InMux I__11031 (
            .O(N__49681),
            .I(N__49665));
    InMux I__11030 (
            .O(N__49678),
            .I(N__49661));
    Span4Mux_h I__11029 (
            .O(N__49675),
            .I(N__49656));
    LocalMux I__11028 (
            .O(N__49672),
            .I(N__49656));
    LocalMux I__11027 (
            .O(N__49665),
            .I(N__49653));
    InMux I__11026 (
            .O(N__49664),
            .I(N__49650));
    LocalMux I__11025 (
            .O(N__49661),
            .I(N__49647));
    Span4Mux_v I__11024 (
            .O(N__49656),
            .I(N__49642));
    Span4Mux_v I__11023 (
            .O(N__49653),
            .I(N__49642));
    LocalMux I__11022 (
            .O(N__49650),
            .I(N__49639));
    Span4Mux_v I__11021 (
            .O(N__49647),
            .I(N__49636));
    Span4Mux_h I__11020 (
            .O(N__49642),
            .I(N__49633));
    Span4Mux_v I__11019 (
            .O(N__49639),
            .I(N__49628));
    Span4Mux_h I__11018 (
            .O(N__49636),
            .I(N__49628));
    Odrv4 I__11017 (
            .O(N__49633),
            .I(\pid_side.pid_preregZ0Z_4 ));
    Odrv4 I__11016 (
            .O(N__49628),
            .I(\pid_side.pid_preregZ0Z_4 ));
    InMux I__11015 (
            .O(N__49623),
            .I(\pid_side.un1_pid_prereg_cry_1_0 ));
    CascadeMux I__11014 (
            .O(N__49620),
            .I(N__49615));
    CascadeMux I__11013 (
            .O(N__49619),
            .I(N__49612));
    CascadeMux I__11012 (
            .O(N__49618),
            .I(N__49608));
    InMux I__11011 (
            .O(N__49615),
            .I(N__49605));
    InMux I__11010 (
            .O(N__49612),
            .I(N__49602));
    InMux I__11009 (
            .O(N__49611),
            .I(N__49599));
    InMux I__11008 (
            .O(N__49608),
            .I(N__49596));
    LocalMux I__11007 (
            .O(N__49605),
            .I(N__49593));
    LocalMux I__11006 (
            .O(N__49602),
            .I(N__49590));
    LocalMux I__11005 (
            .O(N__49599),
            .I(N__49585));
    LocalMux I__11004 (
            .O(N__49596),
            .I(N__49585));
    Span4Mux_v I__11003 (
            .O(N__49593),
            .I(N__49580));
    Span4Mux_v I__11002 (
            .O(N__49590),
            .I(N__49580));
    Span4Mux_v I__11001 (
            .O(N__49585),
            .I(N__49577));
    Odrv4 I__11000 (
            .O(N__49580),
            .I(\pid_side.pid_preregZ0Z_5 ));
    Odrv4 I__10999 (
            .O(N__49577),
            .I(\pid_side.pid_preregZ0Z_5 ));
    InMux I__10998 (
            .O(N__49572),
            .I(\pid_side.un1_pid_prereg_cry_2 ));
    CascadeMux I__10997 (
            .O(N__49569),
            .I(N__49565));
    InMux I__10996 (
            .O(N__49568),
            .I(N__49561));
    InMux I__10995 (
            .O(N__49565),
            .I(N__49556));
    InMux I__10994 (
            .O(N__49564),
            .I(N__49556));
    LocalMux I__10993 (
            .O(N__49561),
            .I(N__49551));
    LocalMux I__10992 (
            .O(N__49556),
            .I(N__49551));
    Span4Mux_h I__10991 (
            .O(N__49551),
            .I(N__49548));
    Odrv4 I__10990 (
            .O(N__49548),
            .I(\pid_side.pid_preregZ0Z_6 ));
    InMux I__10989 (
            .O(N__49545),
            .I(\pid_side.un1_pid_prereg_cry_3 ));
    InMux I__10988 (
            .O(N__49542),
            .I(N__49538));
    CascadeMux I__10987 (
            .O(N__49541),
            .I(N__49534));
    LocalMux I__10986 (
            .O(N__49538),
            .I(N__49531));
    InMux I__10985 (
            .O(N__49537),
            .I(N__49528));
    InMux I__10984 (
            .O(N__49534),
            .I(N__49525));
    Span4Mux_h I__10983 (
            .O(N__49531),
            .I(N__49518));
    LocalMux I__10982 (
            .O(N__49528),
            .I(N__49518));
    LocalMux I__10981 (
            .O(N__49525),
            .I(N__49518));
    Span4Mux_h I__10980 (
            .O(N__49518),
            .I(N__49515));
    Odrv4 I__10979 (
            .O(N__49515),
            .I(\pid_side.pid_preregZ0Z_7 ));
    InMux I__10978 (
            .O(N__49512),
            .I(\pid_side.un1_pid_prereg_cry_4 ));
    InMux I__10977 (
            .O(N__49509),
            .I(N__49504));
    InMux I__10976 (
            .O(N__49508),
            .I(N__49499));
    InMux I__10975 (
            .O(N__49507),
            .I(N__49499));
    LocalMux I__10974 (
            .O(N__49504),
            .I(N__49494));
    LocalMux I__10973 (
            .O(N__49499),
            .I(N__49494));
    Odrv12 I__10972 (
            .O(N__49494),
            .I(\pid_side.pid_preregZ0Z_8 ));
    InMux I__10971 (
            .O(N__49491),
            .I(bfn_20_10_0_));
    InMux I__10970 (
            .O(N__49488),
            .I(N__49483));
    InMux I__10969 (
            .O(N__49487),
            .I(N__49480));
    InMux I__10968 (
            .O(N__49486),
            .I(N__49477));
    LocalMux I__10967 (
            .O(N__49483),
            .I(N__49470));
    LocalMux I__10966 (
            .O(N__49480),
            .I(N__49470));
    LocalMux I__10965 (
            .O(N__49477),
            .I(N__49470));
    Span4Mux_h I__10964 (
            .O(N__49470),
            .I(N__49467));
    Odrv4 I__10963 (
            .O(N__49467),
            .I(\pid_side.pid_preregZ0Z_9 ));
    InMux I__10962 (
            .O(N__49464),
            .I(\pid_side.un1_pid_prereg_cry_6 ));
    InMux I__10961 (
            .O(N__49461),
            .I(N__49457));
    InMux I__10960 (
            .O(N__49460),
            .I(N__49454));
    LocalMux I__10959 (
            .O(N__49457),
            .I(N__49451));
    LocalMux I__10958 (
            .O(N__49454),
            .I(N__49448));
    Span4Mux_v I__10957 (
            .O(N__49451),
            .I(N__49445));
    Span4Mux_v I__10956 (
            .O(N__49448),
            .I(N__49442));
    Sp12to4 I__10955 (
            .O(N__49445),
            .I(N__49439));
    Span4Mux_h I__10954 (
            .O(N__49442),
            .I(N__49436));
    Odrv12 I__10953 (
            .O(N__49439),
            .I(\pid_front.un1_pid_prereg_axb_0 ));
    Odrv4 I__10952 (
            .O(N__49436),
            .I(\pid_front.un1_pid_prereg_axb_0 ));
    InMux I__10951 (
            .O(N__49431),
            .I(N__49428));
    LocalMux I__10950 (
            .O(N__49428),
            .I(N__49424));
    InMux I__10949 (
            .O(N__49427),
            .I(N__49420));
    Span4Mux_h I__10948 (
            .O(N__49424),
            .I(N__49417));
    InMux I__10947 (
            .O(N__49423),
            .I(N__49414));
    LocalMux I__10946 (
            .O(N__49420),
            .I(N__49411));
    Odrv4 I__10945 (
            .O(N__49417),
            .I(\pid_front.pid_preregZ0Z_0 ));
    LocalMux I__10944 (
            .O(N__49414),
            .I(\pid_front.pid_preregZ0Z_0 ));
    Odrv12 I__10943 (
            .O(N__49411),
            .I(\pid_front.pid_preregZ0Z_0 ));
    CascadeMux I__10942 (
            .O(N__49404),
            .I(N__49401));
    InMux I__10941 (
            .O(N__49401),
            .I(N__49397));
    InMux I__10940 (
            .O(N__49400),
            .I(N__49394));
    LocalMux I__10939 (
            .O(N__49397),
            .I(N__49389));
    LocalMux I__10938 (
            .O(N__49394),
            .I(N__49389));
    Span4Mux_v I__10937 (
            .O(N__49389),
            .I(N__49386));
    Span4Mux_h I__10936 (
            .O(N__49386),
            .I(N__49383));
    Span4Mux_h I__10935 (
            .O(N__49383),
            .I(N__49380));
    Odrv4 I__10934 (
            .O(N__49380),
            .I(\pid_front.error_d_reg_prevZ0Z_18 ));
    CEMux I__10933 (
            .O(N__49377),
            .I(N__49317));
    CEMux I__10932 (
            .O(N__49376),
            .I(N__49317));
    CEMux I__10931 (
            .O(N__49375),
            .I(N__49317));
    CEMux I__10930 (
            .O(N__49374),
            .I(N__49317));
    CEMux I__10929 (
            .O(N__49373),
            .I(N__49317));
    CEMux I__10928 (
            .O(N__49372),
            .I(N__49317));
    CEMux I__10927 (
            .O(N__49371),
            .I(N__49317));
    CEMux I__10926 (
            .O(N__49370),
            .I(N__49317));
    CEMux I__10925 (
            .O(N__49369),
            .I(N__49317));
    CEMux I__10924 (
            .O(N__49368),
            .I(N__49317));
    CEMux I__10923 (
            .O(N__49367),
            .I(N__49317));
    CEMux I__10922 (
            .O(N__49366),
            .I(N__49317));
    CEMux I__10921 (
            .O(N__49365),
            .I(N__49317));
    CEMux I__10920 (
            .O(N__49364),
            .I(N__49317));
    CEMux I__10919 (
            .O(N__49363),
            .I(N__49317));
    CEMux I__10918 (
            .O(N__49362),
            .I(N__49317));
    CEMux I__10917 (
            .O(N__49361),
            .I(N__49317));
    CEMux I__10916 (
            .O(N__49360),
            .I(N__49317));
    CEMux I__10915 (
            .O(N__49359),
            .I(N__49317));
    CEMux I__10914 (
            .O(N__49358),
            .I(N__49317));
    GlobalMux I__10913 (
            .O(N__49317),
            .I(N__49314));
    gio2CtrlBuf I__10912 (
            .O(N__49314),
            .I(\pid_front.state_0_g_0 ));
    InMux I__10911 (
            .O(N__49311),
            .I(N__49308));
    LocalMux I__10910 (
            .O(N__49308),
            .I(N__49305));
    Odrv12 I__10909 (
            .O(N__49305),
            .I(\pid_front.O_6 ));
    InMux I__10908 (
            .O(N__49302),
            .I(N__49296));
    InMux I__10907 (
            .O(N__49301),
            .I(N__49296));
    LocalMux I__10906 (
            .O(N__49296),
            .I(N__49292));
    InMux I__10905 (
            .O(N__49295),
            .I(N__49289));
    Span4Mux_h I__10904 (
            .O(N__49292),
            .I(N__49286));
    LocalMux I__10903 (
            .O(N__49289),
            .I(N__49283));
    Span4Mux_h I__10902 (
            .O(N__49286),
            .I(N__49280));
    Span12Mux_v I__10901 (
            .O(N__49283),
            .I(N__49277));
    Odrv4 I__10900 (
            .O(N__49280),
            .I(\pid_front.error_d_regZ0Z_2 ));
    Odrv12 I__10899 (
            .O(N__49277),
            .I(\pid_front.error_d_regZ0Z_2 ));
    IoInMux I__10898 (
            .O(N__49272),
            .I(N__49269));
    LocalMux I__10897 (
            .O(N__49269),
            .I(GB_BUFFER_reset_system_g_THRU_CO));
    InMux I__10896 (
            .O(N__49266),
            .I(N__49263));
    LocalMux I__10895 (
            .O(N__49263),
            .I(N__49260));
    Odrv4 I__10894 (
            .O(N__49260),
            .I(\pid_side.un1_pid_prereg_cry_0_THRU_CO ));
    InMux I__10893 (
            .O(N__49257),
            .I(\pid_side.un1_pid_prereg_cry_0 ));
    InMux I__10892 (
            .O(N__49254),
            .I(N__49251));
    LocalMux I__10891 (
            .O(N__49251),
            .I(N__49248));
    Odrv4 I__10890 (
            .O(N__49248),
            .I(\ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ));
    CascadeMux I__10889 (
            .O(N__49245),
            .I(N__49242));
    InMux I__10888 (
            .O(N__49242),
            .I(N__49239));
    LocalMux I__10887 (
            .O(N__49239),
            .I(N__49236));
    Odrv4 I__10886 (
            .O(N__49236),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ));
    InMux I__10885 (
            .O(N__49233),
            .I(N__49230));
    LocalMux I__10884 (
            .O(N__49230),
            .I(N__49227));
    Span4Mux_h I__10883 (
            .O(N__49227),
            .I(N__49224));
    Odrv4 I__10882 (
            .O(N__49224),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__10881 (
            .O(N__49221),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__10880 (
            .O(N__49218),
            .I(N__49215));
    LocalMux I__10879 (
            .O(N__49215),
            .I(N__49212));
    Span4Mux_h I__10878 (
            .O(N__49212),
            .I(N__49209));
    Odrv4 I__10877 (
            .O(N__49209),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__10876 (
            .O(N__49206),
            .I(N__49203));
    LocalMux I__10875 (
            .O(N__49203),
            .I(N__49200));
    Span4Mux_v I__10874 (
            .O(N__49200),
            .I(N__49197));
    Odrv4 I__10873 (
            .O(N__49197),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__10872 (
            .O(N__49194),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__10871 (
            .O(N__49191),
            .I(N__49188));
    LocalMux I__10870 (
            .O(N__49188),
            .I(N__49185));
    Odrv12 I__10869 (
            .O(N__49185),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__10868 (
            .O(N__49182),
            .I(N__49179));
    LocalMux I__10867 (
            .O(N__49179),
            .I(N__49176));
    Span4Mux_v I__10866 (
            .O(N__49176),
            .I(N__49173));
    Odrv4 I__10865 (
            .O(N__49173),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__10864 (
            .O(N__49170),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__10863 (
            .O(N__49167),
            .I(N__49164));
    LocalMux I__10862 (
            .O(N__49164),
            .I(N__49161));
    Span4Mux_h I__10861 (
            .O(N__49161),
            .I(N__49158));
    Odrv4 I__10860 (
            .O(N__49158),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__10859 (
            .O(N__49155),
            .I(N__49152));
    LocalMux I__10858 (
            .O(N__49152),
            .I(N__49149));
    Span4Mux_v I__10857 (
            .O(N__49149),
            .I(N__49146));
    Odrv4 I__10856 (
            .O(N__49146),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__10855 (
            .O(N__49143),
            .I(bfn_18_17_0_));
    InMux I__10854 (
            .O(N__49140),
            .I(N__49137));
    LocalMux I__10853 (
            .O(N__49137),
            .I(N__49134));
    Span4Mux_h I__10852 (
            .O(N__49134),
            .I(N__49131));
    Odrv4 I__10851 (
            .O(N__49131),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    InMux I__10850 (
            .O(N__49128),
            .I(N__49125));
    LocalMux I__10849 (
            .O(N__49125),
            .I(N__49122));
    Span4Mux_h I__10848 (
            .O(N__49122),
            .I(N__49119));
    Odrv4 I__10847 (
            .O(N__49119),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__10846 (
            .O(N__49116),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__10845 (
            .O(N__49113),
            .I(N__49109));
    InMux I__10844 (
            .O(N__49112),
            .I(N__49106));
    LocalMux I__10843 (
            .O(N__49109),
            .I(N__49102));
    LocalMux I__10842 (
            .O(N__49106),
            .I(N__49099));
    CascadeMux I__10841 (
            .O(N__49105),
            .I(N__49096));
    Span4Mux_v I__10840 (
            .O(N__49102),
            .I(N__49091));
    Span4Mux_h I__10839 (
            .O(N__49099),
            .I(N__49091));
    InMux I__10838 (
            .O(N__49096),
            .I(N__49088));
    Odrv4 I__10837 (
            .O(N__49091),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__10836 (
            .O(N__49088),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    InMux I__10835 (
            .O(N__49083),
            .I(N__49070));
    CascadeMux I__10834 (
            .O(N__49082),
            .I(N__49062));
    InMux I__10833 (
            .O(N__49081),
            .I(N__49053));
    InMux I__10832 (
            .O(N__49080),
            .I(N__49053));
    InMux I__10831 (
            .O(N__49079),
            .I(N__49053));
    InMux I__10830 (
            .O(N__49078),
            .I(N__49044));
    InMux I__10829 (
            .O(N__49077),
            .I(N__49044));
    InMux I__10828 (
            .O(N__49076),
            .I(N__49044));
    InMux I__10827 (
            .O(N__49075),
            .I(N__49044));
    InMux I__10826 (
            .O(N__49074),
            .I(N__49040));
    InMux I__10825 (
            .O(N__49073),
            .I(N__49037));
    LocalMux I__10824 (
            .O(N__49070),
            .I(N__49034));
    InMux I__10823 (
            .O(N__49069),
            .I(N__49027));
    InMux I__10822 (
            .O(N__49068),
            .I(N__49027));
    InMux I__10821 (
            .O(N__49067),
            .I(N__49027));
    CascadeMux I__10820 (
            .O(N__49066),
            .I(N__49018));
    CascadeMux I__10819 (
            .O(N__49065),
            .I(N__49015));
    InMux I__10818 (
            .O(N__49062),
            .I(N__49008));
    InMux I__10817 (
            .O(N__49061),
            .I(N__49008));
    InMux I__10816 (
            .O(N__49060),
            .I(N__49005));
    LocalMux I__10815 (
            .O(N__49053),
            .I(N__49000));
    LocalMux I__10814 (
            .O(N__49044),
            .I(N__49000));
    CascadeMux I__10813 (
            .O(N__49043),
            .I(N__48991));
    LocalMux I__10812 (
            .O(N__49040),
            .I(N__48977));
    LocalMux I__10811 (
            .O(N__49037),
            .I(N__48977));
    Span4Mux_v I__10810 (
            .O(N__49034),
            .I(N__48977));
    LocalMux I__10809 (
            .O(N__49027),
            .I(N__48977));
    InMux I__10808 (
            .O(N__49026),
            .I(N__48972));
    InMux I__10807 (
            .O(N__49025),
            .I(N__48972));
    InMux I__10806 (
            .O(N__49024),
            .I(N__48967));
    InMux I__10805 (
            .O(N__49023),
            .I(N__48967));
    InMux I__10804 (
            .O(N__49022),
            .I(N__48956));
    InMux I__10803 (
            .O(N__49021),
            .I(N__48956));
    InMux I__10802 (
            .O(N__49018),
            .I(N__48956));
    InMux I__10801 (
            .O(N__49015),
            .I(N__48956));
    InMux I__10800 (
            .O(N__49014),
            .I(N__48956));
    InMux I__10799 (
            .O(N__49013),
            .I(N__48953));
    LocalMux I__10798 (
            .O(N__49008),
            .I(N__48950));
    LocalMux I__10797 (
            .O(N__49005),
            .I(N__48945));
    Span4Mux_h I__10796 (
            .O(N__49000),
            .I(N__48945));
    InMux I__10795 (
            .O(N__48999),
            .I(N__48936));
    InMux I__10794 (
            .O(N__48998),
            .I(N__48936));
    InMux I__10793 (
            .O(N__48997),
            .I(N__48936));
    InMux I__10792 (
            .O(N__48996),
            .I(N__48936));
    CascadeMux I__10791 (
            .O(N__48995),
            .I(N__48932));
    InMux I__10790 (
            .O(N__48994),
            .I(N__48928));
    InMux I__10789 (
            .O(N__48991),
            .I(N__48923));
    InMux I__10788 (
            .O(N__48990),
            .I(N__48923));
    InMux I__10787 (
            .O(N__48989),
            .I(N__48914));
    InMux I__10786 (
            .O(N__48988),
            .I(N__48914));
    InMux I__10785 (
            .O(N__48987),
            .I(N__48914));
    InMux I__10784 (
            .O(N__48986),
            .I(N__48914));
    Span4Mux_v I__10783 (
            .O(N__48977),
            .I(N__48909));
    LocalMux I__10782 (
            .O(N__48972),
            .I(N__48909));
    LocalMux I__10781 (
            .O(N__48967),
            .I(N__48904));
    LocalMux I__10780 (
            .O(N__48956),
            .I(N__48904));
    LocalMux I__10779 (
            .O(N__48953),
            .I(N__48895));
    Span4Mux_v I__10778 (
            .O(N__48950),
            .I(N__48895));
    Span4Mux_v I__10777 (
            .O(N__48945),
            .I(N__48895));
    LocalMux I__10776 (
            .O(N__48936),
            .I(N__48895));
    InMux I__10775 (
            .O(N__48935),
            .I(N__48888));
    InMux I__10774 (
            .O(N__48932),
            .I(N__48888));
    InMux I__10773 (
            .O(N__48931),
            .I(N__48888));
    LocalMux I__10772 (
            .O(N__48928),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10771 (
            .O(N__48923),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10770 (
            .O(N__48914),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__10769 (
            .O(N__48909),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__10768 (
            .O(N__48904),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__10767 (
            .O(N__48895),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10766 (
            .O(N__48888),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    InMux I__10765 (
            .O(N__48873),
            .I(N__48858));
    CascadeMux I__10764 (
            .O(N__48872),
            .I(N__48855));
    InMux I__10763 (
            .O(N__48871),
            .I(N__48848));
    InMux I__10762 (
            .O(N__48870),
            .I(N__48841));
    InMux I__10761 (
            .O(N__48869),
            .I(N__48841));
    InMux I__10760 (
            .O(N__48868),
            .I(N__48841));
    CascadeMux I__10759 (
            .O(N__48867),
            .I(N__48838));
    CascadeMux I__10758 (
            .O(N__48866),
            .I(N__48835));
    CascadeMux I__10757 (
            .O(N__48865),
            .I(N__48829));
    CascadeMux I__10756 (
            .O(N__48864),
            .I(N__48826));
    CascadeMux I__10755 (
            .O(N__48863),
            .I(N__48816));
    CascadeMux I__10754 (
            .O(N__48862),
            .I(N__48812));
    CascadeMux I__10753 (
            .O(N__48861),
            .I(N__48809));
    LocalMux I__10752 (
            .O(N__48858),
            .I(N__48805));
    InMux I__10751 (
            .O(N__48855),
            .I(N__48802));
    InMux I__10750 (
            .O(N__48854),
            .I(N__48799));
    InMux I__10749 (
            .O(N__48853),
            .I(N__48786));
    InMux I__10748 (
            .O(N__48852),
            .I(N__48781));
    InMux I__10747 (
            .O(N__48851),
            .I(N__48781));
    LocalMux I__10746 (
            .O(N__48848),
            .I(N__48776));
    LocalMux I__10745 (
            .O(N__48841),
            .I(N__48776));
    InMux I__10744 (
            .O(N__48838),
            .I(N__48769));
    InMux I__10743 (
            .O(N__48835),
            .I(N__48769));
    InMux I__10742 (
            .O(N__48834),
            .I(N__48769));
    InMux I__10741 (
            .O(N__48833),
            .I(N__48764));
    InMux I__10740 (
            .O(N__48832),
            .I(N__48764));
    InMux I__10739 (
            .O(N__48829),
            .I(N__48759));
    InMux I__10738 (
            .O(N__48826),
            .I(N__48759));
    InMux I__10737 (
            .O(N__48825),
            .I(N__48744));
    InMux I__10736 (
            .O(N__48824),
            .I(N__48744));
    InMux I__10735 (
            .O(N__48823),
            .I(N__48744));
    InMux I__10734 (
            .O(N__48822),
            .I(N__48744));
    InMux I__10733 (
            .O(N__48821),
            .I(N__48744));
    InMux I__10732 (
            .O(N__48820),
            .I(N__48744));
    InMux I__10731 (
            .O(N__48819),
            .I(N__48744));
    InMux I__10730 (
            .O(N__48816),
            .I(N__48730));
    InMux I__10729 (
            .O(N__48815),
            .I(N__48730));
    InMux I__10728 (
            .O(N__48812),
            .I(N__48723));
    InMux I__10727 (
            .O(N__48809),
            .I(N__48723));
    InMux I__10726 (
            .O(N__48808),
            .I(N__48723));
    Span4Mux_v I__10725 (
            .O(N__48805),
            .I(N__48718));
    LocalMux I__10724 (
            .O(N__48802),
            .I(N__48718));
    LocalMux I__10723 (
            .O(N__48799),
            .I(N__48715));
    InMux I__10722 (
            .O(N__48798),
            .I(N__48710));
    InMux I__10721 (
            .O(N__48797),
            .I(N__48710));
    CascadeMux I__10720 (
            .O(N__48796),
            .I(N__48706));
    CascadeMux I__10719 (
            .O(N__48795),
            .I(N__48703));
    InMux I__10718 (
            .O(N__48794),
            .I(N__48687));
    InMux I__10717 (
            .O(N__48793),
            .I(N__48687));
    InMux I__10716 (
            .O(N__48792),
            .I(N__48687));
    InMux I__10715 (
            .O(N__48791),
            .I(N__48687));
    InMux I__10714 (
            .O(N__48790),
            .I(N__48682));
    InMux I__10713 (
            .O(N__48789),
            .I(N__48682));
    LocalMux I__10712 (
            .O(N__48786),
            .I(N__48671));
    LocalMux I__10711 (
            .O(N__48781),
            .I(N__48671));
    Span4Mux_v I__10710 (
            .O(N__48776),
            .I(N__48671));
    LocalMux I__10709 (
            .O(N__48769),
            .I(N__48671));
    LocalMux I__10708 (
            .O(N__48764),
            .I(N__48671));
    LocalMux I__10707 (
            .O(N__48759),
            .I(N__48666));
    LocalMux I__10706 (
            .O(N__48744),
            .I(N__48666));
    InMux I__10705 (
            .O(N__48743),
            .I(N__48663));
    InMux I__10704 (
            .O(N__48742),
            .I(N__48654));
    InMux I__10703 (
            .O(N__48741),
            .I(N__48654));
    InMux I__10702 (
            .O(N__48740),
            .I(N__48654));
    InMux I__10701 (
            .O(N__48739),
            .I(N__48654));
    InMux I__10700 (
            .O(N__48738),
            .I(N__48647));
    InMux I__10699 (
            .O(N__48737),
            .I(N__48647));
    InMux I__10698 (
            .O(N__48736),
            .I(N__48647));
    CascadeMux I__10697 (
            .O(N__48735),
            .I(N__48632));
    LocalMux I__10696 (
            .O(N__48730),
            .I(N__48627));
    LocalMux I__10695 (
            .O(N__48723),
            .I(N__48627));
    Span4Mux_v I__10694 (
            .O(N__48718),
            .I(N__48622));
    Span4Mux_v I__10693 (
            .O(N__48715),
            .I(N__48622));
    LocalMux I__10692 (
            .O(N__48710),
            .I(N__48619));
    InMux I__10691 (
            .O(N__48709),
            .I(N__48610));
    InMux I__10690 (
            .O(N__48706),
            .I(N__48610));
    InMux I__10689 (
            .O(N__48703),
            .I(N__48610));
    InMux I__10688 (
            .O(N__48702),
            .I(N__48610));
    InMux I__10687 (
            .O(N__48701),
            .I(N__48599));
    InMux I__10686 (
            .O(N__48700),
            .I(N__48599));
    InMux I__10685 (
            .O(N__48699),
            .I(N__48599));
    InMux I__10684 (
            .O(N__48698),
            .I(N__48599));
    InMux I__10683 (
            .O(N__48697),
            .I(N__48599));
    InMux I__10682 (
            .O(N__48696),
            .I(N__48596));
    LocalMux I__10681 (
            .O(N__48687),
            .I(N__48587));
    LocalMux I__10680 (
            .O(N__48682),
            .I(N__48587));
    Span4Mux_v I__10679 (
            .O(N__48671),
            .I(N__48587));
    Span4Mux_h I__10678 (
            .O(N__48666),
            .I(N__48587));
    LocalMux I__10677 (
            .O(N__48663),
            .I(N__48580));
    LocalMux I__10676 (
            .O(N__48654),
            .I(N__48580));
    LocalMux I__10675 (
            .O(N__48647),
            .I(N__48580));
    InMux I__10674 (
            .O(N__48646),
            .I(N__48571));
    InMux I__10673 (
            .O(N__48645),
            .I(N__48571));
    InMux I__10672 (
            .O(N__48644),
            .I(N__48571));
    InMux I__10671 (
            .O(N__48643),
            .I(N__48571));
    InMux I__10670 (
            .O(N__48642),
            .I(N__48568));
    InMux I__10669 (
            .O(N__48641),
            .I(N__48557));
    InMux I__10668 (
            .O(N__48640),
            .I(N__48557));
    InMux I__10667 (
            .O(N__48639),
            .I(N__48557));
    InMux I__10666 (
            .O(N__48638),
            .I(N__48557));
    InMux I__10665 (
            .O(N__48637),
            .I(N__48557));
    InMux I__10664 (
            .O(N__48636),
            .I(N__48554));
    InMux I__10663 (
            .O(N__48635),
            .I(N__48549));
    InMux I__10662 (
            .O(N__48632),
            .I(N__48549));
    Odrv4 I__10661 (
            .O(N__48627),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10660 (
            .O(N__48622),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10659 (
            .O(N__48619),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10658 (
            .O(N__48610),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10657 (
            .O(N__48599),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10656 (
            .O(N__48596),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10655 (
            .O(N__48587),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10654 (
            .O(N__48580),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10653 (
            .O(N__48571),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10652 (
            .O(N__48568),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10651 (
            .O(N__48557),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10650 (
            .O(N__48554),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10649 (
            .O(N__48549),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    InMux I__10648 (
            .O(N__48522),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__10647 (
            .O(N__48519),
            .I(N__48516));
    LocalMux I__10646 (
            .O(N__48516),
            .I(N__48513));
    Span4Mux_v I__10645 (
            .O(N__48513),
            .I(N__48510));
    Odrv4 I__10644 (
            .O(N__48510),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__10643 (
            .O(N__48507),
            .I(N__48504));
    LocalMux I__10642 (
            .O(N__48504),
            .I(\dron_frame_decoder_1.drone_H_disp_side_5 ));
    InMux I__10641 (
            .O(N__48501),
            .I(N__48498));
    LocalMux I__10640 (
            .O(N__48498),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__10639 (
            .O(N__48495),
            .I(N__48492));
    LocalMux I__10638 (
            .O(N__48492),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__10637 (
            .O(N__48489),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__10636 (
            .O(N__48486),
            .I(N__48483));
    LocalMux I__10635 (
            .O(N__48483),
            .I(\ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ));
    CascadeMux I__10634 (
            .O(N__48480),
            .I(N__48477));
    InMux I__10633 (
            .O(N__48477),
            .I(N__48474));
    LocalMux I__10632 (
            .O(N__48474),
            .I(N__48471));
    Span4Mux_h I__10631 (
            .O(N__48471),
            .I(N__48468));
    Odrv4 I__10630 (
            .O(N__48468),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ));
    InMux I__10629 (
            .O(N__48465),
            .I(N__48462));
    LocalMux I__10628 (
            .O(N__48462),
            .I(N__48459));
    Span4Mux_h I__10627 (
            .O(N__48459),
            .I(N__48456));
    Odrv4 I__10626 (
            .O(N__48456),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__10625 (
            .O(N__48453),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    CascadeMux I__10624 (
            .O(N__48450),
            .I(N__48447));
    InMux I__10623 (
            .O(N__48447),
            .I(N__48444));
    LocalMux I__10622 (
            .O(N__48444),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__10621 (
            .O(N__48441),
            .I(N__48438));
    LocalMux I__10620 (
            .O(N__48438),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__10619 (
            .O(N__48435),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__10618 (
            .O(N__48432),
            .I(N__48429));
    LocalMux I__10617 (
            .O(N__48429),
            .I(N__48426));
    Odrv4 I__10616 (
            .O(N__48426),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__10615 (
            .O(N__48423),
            .I(N__48420));
    LocalMux I__10614 (
            .O(N__48420),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__10613 (
            .O(N__48417),
            .I(bfn_18_16_0_));
    InMux I__10612 (
            .O(N__48414),
            .I(N__48411));
    LocalMux I__10611 (
            .O(N__48411),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    InMux I__10610 (
            .O(N__48408),
            .I(N__48405));
    LocalMux I__10609 (
            .O(N__48405),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__10608 (
            .O(N__48402),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__10607 (
            .O(N__48399),
            .I(N__48396));
    LocalMux I__10606 (
            .O(N__48396),
            .I(N__48393));
    Odrv4 I__10605 (
            .O(N__48393),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    CascadeMux I__10604 (
            .O(N__48390),
            .I(N__48387));
    InMux I__10603 (
            .O(N__48387),
            .I(N__48384));
    LocalMux I__10602 (
            .O(N__48384),
            .I(N__48381));
    Odrv4 I__10601 (
            .O(N__48381),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    InMux I__10600 (
            .O(N__48378),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__10599 (
            .O(N__48375),
            .I(N__48372));
    LocalMux I__10598 (
            .O(N__48372),
            .I(N__48369));
    Odrv4 I__10597 (
            .O(N__48369),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    CascadeMux I__10596 (
            .O(N__48366),
            .I(N__48363));
    InMux I__10595 (
            .O(N__48363),
            .I(N__48360));
    LocalMux I__10594 (
            .O(N__48360),
            .I(N__48357));
    Odrv4 I__10593 (
            .O(N__48357),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__10592 (
            .O(N__48354),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__10591 (
            .O(N__48351),
            .I(N__48348));
    LocalMux I__10590 (
            .O(N__48348),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    CascadeMux I__10589 (
            .O(N__48345),
            .I(N__48342));
    InMux I__10588 (
            .O(N__48342),
            .I(N__48339));
    LocalMux I__10587 (
            .O(N__48339),
            .I(N__48336));
    Odrv4 I__10586 (
            .O(N__48336),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__10585 (
            .O(N__48333),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__10584 (
            .O(N__48330),
            .I(N__48327));
    LocalMux I__10583 (
            .O(N__48327),
            .I(N__48323));
    InMux I__10582 (
            .O(N__48326),
            .I(N__48320));
    Span4Mux_h I__10581 (
            .O(N__48323),
            .I(N__48317));
    LocalMux I__10580 (
            .O(N__48320),
            .I(N__48314));
    Span4Mux_v I__10579 (
            .O(N__48317),
            .I(N__48310));
    Span4Mux_h I__10578 (
            .O(N__48314),
            .I(N__48307));
    InMux I__10577 (
            .O(N__48313),
            .I(N__48304));
    Odrv4 I__10576 (
            .O(N__48310),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    Odrv4 I__10575 (
            .O(N__48307),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    LocalMux I__10574 (
            .O(N__48304),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    CascadeMux I__10573 (
            .O(N__48297),
            .I(N__48293));
    CascadeMux I__10572 (
            .O(N__48296),
            .I(N__48287));
    InMux I__10571 (
            .O(N__48293),
            .I(N__48282));
    InMux I__10570 (
            .O(N__48292),
            .I(N__48279));
    InMux I__10569 (
            .O(N__48291),
            .I(N__48276));
    InMux I__10568 (
            .O(N__48290),
            .I(N__48269));
    InMux I__10567 (
            .O(N__48287),
            .I(N__48269));
    InMux I__10566 (
            .O(N__48286),
            .I(N__48264));
    InMux I__10565 (
            .O(N__48285),
            .I(N__48264));
    LocalMux I__10564 (
            .O(N__48282),
            .I(N__48259));
    LocalMux I__10563 (
            .O(N__48279),
            .I(N__48259));
    LocalMux I__10562 (
            .O(N__48276),
            .I(N__48256));
    InMux I__10561 (
            .O(N__48275),
            .I(N__48251));
    InMux I__10560 (
            .O(N__48274),
            .I(N__48251));
    LocalMux I__10559 (
            .O(N__48269),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    LocalMux I__10558 (
            .O(N__48264),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    Odrv4 I__10557 (
            .O(N__48259),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    Odrv12 I__10556 (
            .O(N__48256),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    LocalMux I__10555 (
            .O(N__48251),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    InMux I__10554 (
            .O(N__48240),
            .I(N__48237));
    LocalMux I__10553 (
            .O(N__48237),
            .I(N__48233));
    InMux I__10552 (
            .O(N__48236),
            .I(N__48229));
    Span4Mux_h I__10551 (
            .O(N__48233),
            .I(N__48226));
    InMux I__10550 (
            .O(N__48232),
            .I(N__48223));
    LocalMux I__10549 (
            .O(N__48229),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv4 I__10548 (
            .O(N__48226),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    LocalMux I__10547 (
            .O(N__48223),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__10546 (
            .O(N__48216),
            .I(N__48213));
    LocalMux I__10545 (
            .O(N__48213),
            .I(N__48210));
    Span4Mux_v I__10544 (
            .O(N__48210),
            .I(N__48207));
    Odrv4 I__10543 (
            .O(N__48207),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ));
    CascadeMux I__10542 (
            .O(N__48204),
            .I(N__48201));
    InMux I__10541 (
            .O(N__48201),
            .I(N__48198));
    LocalMux I__10540 (
            .O(N__48198),
            .I(\ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ));
    InMux I__10539 (
            .O(N__48195),
            .I(N__48192));
    LocalMux I__10538 (
            .O(N__48192),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__10537 (
            .O(N__48189),
            .I(N__48186));
    LocalMux I__10536 (
            .O(N__48186),
            .I(N__48183));
    Span4Mux_h I__10535 (
            .O(N__48183),
            .I(N__48180));
    Odrv4 I__10534 (
            .O(N__48180),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__10533 (
            .O(N__48177),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__10532 (
            .O(N__48174),
            .I(N__48171));
    LocalMux I__10531 (
            .O(N__48171),
            .I(\ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ));
    CascadeMux I__10530 (
            .O(N__48168),
            .I(N__48165));
    InMux I__10529 (
            .O(N__48165),
            .I(N__48162));
    LocalMux I__10528 (
            .O(N__48162),
            .I(N__48159));
    Span4Mux_v I__10527 (
            .O(N__48159),
            .I(N__48156));
    Odrv4 I__10526 (
            .O(N__48156),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ));
    InMux I__10525 (
            .O(N__48153),
            .I(N__48150));
    LocalMux I__10524 (
            .O(N__48150),
            .I(N__48147));
    Span4Mux_v I__10523 (
            .O(N__48147),
            .I(N__48144));
    Odrv4 I__10522 (
            .O(N__48144),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    InMux I__10521 (
            .O(N__48141),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__10520 (
            .O(N__48138),
            .I(N__48135));
    LocalMux I__10519 (
            .O(N__48135),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__10518 (
            .O(N__48132),
            .I(N__48129));
    LocalMux I__10517 (
            .O(N__48129),
            .I(N__48126));
    Span4Mux_h I__10516 (
            .O(N__48126),
            .I(N__48123));
    Odrv4 I__10515 (
            .O(N__48123),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__10514 (
            .O(N__48120),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__10513 (
            .O(N__48117),
            .I(N__48114));
    LocalMux I__10512 (
            .O(N__48114),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__10511 (
            .O(N__48111),
            .I(N__48108));
    LocalMux I__10510 (
            .O(N__48108),
            .I(N__48105));
    Span4Mux_h I__10509 (
            .O(N__48105),
            .I(N__48102));
    Odrv4 I__10508 (
            .O(N__48102),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__10507 (
            .O(N__48099),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__10506 (
            .O(N__48096),
            .I(N__48093));
    LocalMux I__10505 (
            .O(N__48093),
            .I(\pid_side.m9_e_4 ));
    CascadeMux I__10504 (
            .O(N__48090),
            .I(\pid_side.m9_e_5_cascade_ ));
    InMux I__10503 (
            .O(N__48087),
            .I(N__48081));
    InMux I__10502 (
            .O(N__48086),
            .I(N__48074));
    InMux I__10501 (
            .O(N__48085),
            .I(N__48074));
    InMux I__10500 (
            .O(N__48084),
            .I(N__48074));
    LocalMux I__10499 (
            .O(N__48081),
            .I(\pid_side.pid_prereg_esr_RNIFB07Z0Z_20 ));
    LocalMux I__10498 (
            .O(N__48074),
            .I(\pid_side.pid_prereg_esr_RNIFB07Z0Z_20 ));
    CascadeMux I__10497 (
            .O(N__48069),
            .I(\pid_side.pid_prereg_esr_RNIFB07Z0Z_20_cascade_ ));
    InMux I__10496 (
            .O(N__48066),
            .I(N__48063));
    LocalMux I__10495 (
            .O(N__48063),
            .I(N__48059));
    InMux I__10494 (
            .O(N__48062),
            .I(N__48056));
    Span4Mux_h I__10493 (
            .O(N__48059),
            .I(N__48053));
    LocalMux I__10492 (
            .O(N__48056),
            .I(N__48050));
    Span4Mux_h I__10491 (
            .O(N__48053),
            .I(N__48047));
    Span12Mux_v I__10490 (
            .O(N__48050),
            .I(N__48044));
    Span4Mux_v I__10489 (
            .O(N__48047),
            .I(N__48041));
    Odrv12 I__10488 (
            .O(N__48044),
            .I(side_order_13));
    Odrv4 I__10487 (
            .O(N__48041),
            .I(side_order_13));
    CEMux I__10486 (
            .O(N__48036),
            .I(N__48032));
    CEMux I__10485 (
            .O(N__48035),
            .I(N__48029));
    LocalMux I__10484 (
            .O(N__48032),
            .I(N__48026));
    LocalMux I__10483 (
            .O(N__48029),
            .I(N__48022));
    Span4Mux_h I__10482 (
            .O(N__48026),
            .I(N__48017));
    CEMux I__10481 (
            .O(N__48025),
            .I(N__48014));
    Span4Mux_h I__10480 (
            .O(N__48022),
            .I(N__48011));
    CEMux I__10479 (
            .O(N__48021),
            .I(N__48008));
    CEMux I__10478 (
            .O(N__48020),
            .I(N__48005));
    Odrv4 I__10477 (
            .O(N__48017),
            .I(\pid_side.state_0_1 ));
    LocalMux I__10476 (
            .O(N__48014),
            .I(\pid_side.state_0_1 ));
    Odrv4 I__10475 (
            .O(N__48011),
            .I(\pid_side.state_0_1 ));
    LocalMux I__10474 (
            .O(N__48008),
            .I(\pid_side.state_0_1 ));
    LocalMux I__10473 (
            .O(N__48005),
            .I(\pid_side.state_0_1 ));
    SRMux I__10472 (
            .O(N__47994),
            .I(N__47991));
    LocalMux I__10471 (
            .O(N__47991),
            .I(N__47988));
    Span4Mux_v I__10470 (
            .O(N__47988),
            .I(N__47979));
    SRMux I__10469 (
            .O(N__47987),
            .I(N__47976));
    SRMux I__10468 (
            .O(N__47986),
            .I(N__47973));
    SRMux I__10467 (
            .O(N__47985),
            .I(N__47970));
    SRMux I__10466 (
            .O(N__47984),
            .I(N__47967));
    SRMux I__10465 (
            .O(N__47983),
            .I(N__47964));
    InMux I__10464 (
            .O(N__47982),
            .I(N__47961));
    Odrv4 I__10463 (
            .O(N__47979),
            .I(\pid_side.un1_reset_0_i ));
    LocalMux I__10462 (
            .O(N__47976),
            .I(\pid_side.un1_reset_0_i ));
    LocalMux I__10461 (
            .O(N__47973),
            .I(\pid_side.un1_reset_0_i ));
    LocalMux I__10460 (
            .O(N__47970),
            .I(\pid_side.un1_reset_0_i ));
    LocalMux I__10459 (
            .O(N__47967),
            .I(\pid_side.un1_reset_0_i ));
    LocalMux I__10458 (
            .O(N__47964),
            .I(\pid_side.un1_reset_0_i ));
    LocalMux I__10457 (
            .O(N__47961),
            .I(\pid_side.un1_reset_0_i ));
    CascadeMux I__10456 (
            .O(N__47946),
            .I(N__47942));
    InMux I__10455 (
            .O(N__47945),
            .I(N__47939));
    InMux I__10454 (
            .O(N__47942),
            .I(N__47936));
    LocalMux I__10453 (
            .O(N__47939),
            .I(N__47933));
    LocalMux I__10452 (
            .O(N__47936),
            .I(N__47930));
    Span4Mux_v I__10451 (
            .O(N__47933),
            .I(N__47927));
    Span4Mux_v I__10450 (
            .O(N__47930),
            .I(N__47924));
    Sp12to4 I__10449 (
            .O(N__47927),
            .I(N__47921));
    Sp12to4 I__10448 (
            .O(N__47924),
            .I(N__47916));
    Span12Mux_h I__10447 (
            .O(N__47921),
            .I(N__47916));
    Odrv12 I__10446 (
            .O(N__47916),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    InMux I__10445 (
            .O(N__47913),
            .I(N__47909));
    InMux I__10444 (
            .O(N__47912),
            .I(N__47906));
    LocalMux I__10443 (
            .O(N__47909),
            .I(N__47900));
    LocalMux I__10442 (
            .O(N__47906),
            .I(N__47900));
    InMux I__10441 (
            .O(N__47905),
            .I(N__47897));
    Span4Mux_v I__10440 (
            .O(N__47900),
            .I(N__47894));
    LocalMux I__10439 (
            .O(N__47897),
            .I(N__47891));
    Span4Mux_v I__10438 (
            .O(N__47894),
            .I(N__47888));
    Odrv4 I__10437 (
            .O(N__47891),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    Odrv4 I__10436 (
            .O(N__47888),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    InMux I__10435 (
            .O(N__47883),
            .I(N__47880));
    LocalMux I__10434 (
            .O(N__47880),
            .I(N__47877));
    Span4Mux_h I__10433 (
            .O(N__47877),
            .I(N__47874));
    Span4Mux_v I__10432 (
            .O(N__47874),
            .I(N__47866));
    InMux I__10431 (
            .O(N__47873),
            .I(N__47863));
    InMux I__10430 (
            .O(N__47872),
            .I(N__47854));
    InMux I__10429 (
            .O(N__47871),
            .I(N__47854));
    InMux I__10428 (
            .O(N__47870),
            .I(N__47854));
    InMux I__10427 (
            .O(N__47869),
            .I(N__47854));
    Odrv4 I__10426 (
            .O(N__47866),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__10425 (
            .O(N__47863),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__10424 (
            .O(N__47854),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    InMux I__10423 (
            .O(N__47847),
            .I(N__47844));
    LocalMux I__10422 (
            .O(N__47844),
            .I(N__47841));
    Span4Mux_h I__10421 (
            .O(N__47841),
            .I(N__47838));
    Span4Mux_v I__10420 (
            .O(N__47838),
            .I(N__47833));
    InMux I__10419 (
            .O(N__47837),
            .I(N__47828));
    InMux I__10418 (
            .O(N__47836),
            .I(N__47828));
    Odrv4 I__10417 (
            .O(N__47833),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__10416 (
            .O(N__47828),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    InMux I__10415 (
            .O(N__47823),
            .I(N__47819));
    CascadeMux I__10414 (
            .O(N__47822),
            .I(N__47816));
    LocalMux I__10413 (
            .O(N__47819),
            .I(N__47812));
    InMux I__10412 (
            .O(N__47816),
            .I(N__47809));
    InMux I__10411 (
            .O(N__47815),
            .I(N__47806));
    Span4Mux_h I__10410 (
            .O(N__47812),
            .I(N__47803));
    LocalMux I__10409 (
            .O(N__47809),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    LocalMux I__10408 (
            .O(N__47806),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    Odrv4 I__10407 (
            .O(N__47803),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    InMux I__10406 (
            .O(N__47796),
            .I(N__47793));
    LocalMux I__10405 (
            .O(N__47793),
            .I(N__47790));
    Span4Mux_h I__10404 (
            .O(N__47790),
            .I(N__47787));
    Span4Mux_h I__10403 (
            .O(N__47787),
            .I(N__47784));
    Odrv4 I__10402 (
            .O(N__47784),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    IoInMux I__10401 (
            .O(N__47781),
            .I(N__47778));
    LocalMux I__10400 (
            .O(N__47778),
            .I(N__47775));
    Span4Mux_s1_v I__10399 (
            .O(N__47775),
            .I(N__47772));
    Odrv4 I__10398 (
            .O(N__47772),
            .I(\pid_alt.N_664_0 ));
    InMux I__10397 (
            .O(N__47769),
            .I(N__47766));
    LocalMux I__10396 (
            .O(N__47766),
            .I(N__47763));
    Span4Mux_h I__10395 (
            .O(N__47763),
            .I(N__47758));
    InMux I__10394 (
            .O(N__47762),
            .I(N__47755));
    InMux I__10393 (
            .O(N__47761),
            .I(N__47752));
    Odrv4 I__10392 (
            .O(N__47758),
            .I(\pid_side.pid_preregZ0Z_0 ));
    LocalMux I__10391 (
            .O(N__47755),
            .I(\pid_side.pid_preregZ0Z_0 ));
    LocalMux I__10390 (
            .O(N__47752),
            .I(\pid_side.pid_preregZ0Z_0 ));
    InMux I__10389 (
            .O(N__47745),
            .I(N__47742));
    LocalMux I__10388 (
            .O(N__47742),
            .I(N__47738));
    CascadeMux I__10387 (
            .O(N__47741),
            .I(N__47735));
    Span4Mux_h I__10386 (
            .O(N__47738),
            .I(N__47732));
    InMux I__10385 (
            .O(N__47735),
            .I(N__47728));
    Span4Mux_v I__10384 (
            .O(N__47732),
            .I(N__47725));
    InMux I__10383 (
            .O(N__47731),
            .I(N__47722));
    LocalMux I__10382 (
            .O(N__47728),
            .I(\pid_side.pid_preregZ0Z_1 ));
    Odrv4 I__10381 (
            .O(N__47725),
            .I(\pid_side.pid_preregZ0Z_1 ));
    LocalMux I__10380 (
            .O(N__47722),
            .I(\pid_side.pid_preregZ0Z_1 ));
    IoInMux I__10379 (
            .O(N__47715),
            .I(N__47712));
    LocalMux I__10378 (
            .O(N__47712),
            .I(N__47706));
    InMux I__10377 (
            .O(N__47711),
            .I(N__47700));
    InMux I__10376 (
            .O(N__47710),
            .I(N__47700));
    InMux I__10375 (
            .O(N__47709),
            .I(N__47697));
    IoSpan4Mux I__10374 (
            .O(N__47706),
            .I(N__47694));
    InMux I__10373 (
            .O(N__47705),
            .I(N__47691));
    LocalMux I__10372 (
            .O(N__47700),
            .I(N__47688));
    LocalMux I__10371 (
            .O(N__47697),
            .I(N__47685));
    Span4Mux_s2_v I__10370 (
            .O(N__47694),
            .I(N__47681));
    LocalMux I__10369 (
            .O(N__47691),
            .I(N__47678));
    Span4Mux_v I__10368 (
            .O(N__47688),
            .I(N__47674));
    Span4Mux_h I__10367 (
            .O(N__47685),
            .I(N__47671));
    InMux I__10366 (
            .O(N__47684),
            .I(N__47668));
    Span4Mux_v I__10365 (
            .O(N__47681),
            .I(N__47665));
    Span4Mux_h I__10364 (
            .O(N__47678),
            .I(N__47662));
    InMux I__10363 (
            .O(N__47677),
            .I(N__47658));
    Sp12to4 I__10362 (
            .O(N__47674),
            .I(N__47655));
    Sp12to4 I__10361 (
            .O(N__47671),
            .I(N__47652));
    LocalMux I__10360 (
            .O(N__47668),
            .I(N__47649));
    Span4Mux_v I__10359 (
            .O(N__47665),
            .I(N__47644));
    Span4Mux_h I__10358 (
            .O(N__47662),
            .I(N__47644));
    InMux I__10357 (
            .O(N__47661),
            .I(N__47641));
    LocalMux I__10356 (
            .O(N__47658),
            .I(N__47636));
    Span12Mux_h I__10355 (
            .O(N__47655),
            .I(N__47636));
    Span12Mux_v I__10354 (
            .O(N__47652),
            .I(N__47631));
    Span12Mux_v I__10353 (
            .O(N__47649),
            .I(N__47631));
    Odrv4 I__10352 (
            .O(N__47644),
            .I(debug_CH1_0A_c));
    LocalMux I__10351 (
            .O(N__47641),
            .I(debug_CH1_0A_c));
    Odrv12 I__10350 (
            .O(N__47636),
            .I(debug_CH1_0A_c));
    Odrv12 I__10349 (
            .O(N__47631),
            .I(debug_CH1_0A_c));
    CascadeMux I__10348 (
            .O(N__47622),
            .I(N__47614));
    InMux I__10347 (
            .O(N__47621),
            .I(N__47611));
    InMux I__10346 (
            .O(N__47620),
            .I(N__47600));
    InMux I__10345 (
            .O(N__47619),
            .I(N__47600));
    InMux I__10344 (
            .O(N__47618),
            .I(N__47600));
    InMux I__10343 (
            .O(N__47617),
            .I(N__47600));
    InMux I__10342 (
            .O(N__47614),
            .I(N__47600));
    LocalMux I__10341 (
            .O(N__47611),
            .I(N__47597));
    LocalMux I__10340 (
            .O(N__47600),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv12 I__10339 (
            .O(N__47597),
            .I(\pid_side.stateZ0Z_0 ));
    InMux I__10338 (
            .O(N__47592),
            .I(N__47589));
    LocalMux I__10337 (
            .O(N__47589),
            .I(N__47586));
    Odrv4 I__10336 (
            .O(N__47586),
            .I(\pid_side.m18_s_5 ));
    InMux I__10335 (
            .O(N__47583),
            .I(N__47564));
    InMux I__10334 (
            .O(N__47582),
            .I(N__47564));
    InMux I__10333 (
            .O(N__47581),
            .I(N__47564));
    InMux I__10332 (
            .O(N__47580),
            .I(N__47564));
    InMux I__10331 (
            .O(N__47579),
            .I(N__47564));
    InMux I__10330 (
            .O(N__47578),
            .I(N__47564));
    InMux I__10329 (
            .O(N__47577),
            .I(N__47561));
    LocalMux I__10328 (
            .O(N__47564),
            .I(N__47558));
    LocalMux I__10327 (
            .O(N__47561),
            .I(N__47555));
    Span4Mux_h I__10326 (
            .O(N__47558),
            .I(N__47548));
    Span4Mux_h I__10325 (
            .O(N__47555),
            .I(N__47545));
    InMux I__10324 (
            .O(N__47554),
            .I(N__47540));
    InMux I__10323 (
            .O(N__47553),
            .I(N__47540));
    InMux I__10322 (
            .O(N__47552),
            .I(N__47537));
    InMux I__10321 (
            .O(N__47551),
            .I(N__47534));
    Odrv4 I__10320 (
            .O(N__47548),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__10319 (
            .O(N__47545),
            .I(\pid_side.stateZ0Z_1 ));
    LocalMux I__10318 (
            .O(N__47540),
            .I(\pid_side.stateZ0Z_1 ));
    LocalMux I__10317 (
            .O(N__47537),
            .I(\pid_side.stateZ0Z_1 ));
    LocalMux I__10316 (
            .O(N__47534),
            .I(\pid_side.stateZ0Z_1 ));
    InMux I__10315 (
            .O(N__47523),
            .I(N__47520));
    LocalMux I__10314 (
            .O(N__47520),
            .I(\pid_side.un1_reset_0_i_rn_0 ));
    InMux I__10313 (
            .O(N__47517),
            .I(N__47514));
    LocalMux I__10312 (
            .O(N__47514),
            .I(\pid_side.m26_e_1 ));
    InMux I__10311 (
            .O(N__47511),
            .I(N__47508));
    LocalMux I__10310 (
            .O(N__47508),
            .I(N__47505));
    Span4Mux_v I__10309 (
            .O(N__47505),
            .I(N__47502));
    Odrv4 I__10308 (
            .O(N__47502),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ));
    InMux I__10307 (
            .O(N__47499),
            .I(N__47496));
    LocalMux I__10306 (
            .O(N__47496),
            .I(N__47493));
    Odrv4 I__10305 (
            .O(N__47493),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__10304 (
            .O(N__47490),
            .I(N__47487));
    LocalMux I__10303 (
            .O(N__47487),
            .I(N__47484));
    Span4Mux_v I__10302 (
            .O(N__47484),
            .I(N__47480));
    InMux I__10301 (
            .O(N__47483),
            .I(N__47477));
    Span4Mux_v I__10300 (
            .O(N__47480),
            .I(N__47472));
    LocalMux I__10299 (
            .O(N__47477),
            .I(N__47472));
    Odrv4 I__10298 (
            .O(N__47472),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    InMux I__10297 (
            .O(N__47469),
            .I(N__47458));
    InMux I__10296 (
            .O(N__47468),
            .I(N__47453));
    InMux I__10295 (
            .O(N__47467),
            .I(N__47448));
    InMux I__10294 (
            .O(N__47466),
            .I(N__47448));
    InMux I__10293 (
            .O(N__47465),
            .I(N__47441));
    InMux I__10292 (
            .O(N__47464),
            .I(N__47441));
    InMux I__10291 (
            .O(N__47463),
            .I(N__47441));
    InMux I__10290 (
            .O(N__47462),
            .I(N__47436));
    InMux I__10289 (
            .O(N__47461),
            .I(N__47436));
    LocalMux I__10288 (
            .O(N__47458),
            .I(N__47433));
    InMux I__10287 (
            .O(N__47457),
            .I(N__47428));
    InMux I__10286 (
            .O(N__47456),
            .I(N__47428));
    LocalMux I__10285 (
            .O(N__47453),
            .I(N__47425));
    LocalMux I__10284 (
            .O(N__47448),
            .I(N__47410));
    LocalMux I__10283 (
            .O(N__47441),
            .I(N__47410));
    LocalMux I__10282 (
            .O(N__47436),
            .I(N__47410));
    Span4Mux_h I__10281 (
            .O(N__47433),
            .I(N__47407));
    LocalMux I__10280 (
            .O(N__47428),
            .I(N__47404));
    Span4Mux_h I__10279 (
            .O(N__47425),
            .I(N__47401));
    InMux I__10278 (
            .O(N__47424),
            .I(N__47394));
    InMux I__10277 (
            .O(N__47423),
            .I(N__47394));
    InMux I__10276 (
            .O(N__47422),
            .I(N__47394));
    InMux I__10275 (
            .O(N__47421),
            .I(N__47387));
    InMux I__10274 (
            .O(N__47420),
            .I(N__47387));
    InMux I__10273 (
            .O(N__47419),
            .I(N__47387));
    InMux I__10272 (
            .O(N__47418),
            .I(N__47384));
    InMux I__10271 (
            .O(N__47417),
            .I(N__47381));
    Span4Mux_v I__10270 (
            .O(N__47410),
            .I(N__47378));
    Span4Mux_v I__10269 (
            .O(N__47407),
            .I(N__47375));
    Span4Mux_h I__10268 (
            .O(N__47404),
            .I(N__47372));
    Span4Mux_v I__10267 (
            .O(N__47401),
            .I(N__47369));
    LocalMux I__10266 (
            .O(N__47394),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__10265 (
            .O(N__47387),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__10264 (
            .O(N__47384),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__10263 (
            .O(N__47381),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__10262 (
            .O(N__47378),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__10261 (
            .O(N__47375),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__10260 (
            .O(N__47372),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__10259 (
            .O(N__47369),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    CascadeMux I__10258 (
            .O(N__47352),
            .I(N__47340));
    CascadeMux I__10257 (
            .O(N__47351),
            .I(N__47337));
    CascadeMux I__10256 (
            .O(N__47350),
            .I(N__47334));
    CascadeMux I__10255 (
            .O(N__47349),
            .I(N__47331));
    CascadeMux I__10254 (
            .O(N__47348),
            .I(N__47328));
    CascadeMux I__10253 (
            .O(N__47347),
            .I(N__47324));
    CascadeMux I__10252 (
            .O(N__47346),
            .I(N__47321));
    InMux I__10251 (
            .O(N__47345),
            .I(N__47308));
    InMux I__10250 (
            .O(N__47344),
            .I(N__47308));
    InMux I__10249 (
            .O(N__47343),
            .I(N__47308));
    InMux I__10248 (
            .O(N__47340),
            .I(N__47301));
    InMux I__10247 (
            .O(N__47337),
            .I(N__47301));
    InMux I__10246 (
            .O(N__47334),
            .I(N__47301));
    InMux I__10245 (
            .O(N__47331),
            .I(N__47298));
    InMux I__10244 (
            .O(N__47328),
            .I(N__47295));
    InMux I__10243 (
            .O(N__47327),
            .I(N__47292));
    InMux I__10242 (
            .O(N__47324),
            .I(N__47287));
    InMux I__10241 (
            .O(N__47321),
            .I(N__47287));
    CascadeMux I__10240 (
            .O(N__47320),
            .I(N__47284));
    CascadeMux I__10239 (
            .O(N__47319),
            .I(N__47281));
    CascadeMux I__10238 (
            .O(N__47318),
            .I(N__47278));
    CascadeMux I__10237 (
            .O(N__47317),
            .I(N__47274));
    CascadeMux I__10236 (
            .O(N__47316),
            .I(N__47271));
    CascadeMux I__10235 (
            .O(N__47315),
            .I(N__47268));
    LocalMux I__10234 (
            .O(N__47308),
            .I(N__47265));
    LocalMux I__10233 (
            .O(N__47301),
            .I(N__47256));
    LocalMux I__10232 (
            .O(N__47298),
            .I(N__47256));
    LocalMux I__10231 (
            .O(N__47295),
            .I(N__47256));
    LocalMux I__10230 (
            .O(N__47292),
            .I(N__47256));
    LocalMux I__10229 (
            .O(N__47287),
            .I(N__47253));
    InMux I__10228 (
            .O(N__47284),
            .I(N__47248));
    InMux I__10227 (
            .O(N__47281),
            .I(N__47248));
    InMux I__10226 (
            .O(N__47278),
            .I(N__47245));
    InMux I__10225 (
            .O(N__47277),
            .I(N__47242));
    InMux I__10224 (
            .O(N__47274),
            .I(N__47236));
    InMux I__10223 (
            .O(N__47271),
            .I(N__47236));
    InMux I__10222 (
            .O(N__47268),
            .I(N__47233));
    Span4Mux_v I__10221 (
            .O(N__47265),
            .I(N__47230));
    Span4Mux_v I__10220 (
            .O(N__47256),
            .I(N__47225));
    Span4Mux_h I__10219 (
            .O(N__47253),
            .I(N__47225));
    LocalMux I__10218 (
            .O(N__47248),
            .I(N__47218));
    LocalMux I__10217 (
            .O(N__47245),
            .I(N__47218));
    LocalMux I__10216 (
            .O(N__47242),
            .I(N__47218));
    InMux I__10215 (
            .O(N__47241),
            .I(N__47215));
    LocalMux I__10214 (
            .O(N__47236),
            .I(N__47210));
    LocalMux I__10213 (
            .O(N__47233),
            .I(N__47210));
    Odrv4 I__10212 (
            .O(N__47230),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__10211 (
            .O(N__47225),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv12 I__10210 (
            .O(N__47218),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__10209 (
            .O(N__47215),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__10208 (
            .O(N__47210),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    InMux I__10207 (
            .O(N__47199),
            .I(N__47196));
    LocalMux I__10206 (
            .O(N__47196),
            .I(N__47193));
    Odrv4 I__10205 (
            .O(N__47193),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__10204 (
            .O(N__47190),
            .I(N__47181));
    InMux I__10203 (
            .O(N__47189),
            .I(N__47181));
    InMux I__10202 (
            .O(N__47188),
            .I(N__47181));
    LocalMux I__10201 (
            .O(N__47181),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__10200 (
            .O(N__47178),
            .I(N__47174));
    InMux I__10199 (
            .O(N__47177),
            .I(N__47166));
    LocalMux I__10198 (
            .O(N__47174),
            .I(N__47158));
    InMux I__10197 (
            .O(N__47173),
            .I(N__47153));
    InMux I__10196 (
            .O(N__47172),
            .I(N__47153));
    InMux I__10195 (
            .O(N__47171),
            .I(N__47147));
    InMux I__10194 (
            .O(N__47170),
            .I(N__47144));
    InMux I__10193 (
            .O(N__47169),
            .I(N__47141));
    LocalMux I__10192 (
            .O(N__47166),
            .I(N__47138));
    InMux I__10191 (
            .O(N__47165),
            .I(N__47135));
    InMux I__10190 (
            .O(N__47164),
            .I(N__47132));
    InMux I__10189 (
            .O(N__47163),
            .I(N__47129));
    InMux I__10188 (
            .O(N__47162),
            .I(N__47123));
    InMux I__10187 (
            .O(N__47161),
            .I(N__47120));
    Span4Mux_h I__10186 (
            .O(N__47158),
            .I(N__47115));
    LocalMux I__10185 (
            .O(N__47153),
            .I(N__47115));
    InMux I__10184 (
            .O(N__47152),
            .I(N__47110));
    InMux I__10183 (
            .O(N__47151),
            .I(N__47110));
    InMux I__10182 (
            .O(N__47150),
            .I(N__47106));
    LocalMux I__10181 (
            .O(N__47147),
            .I(N__47093));
    LocalMux I__10180 (
            .O(N__47144),
            .I(N__47093));
    LocalMux I__10179 (
            .O(N__47141),
            .I(N__47093));
    Span4Mux_v I__10178 (
            .O(N__47138),
            .I(N__47093));
    LocalMux I__10177 (
            .O(N__47135),
            .I(N__47093));
    LocalMux I__10176 (
            .O(N__47132),
            .I(N__47093));
    LocalMux I__10175 (
            .O(N__47129),
            .I(N__47090));
    InMux I__10174 (
            .O(N__47128),
            .I(N__47087));
    InMux I__10173 (
            .O(N__47127),
            .I(N__47084));
    InMux I__10172 (
            .O(N__47126),
            .I(N__47081));
    LocalMux I__10171 (
            .O(N__47123),
            .I(N__47072));
    LocalMux I__10170 (
            .O(N__47120),
            .I(N__47072));
    Span4Mux_v I__10169 (
            .O(N__47115),
            .I(N__47072));
    LocalMux I__10168 (
            .O(N__47110),
            .I(N__47072));
    InMux I__10167 (
            .O(N__47109),
            .I(N__47069));
    LocalMux I__10166 (
            .O(N__47106),
            .I(N__47064));
    Span4Mux_v I__10165 (
            .O(N__47093),
            .I(N__47064));
    Span4Mux_h I__10164 (
            .O(N__47090),
            .I(N__47061));
    LocalMux I__10163 (
            .O(N__47087),
            .I(N__47054));
    LocalMux I__10162 (
            .O(N__47084),
            .I(N__47054));
    LocalMux I__10161 (
            .O(N__47081),
            .I(N__47054));
    Span4Mux_v I__10160 (
            .O(N__47072),
            .I(N__47051));
    LocalMux I__10159 (
            .O(N__47069),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__10158 (
            .O(N__47064),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__10157 (
            .O(N__47061),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__10156 (
            .O(N__47054),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__10155 (
            .O(N__47051),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__10154 (
            .O(N__47040),
            .I(N__47036));
    InMux I__10153 (
            .O(N__47039),
            .I(N__47033));
    LocalMux I__10152 (
            .O(N__47036),
            .I(N__47029));
    LocalMux I__10151 (
            .O(N__47033),
            .I(N__47026));
    CascadeMux I__10150 (
            .O(N__47032),
            .I(N__47023));
    Span4Mux_h I__10149 (
            .O(N__47029),
            .I(N__47020));
    Span4Mux_h I__10148 (
            .O(N__47026),
            .I(N__47017));
    InMux I__10147 (
            .O(N__47023),
            .I(N__47014));
    Span4Mux_h I__10146 (
            .O(N__47020),
            .I(N__47009));
    Span4Mux_h I__10145 (
            .O(N__47017),
            .I(N__47009));
    LocalMux I__10144 (
            .O(N__47014),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    Odrv4 I__10143 (
            .O(N__47009),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    InMux I__10142 (
            .O(N__47004),
            .I(N__47001));
    LocalMux I__10141 (
            .O(N__47001),
            .I(N__46997));
    InMux I__10140 (
            .O(N__47000),
            .I(N__46994));
    Span4Mux_v I__10139 (
            .O(N__46997),
            .I(N__46988));
    LocalMux I__10138 (
            .O(N__46994),
            .I(N__46988));
    InMux I__10137 (
            .O(N__46993),
            .I(N__46985));
    Span4Mux_h I__10136 (
            .O(N__46988),
            .I(N__46982));
    LocalMux I__10135 (
            .O(N__46985),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv4 I__10134 (
            .O(N__46982),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    InMux I__10133 (
            .O(N__46977),
            .I(N__46974));
    LocalMux I__10132 (
            .O(N__46974),
            .I(N__46971));
    Odrv12 I__10131 (
            .O(N__46971),
            .I(\ppm_encoder_1.N_288 ));
    InMux I__10130 (
            .O(N__46968),
            .I(N__46965));
    LocalMux I__10129 (
            .O(N__46965),
            .I(N__46962));
    Odrv4 I__10128 (
            .O(N__46962),
            .I(\ppm_encoder_1.N_290 ));
    InMux I__10127 (
            .O(N__46959),
            .I(N__46956));
    LocalMux I__10126 (
            .O(N__46956),
            .I(N__46953));
    Span4Mux_h I__10125 (
            .O(N__46953),
            .I(N__46948));
    InMux I__10124 (
            .O(N__46952),
            .I(N__46945));
    InMux I__10123 (
            .O(N__46951),
            .I(N__46942));
    Span4Mux_v I__10122 (
            .O(N__46948),
            .I(N__46937));
    LocalMux I__10121 (
            .O(N__46945),
            .I(N__46937));
    LocalMux I__10120 (
            .O(N__46942),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    Odrv4 I__10119 (
            .O(N__46937),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    InMux I__10118 (
            .O(N__46932),
            .I(N__46929));
    LocalMux I__10117 (
            .O(N__46929),
            .I(N__46926));
    Span4Mux_v I__10116 (
            .O(N__46926),
            .I(N__46923));
    Odrv4 I__10115 (
            .O(N__46923),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ));
    InMux I__10114 (
            .O(N__46920),
            .I(N__46914));
    InMux I__10113 (
            .O(N__46919),
            .I(N__46914));
    LocalMux I__10112 (
            .O(N__46914),
            .I(N__46911));
    Odrv12 I__10111 (
            .O(N__46911),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    InMux I__10110 (
            .O(N__46908),
            .I(N__46901));
    InMux I__10109 (
            .O(N__46907),
            .I(N__46901));
    CascadeMux I__10108 (
            .O(N__46906),
            .I(N__46897));
    LocalMux I__10107 (
            .O(N__46901),
            .I(N__46894));
    InMux I__10106 (
            .O(N__46900),
            .I(N__46891));
    InMux I__10105 (
            .O(N__46897),
            .I(N__46888));
    Span4Mux_h I__10104 (
            .O(N__46894),
            .I(N__46885));
    LocalMux I__10103 (
            .O(N__46891),
            .I(N__46880));
    LocalMux I__10102 (
            .O(N__46888),
            .I(N__46880));
    Span4Mux_v I__10101 (
            .O(N__46885),
            .I(N__46875));
    Span4Mux_v I__10100 (
            .O(N__46880),
            .I(N__46875));
    Span4Mux_v I__10099 (
            .O(N__46875),
            .I(N__46872));
    Odrv4 I__10098 (
            .O(N__46872),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ));
    CascadeMux I__10097 (
            .O(N__46869),
            .I(N__46866));
    InMux I__10096 (
            .O(N__46866),
            .I(N__46862));
    InMux I__10095 (
            .O(N__46865),
            .I(N__46859));
    LocalMux I__10094 (
            .O(N__46862),
            .I(N__46856));
    LocalMux I__10093 (
            .O(N__46859),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    Odrv12 I__10092 (
            .O(N__46856),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    InMux I__10091 (
            .O(N__46851),
            .I(N__46847));
    InMux I__10090 (
            .O(N__46850),
            .I(N__46844));
    LocalMux I__10089 (
            .O(N__46847),
            .I(N__46841));
    LocalMux I__10088 (
            .O(N__46844),
            .I(N__46838));
    Span4Mux_v I__10087 (
            .O(N__46841),
            .I(N__46835));
    Span12Mux_v I__10086 (
            .O(N__46838),
            .I(N__46832));
    Span4Mux_h I__10085 (
            .O(N__46835),
            .I(N__46829));
    Odrv12 I__10084 (
            .O(N__46832),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    Odrv4 I__10083 (
            .O(N__46829),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    InMux I__10082 (
            .O(N__46824),
            .I(N__46821));
    LocalMux I__10081 (
            .O(N__46821),
            .I(N__46818));
    Span4Mux_h I__10080 (
            .O(N__46818),
            .I(N__46814));
    CascadeMux I__10079 (
            .O(N__46817),
            .I(N__46811));
    Span4Mux_v I__10078 (
            .O(N__46814),
            .I(N__46808));
    InMux I__10077 (
            .O(N__46811),
            .I(N__46805));
    Odrv4 I__10076 (
            .O(N__46808),
            .I(scaler_4_data_4));
    LocalMux I__10075 (
            .O(N__46805),
            .I(scaler_4_data_4));
    InMux I__10074 (
            .O(N__46800),
            .I(N__46797));
    LocalMux I__10073 (
            .O(N__46797),
            .I(N__46793));
    InMux I__10072 (
            .O(N__46796),
            .I(N__46790));
    Span4Mux_h I__10071 (
            .O(N__46793),
            .I(N__46787));
    LocalMux I__10070 (
            .O(N__46790),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    Odrv4 I__10069 (
            .O(N__46787),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    CEMux I__10068 (
            .O(N__46782),
            .I(N__46778));
    CEMux I__10067 (
            .O(N__46781),
            .I(N__46773));
    LocalMux I__10066 (
            .O(N__46778),
            .I(N__46770));
    CEMux I__10065 (
            .O(N__46777),
            .I(N__46767));
    CEMux I__10064 (
            .O(N__46776),
            .I(N__46764));
    LocalMux I__10063 (
            .O(N__46773),
            .I(N__46759));
    Span4Mux_h I__10062 (
            .O(N__46770),
            .I(N__46754));
    LocalMux I__10061 (
            .O(N__46767),
            .I(N__46754));
    LocalMux I__10060 (
            .O(N__46764),
            .I(N__46751));
    CEMux I__10059 (
            .O(N__46763),
            .I(N__46748));
    CEMux I__10058 (
            .O(N__46762),
            .I(N__46745));
    Span4Mux_v I__10057 (
            .O(N__46759),
            .I(N__46742));
    Span4Mux_v I__10056 (
            .O(N__46754),
            .I(N__46735));
    Span4Mux_v I__10055 (
            .O(N__46751),
            .I(N__46735));
    LocalMux I__10054 (
            .O(N__46748),
            .I(N__46735));
    LocalMux I__10053 (
            .O(N__46745),
            .I(N__46732));
    Span4Mux_h I__10052 (
            .O(N__46742),
            .I(N__46727));
    Span4Mux_h I__10051 (
            .O(N__46735),
            .I(N__46727));
    Span4Mux_v I__10050 (
            .O(N__46732),
            .I(N__46724));
    Span4Mux_h I__10049 (
            .O(N__46727),
            .I(N__46721));
    Odrv4 I__10048 (
            .O(N__46724),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__10047 (
            .O(N__46721),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    InMux I__10046 (
            .O(N__46716),
            .I(N__46713));
    LocalMux I__10045 (
            .O(N__46713),
            .I(N__46709));
    InMux I__10044 (
            .O(N__46712),
            .I(N__46705));
    Span12Mux_v I__10043 (
            .O(N__46709),
            .I(N__46702));
    InMux I__10042 (
            .O(N__46708),
            .I(N__46699));
    LocalMux I__10041 (
            .O(N__46705),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv12 I__10040 (
            .O(N__46702),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    LocalMux I__10039 (
            .O(N__46699),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    CascadeMux I__10038 (
            .O(N__46692),
            .I(\ppm_encoder_1.N_314_cascade_ ));
    CascadeMux I__10037 (
            .O(N__46689),
            .I(N__46686));
    InMux I__10036 (
            .O(N__46686),
            .I(N__46677));
    InMux I__10035 (
            .O(N__46685),
            .I(N__46677));
    InMux I__10034 (
            .O(N__46684),
            .I(N__46677));
    LocalMux I__10033 (
            .O(N__46677),
            .I(N__46673));
    InMux I__10032 (
            .O(N__46676),
            .I(N__46670));
    Sp12to4 I__10031 (
            .O(N__46673),
            .I(N__46665));
    LocalMux I__10030 (
            .O(N__46670),
            .I(N__46665));
    Span12Mux_s10_h I__10029 (
            .O(N__46665),
            .I(N__46661));
    InMux I__10028 (
            .O(N__46664),
            .I(N__46658));
    Odrv12 I__10027 (
            .O(N__46661),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    LocalMux I__10026 (
            .O(N__46658),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    InMux I__10025 (
            .O(N__46653),
            .I(N__46650));
    LocalMux I__10024 (
            .O(N__46650),
            .I(N__46647));
    Span4Mux_h I__10023 (
            .O(N__46647),
            .I(N__46644));
    Odrv4 I__10022 (
            .O(N__46644),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ));
    InMux I__10021 (
            .O(N__46641),
            .I(N__46638));
    LocalMux I__10020 (
            .O(N__46638),
            .I(N__46634));
    InMux I__10019 (
            .O(N__46637),
            .I(N__46631));
    Span4Mux_h I__10018 (
            .O(N__46634),
            .I(N__46628));
    LocalMux I__10017 (
            .O(N__46631),
            .I(N__46625));
    Span4Mux_v I__10016 (
            .O(N__46628),
            .I(N__46620));
    Span4Mux_v I__10015 (
            .O(N__46625),
            .I(N__46620));
    Odrv4 I__10014 (
            .O(N__46620),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    InMux I__10013 (
            .O(N__46617),
            .I(N__46614));
    LocalMux I__10012 (
            .O(N__46614),
            .I(N__46611));
    Odrv4 I__10011 (
            .O(N__46611),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__10010 (
            .O(N__46608),
            .I(N__46605));
    LocalMux I__10009 (
            .O(N__46605),
            .I(N__46601));
    InMux I__10008 (
            .O(N__46604),
            .I(N__46598));
    Span4Mux_h I__10007 (
            .O(N__46601),
            .I(N__46595));
    LocalMux I__10006 (
            .O(N__46598),
            .I(N__46592));
    Odrv4 I__10005 (
            .O(N__46595),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    Odrv4 I__10004 (
            .O(N__46592),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    InMux I__10003 (
            .O(N__46587),
            .I(N__46578));
    InMux I__10002 (
            .O(N__46586),
            .I(N__46578));
    InMux I__10001 (
            .O(N__46585),
            .I(N__46578));
    LocalMux I__10000 (
            .O(N__46578),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__9999 (
            .O(N__46575),
            .I(N__46561));
    InMux I__9998 (
            .O(N__46574),
            .I(N__46558));
    InMux I__9997 (
            .O(N__46573),
            .I(N__46555));
    CascadeMux I__9996 (
            .O(N__46572),
            .I(N__46550));
    InMux I__9995 (
            .O(N__46571),
            .I(N__46547));
    InMux I__9994 (
            .O(N__46570),
            .I(N__46544));
    InMux I__9993 (
            .O(N__46569),
            .I(N__46541));
    InMux I__9992 (
            .O(N__46568),
            .I(N__46536));
    InMux I__9991 (
            .O(N__46567),
            .I(N__46536));
    InMux I__9990 (
            .O(N__46566),
            .I(N__46531));
    InMux I__9989 (
            .O(N__46565),
            .I(N__46531));
    InMux I__9988 (
            .O(N__46564),
            .I(N__46528));
    LocalMux I__9987 (
            .O(N__46561),
            .I(N__46525));
    LocalMux I__9986 (
            .O(N__46558),
            .I(N__46520));
    LocalMux I__9985 (
            .O(N__46555),
            .I(N__46520));
    InMux I__9984 (
            .O(N__46554),
            .I(N__46513));
    InMux I__9983 (
            .O(N__46553),
            .I(N__46513));
    InMux I__9982 (
            .O(N__46550),
            .I(N__46513));
    LocalMux I__9981 (
            .O(N__46547),
            .I(N__46510));
    LocalMux I__9980 (
            .O(N__46544),
            .I(N__46505));
    LocalMux I__9979 (
            .O(N__46541),
            .I(N__46505));
    LocalMux I__9978 (
            .O(N__46536),
            .I(N__46502));
    LocalMux I__9977 (
            .O(N__46531),
            .I(N__46498));
    LocalMux I__9976 (
            .O(N__46528),
            .I(N__46495));
    Span4Mux_v I__9975 (
            .O(N__46525),
            .I(N__46492));
    Span4Mux_v I__9974 (
            .O(N__46520),
            .I(N__46485));
    LocalMux I__9973 (
            .O(N__46513),
            .I(N__46485));
    Span4Mux_h I__9972 (
            .O(N__46510),
            .I(N__46485));
    Span4Mux_v I__9971 (
            .O(N__46505),
            .I(N__46480));
    Span4Mux_h I__9970 (
            .O(N__46502),
            .I(N__46480));
    InMux I__9969 (
            .O(N__46501),
            .I(N__46477));
    Span4Mux_v I__9968 (
            .O(N__46498),
            .I(N__46470));
    Span4Mux_v I__9967 (
            .O(N__46495),
            .I(N__46470));
    Span4Mux_h I__9966 (
            .O(N__46492),
            .I(N__46470));
    Span4Mux_v I__9965 (
            .O(N__46485),
            .I(N__46467));
    Span4Mux_v I__9964 (
            .O(N__46480),
            .I(N__46464));
    LocalMux I__9963 (
            .O(N__46477),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__9962 (
            .O(N__46470),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__9961 (
            .O(N__46467),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__9960 (
            .O(N__46464),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    CascadeMux I__9959 (
            .O(N__46455),
            .I(N__46450));
    CascadeMux I__9958 (
            .O(N__46454),
            .I(N__46441));
    CascadeMux I__9957 (
            .O(N__46453),
            .I(N__46438));
    InMux I__9956 (
            .O(N__46450),
            .I(N__46433));
    InMux I__9955 (
            .O(N__46449),
            .I(N__46426));
    InMux I__9954 (
            .O(N__46448),
            .I(N__46426));
    InMux I__9953 (
            .O(N__46447),
            .I(N__46426));
    CascadeMux I__9952 (
            .O(N__46446),
            .I(N__46423));
    CascadeMux I__9951 (
            .O(N__46445),
            .I(N__46420));
    CascadeMux I__9950 (
            .O(N__46444),
            .I(N__46417));
    InMux I__9949 (
            .O(N__46441),
            .I(N__46414));
    InMux I__9948 (
            .O(N__46438),
            .I(N__46411));
    CascadeMux I__9947 (
            .O(N__46437),
            .I(N__46408));
    InMux I__9946 (
            .O(N__46436),
            .I(N__46404));
    LocalMux I__9945 (
            .O(N__46433),
            .I(N__46399));
    LocalMux I__9944 (
            .O(N__46426),
            .I(N__46399));
    InMux I__9943 (
            .O(N__46423),
            .I(N__46396));
    InMux I__9942 (
            .O(N__46420),
            .I(N__46393));
    InMux I__9941 (
            .O(N__46417),
            .I(N__46390));
    LocalMux I__9940 (
            .O(N__46414),
            .I(N__46383));
    LocalMux I__9939 (
            .O(N__46411),
            .I(N__46383));
    InMux I__9938 (
            .O(N__46408),
            .I(N__46378));
    InMux I__9937 (
            .O(N__46407),
            .I(N__46378));
    LocalMux I__9936 (
            .O(N__46404),
            .I(N__46371));
    Span4Mux_v I__9935 (
            .O(N__46399),
            .I(N__46371));
    LocalMux I__9934 (
            .O(N__46396),
            .I(N__46371));
    LocalMux I__9933 (
            .O(N__46393),
            .I(N__46366));
    LocalMux I__9932 (
            .O(N__46390),
            .I(N__46366));
    InMux I__9931 (
            .O(N__46389),
            .I(N__46361));
    InMux I__9930 (
            .O(N__46388),
            .I(N__46361));
    Span4Mux_v I__9929 (
            .O(N__46383),
            .I(N__46357));
    LocalMux I__9928 (
            .O(N__46378),
            .I(N__46354));
    Span4Mux_v I__9927 (
            .O(N__46371),
            .I(N__46349));
    Span4Mux_v I__9926 (
            .O(N__46366),
            .I(N__46344));
    LocalMux I__9925 (
            .O(N__46361),
            .I(N__46344));
    InMux I__9924 (
            .O(N__46360),
            .I(N__46341));
    Span4Mux_h I__9923 (
            .O(N__46357),
            .I(N__46336));
    Span4Mux_h I__9922 (
            .O(N__46354),
            .I(N__46336));
    CascadeMux I__9921 (
            .O(N__46353),
            .I(N__46333));
    InMux I__9920 (
            .O(N__46352),
            .I(N__46329));
    Span4Mux_h I__9919 (
            .O(N__46349),
            .I(N__46326));
    Sp12to4 I__9918 (
            .O(N__46344),
            .I(N__46323));
    LocalMux I__9917 (
            .O(N__46341),
            .I(N__46318));
    Span4Mux_v I__9916 (
            .O(N__46336),
            .I(N__46318));
    InMux I__9915 (
            .O(N__46333),
            .I(N__46313));
    InMux I__9914 (
            .O(N__46332),
            .I(N__46313));
    LocalMux I__9913 (
            .O(N__46329),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__9912 (
            .O(N__46326),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv12 I__9911 (
            .O(N__46323),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__9910 (
            .O(N__46318),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__9909 (
            .O(N__46313),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__9908 (
            .O(N__46302),
            .I(N__46298));
    InMux I__9907 (
            .O(N__46301),
            .I(N__46295));
    LocalMux I__9906 (
            .O(N__46298),
            .I(N__46292));
    LocalMux I__9905 (
            .O(N__46295),
            .I(N__46288));
    Span4Mux_v I__9904 (
            .O(N__46292),
            .I(N__46285));
    InMux I__9903 (
            .O(N__46291),
            .I(N__46282));
    Span12Mux_v I__9902 (
            .O(N__46288),
            .I(N__46279));
    Span4Mux_v I__9901 (
            .O(N__46285),
            .I(N__46276));
    LocalMux I__9900 (
            .O(N__46282),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv12 I__9899 (
            .O(N__46279),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__9898 (
            .O(N__46276),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    InMux I__9897 (
            .O(N__46269),
            .I(N__46266));
    LocalMux I__9896 (
            .O(N__46266),
            .I(N__46263));
    Span4Mux_h I__9895 (
            .O(N__46263),
            .I(N__46260));
    Odrv4 I__9894 (
            .O(N__46260),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__9893 (
            .O(N__46257),
            .I(N__46254));
    LocalMux I__9892 (
            .O(N__46254),
            .I(N__46250));
    InMux I__9891 (
            .O(N__46253),
            .I(N__46247));
    Span4Mux_v I__9890 (
            .O(N__46250),
            .I(N__46242));
    LocalMux I__9889 (
            .O(N__46247),
            .I(N__46242));
    Span4Mux_h I__9888 (
            .O(N__46242),
            .I(N__46239));
    Odrv4 I__9887 (
            .O(N__46239),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    InMux I__9886 (
            .O(N__46236),
            .I(N__46233));
    LocalMux I__9885 (
            .O(N__46233),
            .I(N__46228));
    InMux I__9884 (
            .O(N__46232),
            .I(N__46225));
    CascadeMux I__9883 (
            .O(N__46231),
            .I(N__46222));
    Span4Mux_v I__9882 (
            .O(N__46228),
            .I(N__46219));
    LocalMux I__9881 (
            .O(N__46225),
            .I(N__46216));
    InMux I__9880 (
            .O(N__46222),
            .I(N__46213));
    Span4Mux_h I__9879 (
            .O(N__46219),
            .I(N__46208));
    Span4Mux_v I__9878 (
            .O(N__46216),
            .I(N__46208));
    LocalMux I__9877 (
            .O(N__46213),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__9876 (
            .O(N__46208),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    CascadeMux I__9875 (
            .O(N__46203),
            .I(N__46200));
    InMux I__9874 (
            .O(N__46200),
            .I(N__46191));
    InMux I__9873 (
            .O(N__46199),
            .I(N__46191));
    InMux I__9872 (
            .O(N__46198),
            .I(N__46191));
    LocalMux I__9871 (
            .O(N__46191),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__9870 (
            .O(N__46188),
            .I(N__46185));
    LocalMux I__9869 (
            .O(N__46185),
            .I(N__46182));
    Span4Mux_v I__9868 (
            .O(N__46182),
            .I(N__46179));
    Span4Mux_v I__9867 (
            .O(N__46179),
            .I(N__46176));
    Odrv4 I__9866 (
            .O(N__46176),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ));
    InMux I__9865 (
            .O(N__46173),
            .I(N__46170));
    LocalMux I__9864 (
            .O(N__46170),
            .I(N__46167));
    Span4Mux_h I__9863 (
            .O(N__46167),
            .I(N__46164));
    Odrv4 I__9862 (
            .O(N__46164),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__9861 (
            .O(N__46161),
            .I(N__46157));
    InMux I__9860 (
            .O(N__46160),
            .I(N__46154));
    LocalMux I__9859 (
            .O(N__46157),
            .I(N__46151));
    LocalMux I__9858 (
            .O(N__46154),
            .I(N__46148));
    Span4Mux_h I__9857 (
            .O(N__46151),
            .I(N__46143));
    Span4Mux_h I__9856 (
            .O(N__46148),
            .I(N__46143));
    Odrv4 I__9855 (
            .O(N__46143),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    CascadeMux I__9854 (
            .O(N__46140),
            .I(N__46137));
    InMux I__9853 (
            .O(N__46137),
            .I(N__46134));
    LocalMux I__9852 (
            .O(N__46134),
            .I(N__46131));
    Span4Mux_h I__9851 (
            .O(N__46131),
            .I(N__46128));
    Span4Mux_h I__9850 (
            .O(N__46128),
            .I(N__46123));
    InMux I__9849 (
            .O(N__46127),
            .I(N__46118));
    InMux I__9848 (
            .O(N__46126),
            .I(N__46118));
    Odrv4 I__9847 (
            .O(N__46123),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    LocalMux I__9846 (
            .O(N__46118),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    InMux I__9845 (
            .O(N__46113),
            .I(N__46109));
    InMux I__9844 (
            .O(N__46112),
            .I(N__46105));
    LocalMux I__9843 (
            .O(N__46109),
            .I(N__46102));
    InMux I__9842 (
            .O(N__46108),
            .I(N__46099));
    LocalMux I__9841 (
            .O(N__46105),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    Odrv4 I__9840 (
            .O(N__46102),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    LocalMux I__9839 (
            .O(N__46099),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__9838 (
            .O(N__46092),
            .I(N__46089));
    LocalMux I__9837 (
            .O(N__46089),
            .I(N__46086));
    Span4Mux_v I__9836 (
            .O(N__46086),
            .I(N__46083));
    Odrv4 I__9835 (
            .O(N__46083),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ));
    InMux I__9834 (
            .O(N__46080),
            .I(N__46077));
    LocalMux I__9833 (
            .O(N__46077),
            .I(\ppm_encoder_1.un1_init_pulses_10_0 ));
    CascadeMux I__9832 (
            .O(N__46074),
            .I(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ));
    CascadeMux I__9831 (
            .O(N__46071),
            .I(N__46067));
    InMux I__9830 (
            .O(N__46070),
            .I(N__46064));
    InMux I__9829 (
            .O(N__46067),
            .I(N__46059));
    LocalMux I__9828 (
            .O(N__46064),
            .I(N__46056));
    InMux I__9827 (
            .O(N__46063),
            .I(N__46051));
    InMux I__9826 (
            .O(N__46062),
            .I(N__46051));
    LocalMux I__9825 (
            .O(N__46059),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv4 I__9824 (
            .O(N__46056),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    LocalMux I__9823 (
            .O(N__46051),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    CascadeMux I__9822 (
            .O(N__46044),
            .I(N__46041));
    InMux I__9821 (
            .O(N__46041),
            .I(N__46037));
    InMux I__9820 (
            .O(N__46040),
            .I(N__46033));
    LocalMux I__9819 (
            .O(N__46037),
            .I(N__46030));
    InMux I__9818 (
            .O(N__46036),
            .I(N__46027));
    LocalMux I__9817 (
            .O(N__46033),
            .I(N__46022));
    Span4Mux_h I__9816 (
            .O(N__46030),
            .I(N__46022));
    LocalMux I__9815 (
            .O(N__46027),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    Odrv4 I__9814 (
            .O(N__46022),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    InMux I__9813 (
            .O(N__46017),
            .I(N__46014));
    LocalMux I__9812 (
            .O(N__46014),
            .I(N__46011));
    Span4Mux_h I__9811 (
            .O(N__46011),
            .I(N__46008));
    Odrv4 I__9810 (
            .O(N__46008),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__9809 (
            .O(N__46005),
            .I(N__46001));
    InMux I__9808 (
            .O(N__46004),
            .I(N__45998));
    LocalMux I__9807 (
            .O(N__46001),
            .I(N__45995));
    LocalMux I__9806 (
            .O(N__45998),
            .I(N__45992));
    Span4Mux_v I__9805 (
            .O(N__45995),
            .I(N__45989));
    Odrv12 I__9804 (
            .O(N__45992),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    Odrv4 I__9803 (
            .O(N__45989),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    InMux I__9802 (
            .O(N__45984),
            .I(N__45975));
    InMux I__9801 (
            .O(N__45983),
            .I(N__45975));
    InMux I__9800 (
            .O(N__45982),
            .I(N__45975));
    LocalMux I__9799 (
            .O(N__45975),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    InMux I__9798 (
            .O(N__45972),
            .I(N__45968));
    InMux I__9797 (
            .O(N__45971),
            .I(N__45965));
    LocalMux I__9796 (
            .O(N__45968),
            .I(N__45960));
    LocalMux I__9795 (
            .O(N__45965),
            .I(N__45960));
    Span4Mux_h I__9794 (
            .O(N__45960),
            .I(N__45957));
    Span4Mux_h I__9793 (
            .O(N__45957),
            .I(N__45954));
    Odrv4 I__9792 (
            .O(N__45954),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    InMux I__9791 (
            .O(N__45951),
            .I(N__45948));
    LocalMux I__9790 (
            .O(N__45948),
            .I(N__45945));
    Span4Mux_h I__9789 (
            .O(N__45945),
            .I(N__45942));
    Span4Mux_v I__9788 (
            .O(N__45942),
            .I(N__45939));
    Odrv4 I__9787 (
            .O(N__45939),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ));
    InMux I__9786 (
            .O(N__45936),
            .I(N__45933));
    LocalMux I__9785 (
            .O(N__45933),
            .I(N__45930));
    Span4Mux_h I__9784 (
            .O(N__45930),
            .I(N__45927));
    Odrv4 I__9783 (
            .O(N__45927),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__9782 (
            .O(N__45924),
            .I(N__45920));
    InMux I__9781 (
            .O(N__45923),
            .I(N__45917));
    LocalMux I__9780 (
            .O(N__45920),
            .I(N__45914));
    LocalMux I__9779 (
            .O(N__45917),
            .I(N__45911));
    Span4Mux_v I__9778 (
            .O(N__45914),
            .I(N__45908));
    Span4Mux_h I__9777 (
            .O(N__45911),
            .I(N__45905));
    Odrv4 I__9776 (
            .O(N__45908),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    Odrv4 I__9775 (
            .O(N__45905),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    InMux I__9774 (
            .O(N__45900),
            .I(N__45897));
    LocalMux I__9773 (
            .O(N__45897),
            .I(N__45894));
    Span4Mux_v I__9772 (
            .O(N__45894),
            .I(N__45889));
    InMux I__9771 (
            .O(N__45893),
            .I(N__45884));
    InMux I__9770 (
            .O(N__45892),
            .I(N__45884));
    Odrv4 I__9769 (
            .O(N__45889),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    LocalMux I__9768 (
            .O(N__45884),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    InMux I__9767 (
            .O(N__45879),
            .I(N__45875));
    CascadeMux I__9766 (
            .O(N__45878),
            .I(N__45871));
    LocalMux I__9765 (
            .O(N__45875),
            .I(N__45867));
    InMux I__9764 (
            .O(N__45874),
            .I(N__45862));
    InMux I__9763 (
            .O(N__45871),
            .I(N__45862));
    InMux I__9762 (
            .O(N__45870),
            .I(N__45859));
    Span4Mux_h I__9761 (
            .O(N__45867),
            .I(N__45856));
    LocalMux I__9760 (
            .O(N__45862),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    LocalMux I__9759 (
            .O(N__45859),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    Odrv4 I__9758 (
            .O(N__45856),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    InMux I__9757 (
            .O(N__45849),
            .I(N__45846));
    LocalMux I__9756 (
            .O(N__45846),
            .I(N__45843));
    Span4Mux_h I__9755 (
            .O(N__45843),
            .I(N__45840));
    Span4Mux_v I__9754 (
            .O(N__45840),
            .I(N__45837));
    Odrv4 I__9753 (
            .O(N__45837),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__9752 (
            .O(N__45834),
            .I(N__45830));
    InMux I__9751 (
            .O(N__45833),
            .I(N__45827));
    LocalMux I__9750 (
            .O(N__45830),
            .I(N__45822));
    LocalMux I__9749 (
            .O(N__45827),
            .I(N__45822));
    Span4Mux_v I__9748 (
            .O(N__45822),
            .I(N__45819));
    Odrv4 I__9747 (
            .O(N__45819),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    CascadeMux I__9746 (
            .O(N__45816),
            .I(N__45813));
    InMux I__9745 (
            .O(N__45813),
            .I(N__45810));
    LocalMux I__9744 (
            .O(N__45810),
            .I(N__45807));
    Span4Mux_h I__9743 (
            .O(N__45807),
            .I(N__45804));
    Span4Mux_v I__9742 (
            .O(N__45804),
            .I(N__45801));
    Odrv4 I__9741 (
            .O(N__45801),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ));
    CascadeMux I__9740 (
            .O(N__45798),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_ ));
    InMux I__9739 (
            .O(N__45795),
            .I(N__45792));
    LocalMux I__9738 (
            .O(N__45792),
            .I(N__45789));
    Span4Mux_v I__9737 (
            .O(N__45789),
            .I(N__45786));
    Odrv4 I__9736 (
            .O(N__45786),
            .I(\ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ));
    InMux I__9735 (
            .O(N__45783),
            .I(N__45780));
    LocalMux I__9734 (
            .O(N__45780),
            .I(N__45775));
    InMux I__9733 (
            .O(N__45779),
            .I(N__45772));
    InMux I__9732 (
            .O(N__45778),
            .I(N__45769));
    Span4Mux_v I__9731 (
            .O(N__45775),
            .I(N__45766));
    LocalMux I__9730 (
            .O(N__45772),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__9729 (
            .O(N__45769),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    Odrv4 I__9728 (
            .O(N__45766),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    InMux I__9727 (
            .O(N__45759),
            .I(N__45756));
    LocalMux I__9726 (
            .O(N__45756),
            .I(N__45753));
    Span12Mux_h I__9725 (
            .O(N__45753),
            .I(N__45748));
    InMux I__9724 (
            .O(N__45752),
            .I(N__45745));
    InMux I__9723 (
            .O(N__45751),
            .I(N__45742));
    Odrv12 I__9722 (
            .O(N__45748),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__9721 (
            .O(N__45745),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__9720 (
            .O(N__45742),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    CascadeMux I__9719 (
            .O(N__45735),
            .I(N__45732));
    InMux I__9718 (
            .O(N__45732),
            .I(N__45729));
    LocalMux I__9717 (
            .O(N__45729),
            .I(\pid_side.m26_e_5 ));
    CascadeMux I__9716 (
            .O(N__45726),
            .I(\pid_side.pid_prereg_esr_RNIGJDR1Z0Z_10_cascade_ ));
    InMux I__9715 (
            .O(N__45723),
            .I(N__45720));
    LocalMux I__9714 (
            .O(N__45720),
            .I(\pid_side.m18_s_4 ));
    CascadeMux I__9713 (
            .O(N__45717),
            .I(\pid_side.pid_prereg_esr_RNIQBAH2Z0Z_23_cascade_ ));
    InMux I__9712 (
            .O(N__45714),
            .I(N__45711));
    LocalMux I__9711 (
            .O(N__45711),
            .I(N__45708));
    Odrv4 I__9710 (
            .O(N__45708),
            .I(\pid_side.un1_reset_0_i_sn ));
    CascadeMux I__9709 (
            .O(N__45705),
            .I(\pid_side.i19_mux_cascade_ ));
    InMux I__9708 (
            .O(N__45702),
            .I(N__45691));
    InMux I__9707 (
            .O(N__45701),
            .I(N__45688));
    InMux I__9706 (
            .O(N__45700),
            .I(N__45675));
    InMux I__9705 (
            .O(N__45699),
            .I(N__45675));
    InMux I__9704 (
            .O(N__45698),
            .I(N__45675));
    InMux I__9703 (
            .O(N__45697),
            .I(N__45675));
    InMux I__9702 (
            .O(N__45696),
            .I(N__45675));
    InMux I__9701 (
            .O(N__45695),
            .I(N__45675));
    InMux I__9700 (
            .O(N__45694),
            .I(N__45672));
    LocalMux I__9699 (
            .O(N__45691),
            .I(\pid_side.pid_prereg_esr_RNIEUA9Z0Z_12 ));
    LocalMux I__9698 (
            .O(N__45688),
            .I(\pid_side.pid_prereg_esr_RNIEUA9Z0Z_12 ));
    LocalMux I__9697 (
            .O(N__45675),
            .I(\pid_side.pid_prereg_esr_RNIEUA9Z0Z_12 ));
    LocalMux I__9696 (
            .O(N__45672),
            .I(\pid_side.pid_prereg_esr_RNIEUA9Z0Z_12 ));
    InMux I__9695 (
            .O(N__45663),
            .I(N__45658));
    InMux I__9694 (
            .O(N__45662),
            .I(N__45653));
    InMux I__9693 (
            .O(N__45661),
            .I(N__45653));
    LocalMux I__9692 (
            .O(N__45658),
            .I(\pid_side.N_11_0 ));
    LocalMux I__9691 (
            .O(N__45653),
            .I(\pid_side.N_11_0 ));
    CascadeMux I__9690 (
            .O(N__45648),
            .I(\pid_side.pid_prereg_esr_RNIEUA9Z0Z_12_cascade_ ));
    InMux I__9689 (
            .O(N__45645),
            .I(N__45638));
    InMux I__9688 (
            .O(N__45644),
            .I(N__45638));
    InMux I__9687 (
            .O(N__45643),
            .I(N__45635));
    LocalMux I__9686 (
            .O(N__45638),
            .I(N__45632));
    LocalMux I__9685 (
            .O(N__45635),
            .I(\pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10 ));
    Odrv4 I__9684 (
            .O(N__45632),
            .I(\pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10 ));
    InMux I__9683 (
            .O(N__45627),
            .I(N__45618));
    InMux I__9682 (
            .O(N__45626),
            .I(N__45618));
    InMux I__9681 (
            .O(N__45625),
            .I(N__45618));
    LocalMux I__9680 (
            .O(N__45618),
            .I(N__45615));
    Span4Mux_h I__9679 (
            .O(N__45615),
            .I(N__45610));
    InMux I__9678 (
            .O(N__45614),
            .I(N__45607));
    InMux I__9677 (
            .O(N__45613),
            .I(N__45604));
    Odrv4 I__9676 (
            .O(N__45610),
            .I(\pid_side.N_82_mux ));
    LocalMux I__9675 (
            .O(N__45607),
            .I(\pid_side.N_82_mux ));
    LocalMux I__9674 (
            .O(N__45604),
            .I(\pid_side.N_82_mux ));
    InMux I__9673 (
            .O(N__45597),
            .I(N__45594));
    LocalMux I__9672 (
            .O(N__45594),
            .I(N__45591));
    Span4Mux_h I__9671 (
            .O(N__45591),
            .I(N__45587));
    InMux I__9670 (
            .O(N__45590),
            .I(N__45584));
    Span4Mux_v I__9669 (
            .O(N__45587),
            .I(N__45581));
    LocalMux I__9668 (
            .O(N__45584),
            .I(N__45578));
    Span4Mux_h I__9667 (
            .O(N__45581),
            .I(N__45575));
    Odrv4 I__9666 (
            .O(N__45578),
            .I(side_order_12));
    Odrv4 I__9665 (
            .O(N__45575),
            .I(side_order_12));
    InMux I__9664 (
            .O(N__45570),
            .I(N__45567));
    LocalMux I__9663 (
            .O(N__45567),
            .I(N__45564));
    Odrv4 I__9662 (
            .O(N__45564),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0 ));
    CascadeMux I__9661 (
            .O(N__45561),
            .I(N__45554));
    CascadeMux I__9660 (
            .O(N__45560),
            .I(N__45550));
    InMux I__9659 (
            .O(N__45559),
            .I(N__45547));
    CascadeMux I__9658 (
            .O(N__45558),
            .I(N__45542));
    InMux I__9657 (
            .O(N__45557),
            .I(N__45539));
    InMux I__9656 (
            .O(N__45554),
            .I(N__45536));
    InMux I__9655 (
            .O(N__45553),
            .I(N__45533));
    InMux I__9654 (
            .O(N__45550),
            .I(N__45529));
    LocalMux I__9653 (
            .O(N__45547),
            .I(N__45526));
    InMux I__9652 (
            .O(N__45546),
            .I(N__45523));
    CascadeMux I__9651 (
            .O(N__45545),
            .I(N__45520));
    InMux I__9650 (
            .O(N__45542),
            .I(N__45517));
    LocalMux I__9649 (
            .O(N__45539),
            .I(N__45510));
    LocalMux I__9648 (
            .O(N__45536),
            .I(N__45505));
    LocalMux I__9647 (
            .O(N__45533),
            .I(N__45505));
    CascadeMux I__9646 (
            .O(N__45532),
            .I(N__45500));
    LocalMux I__9645 (
            .O(N__45529),
            .I(N__45493));
    Span4Mux_h I__9644 (
            .O(N__45526),
            .I(N__45493));
    LocalMux I__9643 (
            .O(N__45523),
            .I(N__45493));
    InMux I__9642 (
            .O(N__45520),
            .I(N__45490));
    LocalMux I__9641 (
            .O(N__45517),
            .I(N__45487));
    InMux I__9640 (
            .O(N__45516),
            .I(N__45484));
    CascadeMux I__9639 (
            .O(N__45515),
            .I(N__45480));
    CascadeMux I__9638 (
            .O(N__45514),
            .I(N__45477));
    InMux I__9637 (
            .O(N__45513),
            .I(N__45474));
    Span4Mux_v I__9636 (
            .O(N__45510),
            .I(N__45469));
    Span4Mux_v I__9635 (
            .O(N__45505),
            .I(N__45469));
    InMux I__9634 (
            .O(N__45504),
            .I(N__45464));
    InMux I__9633 (
            .O(N__45503),
            .I(N__45464));
    InMux I__9632 (
            .O(N__45500),
            .I(N__45461));
    Span4Mux_v I__9631 (
            .O(N__45493),
            .I(N__45452));
    LocalMux I__9630 (
            .O(N__45490),
            .I(N__45452));
    Span4Mux_h I__9629 (
            .O(N__45487),
            .I(N__45452));
    LocalMux I__9628 (
            .O(N__45484),
            .I(N__45452));
    InMux I__9627 (
            .O(N__45483),
            .I(N__45449));
    InMux I__9626 (
            .O(N__45480),
            .I(N__45444));
    InMux I__9625 (
            .O(N__45477),
            .I(N__45444));
    LocalMux I__9624 (
            .O(N__45474),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__9623 (
            .O(N__45469),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__9622 (
            .O(N__45464),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__9621 (
            .O(N__45461),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__9620 (
            .O(N__45452),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__9619 (
            .O(N__45449),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__9618 (
            .O(N__45444),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    InMux I__9617 (
            .O(N__45429),
            .I(N__45425));
    InMux I__9616 (
            .O(N__45428),
            .I(N__45422));
    LocalMux I__9615 (
            .O(N__45425),
            .I(N__45419));
    LocalMux I__9614 (
            .O(N__45422),
            .I(N__45416));
    Span12Mux_h I__9613 (
            .O(N__45419),
            .I(N__45413));
    Span4Mux_h I__9612 (
            .O(N__45416),
            .I(N__45410));
    Odrv12 I__9611 (
            .O(N__45413),
            .I(front_order_0));
    Odrv4 I__9610 (
            .O(N__45410),
            .I(front_order_0));
    InMux I__9609 (
            .O(N__45405),
            .I(N__45391));
    CascadeMux I__9608 (
            .O(N__45404),
            .I(N__45382));
    CascadeMux I__9607 (
            .O(N__45403),
            .I(N__45377));
    CascadeMux I__9606 (
            .O(N__45402),
            .I(N__45367));
    CascadeMux I__9605 (
            .O(N__45401),
            .I(N__45364));
    CascadeMux I__9604 (
            .O(N__45400),
            .I(N__45359));
    CascadeMux I__9603 (
            .O(N__45399),
            .I(N__45355));
    CascadeMux I__9602 (
            .O(N__45398),
            .I(N__45351));
    CascadeMux I__9601 (
            .O(N__45397),
            .I(N__45348));
    CascadeMux I__9600 (
            .O(N__45396),
            .I(N__45345));
    CascadeMux I__9599 (
            .O(N__45395),
            .I(N__45337));
    CascadeMux I__9598 (
            .O(N__45394),
            .I(N__45334));
    LocalMux I__9597 (
            .O(N__45391),
            .I(N__45330));
    InMux I__9596 (
            .O(N__45390),
            .I(N__45325));
    InMux I__9595 (
            .O(N__45389),
            .I(N__45325));
    CascadeMux I__9594 (
            .O(N__45388),
            .I(N__45322));
    CascadeMux I__9593 (
            .O(N__45387),
            .I(N__45318));
    CascadeMux I__9592 (
            .O(N__45386),
            .I(N__45315));
    InMux I__9591 (
            .O(N__45385),
            .I(N__45311));
    InMux I__9590 (
            .O(N__45382),
            .I(N__45306));
    InMux I__9589 (
            .O(N__45381),
            .I(N__45306));
    InMux I__9588 (
            .O(N__45380),
            .I(N__45299));
    InMux I__9587 (
            .O(N__45377),
            .I(N__45299));
    InMux I__9586 (
            .O(N__45376),
            .I(N__45299));
    CascadeMux I__9585 (
            .O(N__45375),
            .I(N__45291));
    CascadeMux I__9584 (
            .O(N__45374),
            .I(N__45288));
    CascadeMux I__9583 (
            .O(N__45373),
            .I(N__45285));
    CascadeMux I__9582 (
            .O(N__45372),
            .I(N__45282));
    CascadeMux I__9581 (
            .O(N__45371),
            .I(N__45279));
    CascadeMux I__9580 (
            .O(N__45370),
            .I(N__45276));
    InMux I__9579 (
            .O(N__45367),
            .I(N__45273));
    InMux I__9578 (
            .O(N__45364),
            .I(N__45270));
    InMux I__9577 (
            .O(N__45363),
            .I(N__45267));
    InMux I__9576 (
            .O(N__45362),
            .I(N__45262));
    InMux I__9575 (
            .O(N__45359),
            .I(N__45262));
    InMux I__9574 (
            .O(N__45358),
            .I(N__45257));
    InMux I__9573 (
            .O(N__45355),
            .I(N__45257));
    InMux I__9572 (
            .O(N__45354),
            .I(N__45252));
    InMux I__9571 (
            .O(N__45351),
            .I(N__45252));
    InMux I__9570 (
            .O(N__45348),
            .I(N__45241));
    InMux I__9569 (
            .O(N__45345),
            .I(N__45241));
    InMux I__9568 (
            .O(N__45344),
            .I(N__45241));
    InMux I__9567 (
            .O(N__45343),
            .I(N__45241));
    InMux I__9566 (
            .O(N__45342),
            .I(N__45241));
    InMux I__9565 (
            .O(N__45341),
            .I(N__45230));
    InMux I__9564 (
            .O(N__45340),
            .I(N__45230));
    InMux I__9563 (
            .O(N__45337),
            .I(N__45230));
    InMux I__9562 (
            .O(N__45334),
            .I(N__45230));
    InMux I__9561 (
            .O(N__45333),
            .I(N__45230));
    Span4Mux_v I__9560 (
            .O(N__45330),
            .I(N__45225));
    LocalMux I__9559 (
            .O(N__45325),
            .I(N__45225));
    InMux I__9558 (
            .O(N__45322),
            .I(N__45222));
    InMux I__9557 (
            .O(N__45321),
            .I(N__45215));
    InMux I__9556 (
            .O(N__45318),
            .I(N__45215));
    InMux I__9555 (
            .O(N__45315),
            .I(N__45215));
    CascadeMux I__9554 (
            .O(N__45314),
            .I(N__45212));
    LocalMux I__9553 (
            .O(N__45311),
            .I(N__45209));
    LocalMux I__9552 (
            .O(N__45306),
            .I(N__45204));
    LocalMux I__9551 (
            .O(N__45299),
            .I(N__45204));
    CascadeMux I__9550 (
            .O(N__45298),
            .I(N__45197));
    CascadeMux I__9549 (
            .O(N__45297),
            .I(N__45194));
    CascadeMux I__9548 (
            .O(N__45296),
            .I(N__45191));
    CascadeMux I__9547 (
            .O(N__45295),
            .I(N__45187));
    InMux I__9546 (
            .O(N__45294),
            .I(N__45181));
    InMux I__9545 (
            .O(N__45291),
            .I(N__45181));
    InMux I__9544 (
            .O(N__45288),
            .I(N__45174));
    InMux I__9543 (
            .O(N__45285),
            .I(N__45174));
    InMux I__9542 (
            .O(N__45282),
            .I(N__45174));
    InMux I__9541 (
            .O(N__45279),
            .I(N__45169));
    InMux I__9540 (
            .O(N__45276),
            .I(N__45169));
    LocalMux I__9539 (
            .O(N__45273),
            .I(N__45164));
    LocalMux I__9538 (
            .O(N__45270),
            .I(N__45164));
    LocalMux I__9537 (
            .O(N__45267),
            .I(N__45159));
    LocalMux I__9536 (
            .O(N__45262),
            .I(N__45159));
    LocalMux I__9535 (
            .O(N__45257),
            .I(N__45144));
    LocalMux I__9534 (
            .O(N__45252),
            .I(N__45144));
    LocalMux I__9533 (
            .O(N__45241),
            .I(N__45144));
    LocalMux I__9532 (
            .O(N__45230),
            .I(N__45144));
    Span4Mux_h I__9531 (
            .O(N__45225),
            .I(N__45144));
    LocalMux I__9530 (
            .O(N__45222),
            .I(N__45144));
    LocalMux I__9529 (
            .O(N__45215),
            .I(N__45144));
    InMux I__9528 (
            .O(N__45212),
            .I(N__45141));
    Span4Mux_h I__9527 (
            .O(N__45209),
            .I(N__45136));
    Span4Mux_v I__9526 (
            .O(N__45204),
            .I(N__45136));
    InMux I__9525 (
            .O(N__45203),
            .I(N__45133));
    CascadeMux I__9524 (
            .O(N__45202),
            .I(N__45129));
    CascadeMux I__9523 (
            .O(N__45201),
            .I(N__45126));
    InMux I__9522 (
            .O(N__45200),
            .I(N__45115));
    InMux I__9521 (
            .O(N__45197),
            .I(N__45115));
    InMux I__9520 (
            .O(N__45194),
            .I(N__45115));
    InMux I__9519 (
            .O(N__45191),
            .I(N__45115));
    InMux I__9518 (
            .O(N__45190),
            .I(N__45115));
    InMux I__9517 (
            .O(N__45187),
            .I(N__45110));
    InMux I__9516 (
            .O(N__45186),
            .I(N__45110));
    LocalMux I__9515 (
            .O(N__45181),
            .I(N__45107));
    LocalMux I__9514 (
            .O(N__45174),
            .I(N__45098));
    LocalMux I__9513 (
            .O(N__45169),
            .I(N__45098));
    Span4Mux_v I__9512 (
            .O(N__45164),
            .I(N__45098));
    Span4Mux_v I__9511 (
            .O(N__45159),
            .I(N__45098));
    Span4Mux_v I__9510 (
            .O(N__45144),
            .I(N__45095));
    LocalMux I__9509 (
            .O(N__45141),
            .I(N__45088));
    Span4Mux_h I__9508 (
            .O(N__45136),
            .I(N__45088));
    LocalMux I__9507 (
            .O(N__45133),
            .I(N__45088));
    InMux I__9506 (
            .O(N__45132),
            .I(N__45081));
    InMux I__9505 (
            .O(N__45129),
            .I(N__45081));
    InMux I__9504 (
            .O(N__45126),
            .I(N__45081));
    LocalMux I__9503 (
            .O(N__45115),
            .I(N__45076));
    LocalMux I__9502 (
            .O(N__45110),
            .I(N__45076));
    Span4Mux_v I__9501 (
            .O(N__45107),
            .I(N__45071));
    Span4Mux_v I__9500 (
            .O(N__45098),
            .I(N__45071));
    Span4Mux_v I__9499 (
            .O(N__45095),
            .I(N__45066));
    Span4Mux_v I__9498 (
            .O(N__45088),
            .I(N__45066));
    LocalMux I__9497 (
            .O(N__45081),
            .I(pid_altitude_dv));
    Odrv12 I__9496 (
            .O(N__45076),
            .I(pid_altitude_dv));
    Odrv4 I__9495 (
            .O(N__45071),
            .I(pid_altitude_dv));
    Odrv4 I__9494 (
            .O(N__45066),
            .I(pid_altitude_dv));
    InMux I__9493 (
            .O(N__45057),
            .I(N__45053));
    InMux I__9492 (
            .O(N__45056),
            .I(N__45050));
    LocalMux I__9491 (
            .O(N__45053),
            .I(N__45047));
    LocalMux I__9490 (
            .O(N__45050),
            .I(N__45044));
    Span12Mux_h I__9489 (
            .O(N__45047),
            .I(N__45041));
    Span12Mux_s9_h I__9488 (
            .O(N__45044),
            .I(N__45038));
    Odrv12 I__9487 (
            .O(N__45041),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    Odrv12 I__9486 (
            .O(N__45038),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    InMux I__9485 (
            .O(N__45033),
            .I(N__45029));
    CascadeMux I__9484 (
            .O(N__45032),
            .I(N__45026));
    LocalMux I__9483 (
            .O(N__45029),
            .I(N__45022));
    InMux I__9482 (
            .O(N__45026),
            .I(N__45017));
    InMux I__9481 (
            .O(N__45025),
            .I(N__45017));
    Odrv12 I__9480 (
            .O(N__45022),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__9479 (
            .O(N__45017),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__9478 (
            .O(N__45012),
            .I(N__45008));
    CascadeMux I__9477 (
            .O(N__45011),
            .I(N__45005));
    InMux I__9476 (
            .O(N__45008),
            .I(N__45002));
    InMux I__9475 (
            .O(N__45005),
            .I(N__44999));
    LocalMux I__9474 (
            .O(N__45002),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    LocalMux I__9473 (
            .O(N__44999),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__9472 (
            .O(N__44994),
            .I(N__44991));
    LocalMux I__9471 (
            .O(N__44991),
            .I(\pid_side.m32_1 ));
    InMux I__9470 (
            .O(N__44988),
            .I(N__44985));
    LocalMux I__9469 (
            .O(N__44985),
            .I(N__44981));
    InMux I__9468 (
            .O(N__44984),
            .I(N__44975));
    Span4Mux_h I__9467 (
            .O(N__44981),
            .I(N__44972));
    InMux I__9466 (
            .O(N__44980),
            .I(N__44967));
    InMux I__9465 (
            .O(N__44979),
            .I(N__44961));
    InMux I__9464 (
            .O(N__44978),
            .I(N__44961));
    LocalMux I__9463 (
            .O(N__44975),
            .I(N__44958));
    Span4Mux_h I__9462 (
            .O(N__44972),
            .I(N__44955));
    IoInMux I__9461 (
            .O(N__44971),
            .I(N__44952));
    InMux I__9460 (
            .O(N__44970),
            .I(N__44947));
    LocalMux I__9459 (
            .O(N__44967),
            .I(N__44944));
    InMux I__9458 (
            .O(N__44966),
            .I(N__44941));
    LocalMux I__9457 (
            .O(N__44961),
            .I(N__44938));
    Span4Mux_v I__9456 (
            .O(N__44958),
            .I(N__44935));
    Span4Mux_v I__9455 (
            .O(N__44955),
            .I(N__44932));
    LocalMux I__9454 (
            .O(N__44952),
            .I(N__44929));
    InMux I__9453 (
            .O(N__44951),
            .I(N__44925));
    InMux I__9452 (
            .O(N__44950),
            .I(N__44922));
    LocalMux I__9451 (
            .O(N__44947),
            .I(N__44919));
    Span4Mux_h I__9450 (
            .O(N__44944),
            .I(N__44916));
    LocalMux I__9449 (
            .O(N__44941),
            .I(N__44913));
    Span4Mux_v I__9448 (
            .O(N__44938),
            .I(N__44910));
    Span4Mux_v I__9447 (
            .O(N__44935),
            .I(N__44905));
    Span4Mux_v I__9446 (
            .O(N__44932),
            .I(N__44905));
    Span4Mux_s3_v I__9445 (
            .O(N__44929),
            .I(N__44902));
    InMux I__9444 (
            .O(N__44928),
            .I(N__44899));
    LocalMux I__9443 (
            .O(N__44925),
            .I(N__44896));
    LocalMux I__9442 (
            .O(N__44922),
            .I(N__44891));
    Span4Mux_v I__9441 (
            .O(N__44919),
            .I(N__44891));
    Span4Mux_h I__9440 (
            .O(N__44916),
            .I(N__44888));
    Span4Mux_v I__9439 (
            .O(N__44913),
            .I(N__44881));
    Span4Mux_h I__9438 (
            .O(N__44910),
            .I(N__44881));
    Span4Mux_v I__9437 (
            .O(N__44905),
            .I(N__44881));
    Span4Mux_h I__9436 (
            .O(N__44902),
            .I(N__44878));
    LocalMux I__9435 (
            .O(N__44899),
            .I(reset_system));
    Odrv4 I__9434 (
            .O(N__44896),
            .I(reset_system));
    Odrv4 I__9433 (
            .O(N__44891),
            .I(reset_system));
    Odrv4 I__9432 (
            .O(N__44888),
            .I(reset_system));
    Odrv4 I__9431 (
            .O(N__44881),
            .I(reset_system));
    Odrv4 I__9430 (
            .O(N__44878),
            .I(reset_system));
    CascadeMux I__9429 (
            .O(N__44865),
            .I(\pid_side.m26_e_5_cascade_ ));
    CascadeMux I__9428 (
            .O(N__44862),
            .I(\pid_side.N_11_0_cascade_ ));
    CascadeMux I__9427 (
            .O(N__44859),
            .I(N__44855));
    InMux I__9426 (
            .O(N__44858),
            .I(N__44847));
    InMux I__9425 (
            .O(N__44855),
            .I(N__44847));
    InMux I__9424 (
            .O(N__44854),
            .I(N__44847));
    LocalMux I__9423 (
            .O(N__44847),
            .I(N__44844));
    Span4Mux_v I__9422 (
            .O(N__44844),
            .I(N__44840));
    InMux I__9421 (
            .O(N__44843),
            .I(N__44837));
    Odrv4 I__9420 (
            .O(N__44840),
            .I(\pid_side.pid_prereg_esr_RNILRSP2Z0Z_5 ));
    LocalMux I__9419 (
            .O(N__44837),
            .I(\pid_side.pid_prereg_esr_RNILRSP2Z0Z_5 ));
    InMux I__9418 (
            .O(N__44832),
            .I(N__44823));
    InMux I__9417 (
            .O(N__44831),
            .I(N__44823));
    InMux I__9416 (
            .O(N__44830),
            .I(N__44823));
    LocalMux I__9415 (
            .O(N__44823),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    InMux I__9414 (
            .O(N__44820),
            .I(N__44817));
    LocalMux I__9413 (
            .O(N__44817),
            .I(N__44813));
    InMux I__9412 (
            .O(N__44816),
            .I(N__44810));
    Span4Mux_v I__9411 (
            .O(N__44813),
            .I(N__44807));
    LocalMux I__9410 (
            .O(N__44810),
            .I(N__44804));
    Span4Mux_h I__9409 (
            .O(N__44807),
            .I(N__44801));
    Span4Mux_v I__9408 (
            .O(N__44804),
            .I(N__44798));
    Span4Mux_v I__9407 (
            .O(N__44801),
            .I(N__44795));
    Span4Mux_v I__9406 (
            .O(N__44798),
            .I(N__44792));
    Odrv4 I__9405 (
            .O(N__44795),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    Odrv4 I__9404 (
            .O(N__44792),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    InMux I__9403 (
            .O(N__44787),
            .I(N__44784));
    LocalMux I__9402 (
            .O(N__44784),
            .I(N__44781));
    Odrv4 I__9401 (
            .O(N__44781),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__9400 (
            .O(N__44778),
            .I(N__44775));
    LocalMux I__9399 (
            .O(N__44775),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__9398 (
            .O(N__44772),
            .I(N__44766));
    InMux I__9397 (
            .O(N__44771),
            .I(N__44766));
    LocalMux I__9396 (
            .O(N__44766),
            .I(N__44762));
    InMux I__9395 (
            .O(N__44765),
            .I(N__44759));
    Span4Mux_v I__9394 (
            .O(N__44762),
            .I(N__44756));
    LocalMux I__9393 (
            .O(N__44759),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    Odrv4 I__9392 (
            .O(N__44756),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__9391 (
            .O(N__44751),
            .I(N__44748));
    LocalMux I__9390 (
            .O(N__44748),
            .I(N__44745));
    Span4Mux_h I__9389 (
            .O(N__44745),
            .I(N__44742));
    Odrv4 I__9388 (
            .O(N__44742),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ));
    InMux I__9387 (
            .O(N__44739),
            .I(N__44736));
    LocalMux I__9386 (
            .O(N__44736),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ));
    InMux I__9385 (
            .O(N__44733),
            .I(N__44730));
    LocalMux I__9384 (
            .O(N__44730),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    CascadeMux I__9383 (
            .O(N__44727),
            .I(N__44722));
    InMux I__9382 (
            .O(N__44726),
            .I(N__44717));
    InMux I__9381 (
            .O(N__44725),
            .I(N__44714));
    InMux I__9380 (
            .O(N__44722),
            .I(N__44707));
    InMux I__9379 (
            .O(N__44721),
            .I(N__44707));
    InMux I__9378 (
            .O(N__44720),
            .I(N__44707));
    LocalMux I__9377 (
            .O(N__44717),
            .I(N__44698));
    LocalMux I__9376 (
            .O(N__44714),
            .I(N__44698));
    LocalMux I__9375 (
            .O(N__44707),
            .I(N__44695));
    InMux I__9374 (
            .O(N__44706),
            .I(N__44686));
    InMux I__9373 (
            .O(N__44705),
            .I(N__44686));
    InMux I__9372 (
            .O(N__44704),
            .I(N__44686));
    InMux I__9371 (
            .O(N__44703),
            .I(N__44686));
    Span4Mux_v I__9370 (
            .O(N__44698),
            .I(N__44678));
    Span4Mux_v I__9369 (
            .O(N__44695),
            .I(N__44675));
    LocalMux I__9368 (
            .O(N__44686),
            .I(N__44672));
    InMux I__9367 (
            .O(N__44685),
            .I(N__44661));
    InMux I__9366 (
            .O(N__44684),
            .I(N__44661));
    InMux I__9365 (
            .O(N__44683),
            .I(N__44661));
    InMux I__9364 (
            .O(N__44682),
            .I(N__44661));
    InMux I__9363 (
            .O(N__44681),
            .I(N__44661));
    Span4Mux_v I__9362 (
            .O(N__44678),
            .I(N__44657));
    Sp12to4 I__9361 (
            .O(N__44675),
            .I(N__44650));
    Sp12to4 I__9360 (
            .O(N__44672),
            .I(N__44650));
    LocalMux I__9359 (
            .O(N__44661),
            .I(N__44650));
    InMux I__9358 (
            .O(N__44660),
            .I(N__44647));
    Odrv4 I__9357 (
            .O(N__44657),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv12 I__9356 (
            .O(N__44650),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    LocalMux I__9355 (
            .O(N__44647),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    InMux I__9354 (
            .O(N__44640),
            .I(N__44637));
    LocalMux I__9353 (
            .O(N__44637),
            .I(N__44634));
    Odrv12 I__9352 (
            .O(N__44634),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ));
    InMux I__9351 (
            .O(N__44631),
            .I(N__44628));
    LocalMux I__9350 (
            .O(N__44628),
            .I(N__44625));
    Odrv12 I__9349 (
            .O(N__44625),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ));
    CascadeMux I__9348 (
            .O(N__44622),
            .I(N__44619));
    InMux I__9347 (
            .O(N__44619),
            .I(N__44616));
    LocalMux I__9346 (
            .O(N__44616),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    CEMux I__9345 (
            .O(N__44613),
            .I(N__44609));
    CEMux I__9344 (
            .O(N__44612),
            .I(N__44606));
    LocalMux I__9343 (
            .O(N__44609),
            .I(N__44603));
    LocalMux I__9342 (
            .O(N__44606),
            .I(N__44599));
    Span4Mux_h I__9341 (
            .O(N__44603),
            .I(N__44596));
    CEMux I__9340 (
            .O(N__44602),
            .I(N__44593));
    Span4Mux_v I__9339 (
            .O(N__44599),
            .I(N__44589));
    Span4Mux_v I__9338 (
            .O(N__44596),
            .I(N__44584));
    LocalMux I__9337 (
            .O(N__44593),
            .I(N__44584));
    CEMux I__9336 (
            .O(N__44592),
            .I(N__44581));
    Span4Mux_h I__9335 (
            .O(N__44589),
            .I(N__44577));
    Span4Mux_v I__9334 (
            .O(N__44584),
            .I(N__44572));
    LocalMux I__9333 (
            .O(N__44581),
            .I(N__44572));
    CEMux I__9332 (
            .O(N__44580),
            .I(N__44569));
    Span4Mux_v I__9331 (
            .O(N__44577),
            .I(N__44566));
    Span4Mux_h I__9330 (
            .O(N__44572),
            .I(N__44563));
    LocalMux I__9329 (
            .O(N__44569),
            .I(N__44560));
    Odrv4 I__9328 (
            .O(N__44566),
            .I(\ppm_encoder_1.N_2150_0 ));
    Odrv4 I__9327 (
            .O(N__44563),
            .I(\ppm_encoder_1.N_2150_0 ));
    Odrv12 I__9326 (
            .O(N__44560),
            .I(\ppm_encoder_1.N_2150_0 ));
    InMux I__9325 (
            .O(N__44553),
            .I(N__44548));
    InMux I__9324 (
            .O(N__44552),
            .I(N__44545));
    InMux I__9323 (
            .O(N__44551),
            .I(N__44542));
    LocalMux I__9322 (
            .O(N__44548),
            .I(N__44539));
    LocalMux I__9321 (
            .O(N__44545),
            .I(N__44536));
    LocalMux I__9320 (
            .O(N__44542),
            .I(N__44531));
    Span4Mux_v I__9319 (
            .O(N__44539),
            .I(N__44531));
    Span4Mux_h I__9318 (
            .O(N__44536),
            .I(N__44528));
    Odrv4 I__9317 (
            .O(N__44531),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__9316 (
            .O(N__44528),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__9315 (
            .O(N__44523),
            .I(N__44520));
    LocalMux I__9314 (
            .O(N__44520),
            .I(N__44515));
    InMux I__9313 (
            .O(N__44519),
            .I(N__44512));
    InMux I__9312 (
            .O(N__44518),
            .I(N__44509));
    Span4Mux_h I__9311 (
            .O(N__44515),
            .I(N__44506));
    LocalMux I__9310 (
            .O(N__44512),
            .I(N__44503));
    LocalMux I__9309 (
            .O(N__44509),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv4 I__9308 (
            .O(N__44506),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv4 I__9307 (
            .O(N__44503),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    CascadeMux I__9306 (
            .O(N__44496),
            .I(N__44493));
    InMux I__9305 (
            .O(N__44493),
            .I(N__44488));
    InMux I__9304 (
            .O(N__44492),
            .I(N__44485));
    InMux I__9303 (
            .O(N__44491),
            .I(N__44482));
    LocalMux I__9302 (
            .O(N__44488),
            .I(N__44479));
    LocalMux I__9301 (
            .O(N__44485),
            .I(N__44476));
    LocalMux I__9300 (
            .O(N__44482),
            .I(N__44471));
    Span4Mux_v I__9299 (
            .O(N__44479),
            .I(N__44471));
    Span4Mux_h I__9298 (
            .O(N__44476),
            .I(N__44468));
    Odrv4 I__9297 (
            .O(N__44471),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__9296 (
            .O(N__44468),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__9295 (
            .O(N__44463),
            .I(N__44460));
    LocalMux I__9294 (
            .O(N__44460),
            .I(N__44456));
    InMux I__9293 (
            .O(N__44459),
            .I(N__44452));
    Span4Mux_v I__9292 (
            .O(N__44456),
            .I(N__44449));
    InMux I__9291 (
            .O(N__44455),
            .I(N__44446));
    LocalMux I__9290 (
            .O(N__44452),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    Odrv4 I__9289 (
            .O(N__44449),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__9288 (
            .O(N__44446),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    InMux I__9287 (
            .O(N__44439),
            .I(N__44433));
    InMux I__9286 (
            .O(N__44438),
            .I(N__44433));
    LocalMux I__9285 (
            .O(N__44433),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    InMux I__9284 (
            .O(N__44430),
            .I(N__44427));
    LocalMux I__9283 (
            .O(N__44427),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__9282 (
            .O(N__44424),
            .I(N__44421));
    LocalMux I__9281 (
            .O(N__44421),
            .I(N__44418));
    Span4Mux_v I__9280 (
            .O(N__44418),
            .I(N__44414));
    InMux I__9279 (
            .O(N__44417),
            .I(N__44411));
    Odrv4 I__9278 (
            .O(N__44414),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    LocalMux I__9277 (
            .O(N__44411),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    InMux I__9276 (
            .O(N__44406),
            .I(N__44403));
    LocalMux I__9275 (
            .O(N__44403),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__9274 (
            .O(N__44400),
            .I(N__44397));
    LocalMux I__9273 (
            .O(N__44397),
            .I(N__44394));
    Span4Mux_h I__9272 (
            .O(N__44394),
            .I(N__44390));
    InMux I__9271 (
            .O(N__44393),
            .I(N__44387));
    Odrv4 I__9270 (
            .O(N__44390),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    LocalMux I__9269 (
            .O(N__44387),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    InMux I__9268 (
            .O(N__44382),
            .I(N__44379));
    LocalMux I__9267 (
            .O(N__44379),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    InMux I__9266 (
            .O(N__44376),
            .I(N__44373));
    LocalMux I__9265 (
            .O(N__44373),
            .I(N__44369));
    InMux I__9264 (
            .O(N__44372),
            .I(N__44366));
    Span4Mux_h I__9263 (
            .O(N__44369),
            .I(N__44362));
    LocalMux I__9262 (
            .O(N__44366),
            .I(N__44359));
    InMux I__9261 (
            .O(N__44365),
            .I(N__44356));
    Sp12to4 I__9260 (
            .O(N__44362),
            .I(N__44351));
    Sp12to4 I__9259 (
            .O(N__44359),
            .I(N__44351));
    LocalMux I__9258 (
            .O(N__44356),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv12 I__9257 (
            .O(N__44351),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    InMux I__9256 (
            .O(N__44346),
            .I(N__44343));
    LocalMux I__9255 (
            .O(N__44343),
            .I(N__44340));
    Span4Mux_h I__9254 (
            .O(N__44340),
            .I(N__44337));
    Odrv4 I__9253 (
            .O(N__44337),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ));
    InMux I__9252 (
            .O(N__44334),
            .I(N__44331));
    LocalMux I__9251 (
            .O(N__44331),
            .I(N__44328));
    Odrv4 I__9250 (
            .O(N__44328),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__9249 (
            .O(N__44325),
            .I(N__44322));
    LocalMux I__9248 (
            .O(N__44322),
            .I(N__44318));
    InMux I__9247 (
            .O(N__44321),
            .I(N__44315));
    Span4Mux_h I__9246 (
            .O(N__44318),
            .I(N__44312));
    LocalMux I__9245 (
            .O(N__44315),
            .I(N__44309));
    Span4Mux_h I__9244 (
            .O(N__44312),
            .I(N__44304));
    Span4Mux_h I__9243 (
            .O(N__44309),
            .I(N__44304));
    Odrv4 I__9242 (
            .O(N__44304),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    InMux I__9241 (
            .O(N__44301),
            .I(N__44298));
    LocalMux I__9240 (
            .O(N__44298),
            .I(N__44295));
    Span4Mux_v I__9239 (
            .O(N__44295),
            .I(N__44292));
    Span4Mux_v I__9238 (
            .O(N__44292),
            .I(N__44289));
    Odrv4 I__9237 (
            .O(N__44289),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ));
    InMux I__9236 (
            .O(N__44286),
            .I(N__44283));
    LocalMux I__9235 (
            .O(N__44283),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    InMux I__9234 (
            .O(N__44280),
            .I(N__44277));
    LocalMux I__9233 (
            .O(N__44277),
            .I(N__44273));
    InMux I__9232 (
            .O(N__44276),
            .I(N__44270));
    Odrv12 I__9231 (
            .O(N__44273),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    LocalMux I__9230 (
            .O(N__44270),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    InMux I__9229 (
            .O(N__44265),
            .I(N__44262));
    LocalMux I__9228 (
            .O(N__44262),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__9227 (
            .O(N__44259),
            .I(N__44256));
    LocalMux I__9226 (
            .O(N__44256),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    CascadeMux I__9225 (
            .O(N__44253),
            .I(N__44250));
    InMux I__9224 (
            .O(N__44250),
            .I(N__44247));
    LocalMux I__9223 (
            .O(N__44247),
            .I(N__44244));
    Odrv4 I__9222 (
            .O(N__44244),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__9221 (
            .O(N__44241),
            .I(N__44238));
    LocalMux I__9220 (
            .O(N__44238),
            .I(N__44234));
    InMux I__9219 (
            .O(N__44237),
            .I(N__44231));
    Odrv4 I__9218 (
            .O(N__44234),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    LocalMux I__9217 (
            .O(N__44231),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    InMux I__9216 (
            .O(N__44226),
            .I(N__44220));
    InMux I__9215 (
            .O(N__44225),
            .I(N__44220));
    LocalMux I__9214 (
            .O(N__44220),
            .I(N__44217));
    Span4Mux_v I__9213 (
            .O(N__44217),
            .I(N__44213));
    InMux I__9212 (
            .O(N__44216),
            .I(N__44210));
    Span4Mux_h I__9211 (
            .O(N__44213),
            .I(N__44207));
    LocalMux I__9210 (
            .O(N__44210),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv4 I__9209 (
            .O(N__44207),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    CascadeMux I__9208 (
            .O(N__44202),
            .I(N__44196));
    CascadeMux I__9207 (
            .O(N__44201),
            .I(N__44191));
    CascadeMux I__9206 (
            .O(N__44200),
            .I(N__44186));
    CascadeMux I__9205 (
            .O(N__44199),
            .I(N__44183));
    InMux I__9204 (
            .O(N__44196),
            .I(N__44180));
    InMux I__9203 (
            .O(N__44195),
            .I(N__44177));
    InMux I__9202 (
            .O(N__44194),
            .I(N__44174));
    InMux I__9201 (
            .O(N__44191),
            .I(N__44171));
    CascadeMux I__9200 (
            .O(N__44190),
            .I(N__44167));
    InMux I__9199 (
            .O(N__44189),
            .I(N__44163));
    InMux I__9198 (
            .O(N__44186),
            .I(N__44160));
    InMux I__9197 (
            .O(N__44183),
            .I(N__44156));
    LocalMux I__9196 (
            .O(N__44180),
            .I(N__44153));
    LocalMux I__9195 (
            .O(N__44177),
            .I(N__44148));
    LocalMux I__9194 (
            .O(N__44174),
            .I(N__44148));
    LocalMux I__9193 (
            .O(N__44171),
            .I(N__44145));
    InMux I__9192 (
            .O(N__44170),
            .I(N__44142));
    InMux I__9191 (
            .O(N__44167),
            .I(N__44139));
    InMux I__9190 (
            .O(N__44166),
            .I(N__44136));
    LocalMux I__9189 (
            .O(N__44163),
            .I(N__44133));
    LocalMux I__9188 (
            .O(N__44160),
            .I(N__44130));
    CascadeMux I__9187 (
            .O(N__44159),
            .I(N__44127));
    LocalMux I__9186 (
            .O(N__44156),
            .I(N__44120));
    Span4Mux_v I__9185 (
            .O(N__44153),
            .I(N__44117));
    Span4Mux_v I__9184 (
            .O(N__44148),
            .I(N__44108));
    Span4Mux_h I__9183 (
            .O(N__44145),
            .I(N__44108));
    LocalMux I__9182 (
            .O(N__44142),
            .I(N__44108));
    LocalMux I__9181 (
            .O(N__44139),
            .I(N__44108));
    LocalMux I__9180 (
            .O(N__44136),
            .I(N__44101));
    Span4Mux_h I__9179 (
            .O(N__44133),
            .I(N__44101));
    Span4Mux_h I__9178 (
            .O(N__44130),
            .I(N__44101));
    InMux I__9177 (
            .O(N__44127),
            .I(N__44096));
    InMux I__9176 (
            .O(N__44126),
            .I(N__44096));
    InMux I__9175 (
            .O(N__44125),
            .I(N__44093));
    InMux I__9174 (
            .O(N__44124),
            .I(N__44088));
    InMux I__9173 (
            .O(N__44123),
            .I(N__44088));
    Odrv4 I__9172 (
            .O(N__44120),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__9171 (
            .O(N__44117),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__9170 (
            .O(N__44108),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__9169 (
            .O(N__44101),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__9168 (
            .O(N__44096),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__9167 (
            .O(N__44093),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__9166 (
            .O(N__44088),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    CascadeMux I__9165 (
            .O(N__44073),
            .I(N__44066));
    CascadeMux I__9164 (
            .O(N__44072),
            .I(N__44063));
    CascadeMux I__9163 (
            .O(N__44071),
            .I(N__44060));
    CascadeMux I__9162 (
            .O(N__44070),
            .I(N__44055));
    InMux I__9161 (
            .O(N__44069),
            .I(N__44050));
    InMux I__9160 (
            .O(N__44066),
            .I(N__44045));
    InMux I__9159 (
            .O(N__44063),
            .I(N__44042));
    InMux I__9158 (
            .O(N__44060),
            .I(N__44039));
    InMux I__9157 (
            .O(N__44059),
            .I(N__44034));
    InMux I__9156 (
            .O(N__44058),
            .I(N__44034));
    InMux I__9155 (
            .O(N__44055),
            .I(N__44031));
    InMux I__9154 (
            .O(N__44054),
            .I(N__44028));
    InMux I__9153 (
            .O(N__44053),
            .I(N__44025));
    LocalMux I__9152 (
            .O(N__44050),
            .I(N__44022));
    InMux I__9151 (
            .O(N__44049),
            .I(N__44015));
    InMux I__9150 (
            .O(N__44048),
            .I(N__44015));
    LocalMux I__9149 (
            .O(N__44045),
            .I(N__44012));
    LocalMux I__9148 (
            .O(N__44042),
            .I(N__44005));
    LocalMux I__9147 (
            .O(N__44039),
            .I(N__44005));
    LocalMux I__9146 (
            .O(N__44034),
            .I(N__44005));
    LocalMux I__9145 (
            .O(N__44031),
            .I(N__43998));
    LocalMux I__9144 (
            .O(N__44028),
            .I(N__43998));
    LocalMux I__9143 (
            .O(N__44025),
            .I(N__43998));
    Span4Mux_v I__9142 (
            .O(N__44022),
            .I(N__43995));
    InMux I__9141 (
            .O(N__44021),
            .I(N__43992));
    InMux I__9140 (
            .O(N__44020),
            .I(N__43989));
    LocalMux I__9139 (
            .O(N__44015),
            .I(N__43980));
    Span4Mux_h I__9138 (
            .O(N__44012),
            .I(N__43980));
    Span4Mux_v I__9137 (
            .O(N__44005),
            .I(N__43980));
    Span4Mux_v I__9136 (
            .O(N__43998),
            .I(N__43980));
    Odrv4 I__9135 (
            .O(N__43995),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__9134 (
            .O(N__43992),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__9133 (
            .O(N__43989),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__9132 (
            .O(N__43980),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    CascadeMux I__9131 (
            .O(N__43971),
            .I(\ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ));
    CascadeMux I__9130 (
            .O(N__43968),
            .I(N__43965));
    InMux I__9129 (
            .O(N__43965),
            .I(N__43962));
    LocalMux I__9128 (
            .O(N__43962),
            .I(\ppm_encoder_1.elevator_RNIT3R05Z0Z_3 ));
    InMux I__9127 (
            .O(N__43959),
            .I(N__43956));
    LocalMux I__9126 (
            .O(N__43956),
            .I(\ppm_encoder_1.N_289 ));
    CascadeMux I__9125 (
            .O(N__43953),
            .I(N__43949));
    InMux I__9124 (
            .O(N__43952),
            .I(N__43946));
    InMux I__9123 (
            .O(N__43949),
            .I(N__43943));
    LocalMux I__9122 (
            .O(N__43946),
            .I(N__43940));
    LocalMux I__9121 (
            .O(N__43943),
            .I(N__43937));
    Span4Mux_h I__9120 (
            .O(N__43940),
            .I(N__43934));
    Odrv4 I__9119 (
            .O(N__43937),
            .I(side_order_3));
    Odrv4 I__9118 (
            .O(N__43934),
            .I(side_order_3));
    InMux I__9117 (
            .O(N__43929),
            .I(N__43926));
    LocalMux I__9116 (
            .O(N__43926),
            .I(N__43923));
    Span12Mux_v I__9115 (
            .O(N__43923),
            .I(N__43920));
    Odrv12 I__9114 (
            .O(N__43920),
            .I(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ));
    InMux I__9113 (
            .O(N__43917),
            .I(N__43912));
    InMux I__9112 (
            .O(N__43916),
            .I(N__43907));
    InMux I__9111 (
            .O(N__43915),
            .I(N__43907));
    LocalMux I__9110 (
            .O(N__43912),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    LocalMux I__9109 (
            .O(N__43907),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    InMux I__9108 (
            .O(N__43902),
            .I(N__43899));
    LocalMux I__9107 (
            .O(N__43899),
            .I(N__43896));
    Span4Mux_h I__9106 (
            .O(N__43896),
            .I(N__43893));
    Odrv4 I__9105 (
            .O(N__43893),
            .I(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ));
    InMux I__9104 (
            .O(N__43890),
            .I(N__43887));
    LocalMux I__9103 (
            .O(N__43887),
            .I(N__43883));
    InMux I__9102 (
            .O(N__43886),
            .I(N__43880));
    Span4Mux_h I__9101 (
            .O(N__43883),
            .I(N__43875));
    LocalMux I__9100 (
            .O(N__43880),
            .I(N__43875));
    Span4Mux_h I__9099 (
            .O(N__43875),
            .I(N__43872));
    Span4Mux_v I__9098 (
            .O(N__43872),
            .I(N__43869));
    Odrv4 I__9097 (
            .O(N__43869),
            .I(front_order_3));
    InMux I__9096 (
            .O(N__43866),
            .I(N__43857));
    InMux I__9095 (
            .O(N__43865),
            .I(N__43857));
    InMux I__9094 (
            .O(N__43864),
            .I(N__43857));
    LocalMux I__9093 (
            .O(N__43857),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    CascadeMux I__9092 (
            .O(N__43854),
            .I(N__43851));
    InMux I__9091 (
            .O(N__43851),
            .I(N__43848));
    LocalMux I__9090 (
            .O(N__43848),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__9089 (
            .O(N__43845),
            .I(N__43842));
    LocalMux I__9088 (
            .O(N__43842),
            .I(N__43838));
    InMux I__9087 (
            .O(N__43841),
            .I(N__43835));
    Span4Mux_h I__9086 (
            .O(N__43838),
            .I(N__43832));
    LocalMux I__9085 (
            .O(N__43835),
            .I(N__43829));
    Odrv4 I__9084 (
            .O(N__43832),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    Odrv4 I__9083 (
            .O(N__43829),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    InMux I__9082 (
            .O(N__43824),
            .I(N__43821));
    LocalMux I__9081 (
            .O(N__43821),
            .I(N__43818));
    Span4Mux_v I__9080 (
            .O(N__43818),
            .I(N__43815));
    Span4Mux_v I__9079 (
            .O(N__43815),
            .I(N__43812));
    Odrv4 I__9078 (
            .O(N__43812),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    CascadeMux I__9077 (
            .O(N__43809),
            .I(N__43806));
    InMux I__9076 (
            .O(N__43806),
            .I(N__43803));
    LocalMux I__9075 (
            .O(N__43803),
            .I(N__43800));
    Span4Mux_h I__9074 (
            .O(N__43800),
            .I(N__43797));
    Odrv4 I__9073 (
            .O(N__43797),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ));
    InMux I__9072 (
            .O(N__43794),
            .I(N__43789));
    InMux I__9071 (
            .O(N__43793),
            .I(N__43786));
    CascadeMux I__9070 (
            .O(N__43792),
            .I(N__43783));
    LocalMux I__9069 (
            .O(N__43789),
            .I(N__43780));
    LocalMux I__9068 (
            .O(N__43786),
            .I(N__43777));
    InMux I__9067 (
            .O(N__43783),
            .I(N__43774));
    Span4Mux_v I__9066 (
            .O(N__43780),
            .I(N__43771));
    Span4Mux_v I__9065 (
            .O(N__43777),
            .I(N__43768));
    LocalMux I__9064 (
            .O(N__43774),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    Odrv4 I__9063 (
            .O(N__43771),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    Odrv4 I__9062 (
            .O(N__43768),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    CascadeMux I__9061 (
            .O(N__43761),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ));
    CascadeMux I__9060 (
            .O(N__43758),
            .I(N__43755));
    InMux I__9059 (
            .O(N__43755),
            .I(N__43752));
    LocalMux I__9058 (
            .O(N__43752),
            .I(N__43749));
    Odrv4 I__9057 (
            .O(N__43749),
            .I(\ppm_encoder_1.elevator_RNIPVQ05Z0Z_2 ));
    InMux I__9056 (
            .O(N__43746),
            .I(N__43740));
    InMux I__9055 (
            .O(N__43745),
            .I(N__43733));
    InMux I__9054 (
            .O(N__43744),
            .I(N__43733));
    InMux I__9053 (
            .O(N__43743),
            .I(N__43733));
    LocalMux I__9052 (
            .O(N__43740),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__9051 (
            .O(N__43733),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    CascadeMux I__9050 (
            .O(N__43728),
            .I(N__43725));
    InMux I__9049 (
            .O(N__43725),
            .I(N__43719));
    InMux I__9048 (
            .O(N__43724),
            .I(N__43716));
    InMux I__9047 (
            .O(N__43723),
            .I(N__43711));
    InMux I__9046 (
            .O(N__43722),
            .I(N__43711));
    LocalMux I__9045 (
            .O(N__43719),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__9044 (
            .O(N__43716),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__9043 (
            .O(N__43711),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    CascadeMux I__9042 (
            .O(N__43704),
            .I(N__43700));
    InMux I__9041 (
            .O(N__43703),
            .I(N__43696));
    InMux I__9040 (
            .O(N__43700),
            .I(N__43693));
    InMux I__9039 (
            .O(N__43699),
            .I(N__43688));
    LocalMux I__9038 (
            .O(N__43696),
            .I(N__43685));
    LocalMux I__9037 (
            .O(N__43693),
            .I(N__43682));
    InMux I__9036 (
            .O(N__43692),
            .I(N__43677));
    InMux I__9035 (
            .O(N__43691),
            .I(N__43677));
    LocalMux I__9034 (
            .O(N__43688),
            .I(\ppm_encoder_1.N_221 ));
    Odrv4 I__9033 (
            .O(N__43685),
            .I(\ppm_encoder_1.N_221 ));
    Odrv4 I__9032 (
            .O(N__43682),
            .I(\ppm_encoder_1.N_221 ));
    LocalMux I__9031 (
            .O(N__43677),
            .I(\ppm_encoder_1.N_221 ));
    InMux I__9030 (
            .O(N__43668),
            .I(N__43664));
    InMux I__9029 (
            .O(N__43667),
            .I(N__43661));
    LocalMux I__9028 (
            .O(N__43664),
            .I(N__43655));
    LocalMux I__9027 (
            .O(N__43661),
            .I(N__43655));
    InMux I__9026 (
            .O(N__43660),
            .I(N__43652));
    Span4Mux_v I__9025 (
            .O(N__43655),
            .I(N__43649));
    LocalMux I__9024 (
            .O(N__43652),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    Odrv4 I__9023 (
            .O(N__43649),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    CascadeMux I__9022 (
            .O(N__43644),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ));
    CascadeMux I__9021 (
            .O(N__43641),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ));
    InMux I__9020 (
            .O(N__43638),
            .I(N__43635));
    LocalMux I__9019 (
            .O(N__43635),
            .I(N__43632));
    Odrv4 I__9018 (
            .O(N__43632),
            .I(\ppm_encoder_1.elevator_RNIHNQ05Z0Z_0 ));
    InMux I__9017 (
            .O(N__43629),
            .I(N__43625));
    InMux I__9016 (
            .O(N__43628),
            .I(N__43622));
    LocalMux I__9015 (
            .O(N__43625),
            .I(N__43619));
    LocalMux I__9014 (
            .O(N__43622),
            .I(N__43615));
    Span4Mux_h I__9013 (
            .O(N__43619),
            .I(N__43612));
    InMux I__9012 (
            .O(N__43618),
            .I(N__43609));
    Span4Mux_v I__9011 (
            .O(N__43615),
            .I(N__43605));
    Span4Mux_v I__9010 (
            .O(N__43612),
            .I(N__43600));
    LocalMux I__9009 (
            .O(N__43609),
            .I(N__43600));
    InMux I__9008 (
            .O(N__43608),
            .I(N__43597));
    Odrv4 I__9007 (
            .O(N__43605),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv4 I__9006 (
            .O(N__43600),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    LocalMux I__9005 (
            .O(N__43597),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    InMux I__9004 (
            .O(N__43590),
            .I(N__43587));
    LocalMux I__9003 (
            .O(N__43587),
            .I(N__43583));
    InMux I__9002 (
            .O(N__43586),
            .I(N__43580));
    Sp12to4 I__9001 (
            .O(N__43583),
            .I(N__43575));
    LocalMux I__9000 (
            .O(N__43580),
            .I(N__43575));
    Span12Mux_v I__8999 (
            .O(N__43575),
            .I(N__43570));
    InMux I__8998 (
            .O(N__43574),
            .I(N__43565));
    InMux I__8997 (
            .O(N__43573),
            .I(N__43565));
    Odrv12 I__8996 (
            .O(N__43570),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__8995 (
            .O(N__43565),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    CascadeMux I__8994 (
            .O(N__43560),
            .I(N__43557));
    InMux I__8993 (
            .O(N__43557),
            .I(N__43551));
    InMux I__8992 (
            .O(N__43556),
            .I(N__43551));
    LocalMux I__8991 (
            .O(N__43551),
            .I(N__43548));
    Span4Mux_v I__8990 (
            .O(N__43548),
            .I(N__43545));
    Span4Mux_v I__8989 (
            .O(N__43545),
            .I(N__43542));
    Odrv4 I__8988 (
            .O(N__43542),
            .I(\ppm_encoder_1.N_232 ));
    CascadeMux I__8987 (
            .O(N__43539),
            .I(N__43533));
    InMux I__8986 (
            .O(N__43538),
            .I(N__43530));
    InMux I__8985 (
            .O(N__43537),
            .I(N__43527));
    InMux I__8984 (
            .O(N__43536),
            .I(N__43524));
    InMux I__8983 (
            .O(N__43533),
            .I(N__43521));
    LocalMux I__8982 (
            .O(N__43530),
            .I(N__43518));
    LocalMux I__8981 (
            .O(N__43527),
            .I(N__43512));
    LocalMux I__8980 (
            .O(N__43524),
            .I(N__43512));
    LocalMux I__8979 (
            .O(N__43521),
            .I(N__43505));
    Span4Mux_h I__8978 (
            .O(N__43518),
            .I(N__43505));
    InMux I__8977 (
            .O(N__43517),
            .I(N__43502));
    Sp12to4 I__8976 (
            .O(N__43512),
            .I(N__43499));
    InMux I__8975 (
            .O(N__43511),
            .I(N__43494));
    InMux I__8974 (
            .O(N__43510),
            .I(N__43494));
    Odrv4 I__8973 (
            .O(N__43505),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__8972 (
            .O(N__43502),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv12 I__8971 (
            .O(N__43499),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__8970 (
            .O(N__43494),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    InMux I__8969 (
            .O(N__43485),
            .I(N__43476));
    InMux I__8968 (
            .O(N__43484),
            .I(N__43473));
    InMux I__8967 (
            .O(N__43483),
            .I(N__43468));
    InMux I__8966 (
            .O(N__43482),
            .I(N__43468));
    InMux I__8965 (
            .O(N__43481),
            .I(N__43463));
    InMux I__8964 (
            .O(N__43480),
            .I(N__43463));
    InMux I__8963 (
            .O(N__43479),
            .I(N__43460));
    LocalMux I__8962 (
            .O(N__43476),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__8961 (
            .O(N__43473),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__8960 (
            .O(N__43468),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__8959 (
            .O(N__43463),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__8958 (
            .O(N__43460),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    CascadeMux I__8957 (
            .O(N__43449),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_ ));
    CascadeMux I__8956 (
            .O(N__43446),
            .I(N__43442));
    CascadeMux I__8955 (
            .O(N__43445),
            .I(N__43439));
    InMux I__8954 (
            .O(N__43442),
            .I(N__43432));
    InMux I__8953 (
            .O(N__43439),
            .I(N__43429));
    InMux I__8952 (
            .O(N__43438),
            .I(N__43424));
    InMux I__8951 (
            .O(N__43437),
            .I(N__43424));
    InMux I__8950 (
            .O(N__43436),
            .I(N__43419));
    InMux I__8949 (
            .O(N__43435),
            .I(N__43419));
    LocalMux I__8948 (
            .O(N__43432),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__8947 (
            .O(N__43429),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__8946 (
            .O(N__43424),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__8945 (
            .O(N__43419),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    CascadeMux I__8944 (
            .O(N__43410),
            .I(N__43405));
    InMux I__8943 (
            .O(N__43409),
            .I(N__43402));
    InMux I__8942 (
            .O(N__43408),
            .I(N__43399));
    InMux I__8941 (
            .O(N__43405),
            .I(N__43396));
    LocalMux I__8940 (
            .O(N__43402),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__8939 (
            .O(N__43399),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__8938 (
            .O(N__43396),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    InMux I__8937 (
            .O(N__43389),
            .I(N__43384));
    InMux I__8936 (
            .O(N__43388),
            .I(N__43379));
    InMux I__8935 (
            .O(N__43387),
            .I(N__43376));
    LocalMux I__8934 (
            .O(N__43384),
            .I(N__43373));
    InMux I__8933 (
            .O(N__43383),
            .I(N__43368));
    InMux I__8932 (
            .O(N__43382),
            .I(N__43368));
    LocalMux I__8931 (
            .O(N__43379),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__8930 (
            .O(N__43376),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__8929 (
            .O(N__43373),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__8928 (
            .O(N__43368),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    CascadeMux I__8927 (
            .O(N__43359),
            .I(N__43352));
    InMux I__8926 (
            .O(N__43358),
            .I(N__43347));
    InMux I__8925 (
            .O(N__43357),
            .I(N__43344));
    InMux I__8924 (
            .O(N__43356),
            .I(N__43337));
    InMux I__8923 (
            .O(N__43355),
            .I(N__43337));
    InMux I__8922 (
            .O(N__43352),
            .I(N__43337));
    InMux I__8921 (
            .O(N__43351),
            .I(N__43332));
    InMux I__8920 (
            .O(N__43350),
            .I(N__43332));
    LocalMux I__8919 (
            .O(N__43347),
            .I(N__43327));
    LocalMux I__8918 (
            .O(N__43344),
            .I(N__43327));
    LocalMux I__8917 (
            .O(N__43337),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__8916 (
            .O(N__43332),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__8915 (
            .O(N__43327),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    CascadeMux I__8914 (
            .O(N__43320),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ));
    CascadeMux I__8913 (
            .O(N__43317),
            .I(N__43313));
    InMux I__8912 (
            .O(N__43316),
            .I(N__43309));
    InMux I__8911 (
            .O(N__43313),
            .I(N__43306));
    InMux I__8910 (
            .O(N__43312),
            .I(N__43303));
    LocalMux I__8909 (
            .O(N__43309),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    LocalMux I__8908 (
            .O(N__43306),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    LocalMux I__8907 (
            .O(N__43303),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    CascadeMux I__8906 (
            .O(N__43296),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ));
    InMux I__8905 (
            .O(N__43293),
            .I(N__43290));
    LocalMux I__8904 (
            .O(N__43290),
            .I(N__43286));
    InMux I__8903 (
            .O(N__43289),
            .I(N__43283));
    Span12Mux_h I__8902 (
            .O(N__43286),
            .I(N__43280));
    LocalMux I__8901 (
            .O(N__43283),
            .I(side_order_0));
    Odrv12 I__8900 (
            .O(N__43280),
            .I(side_order_0));
    InMux I__8899 (
            .O(N__43275),
            .I(N__43271));
    InMux I__8898 (
            .O(N__43274),
            .I(N__43268));
    LocalMux I__8897 (
            .O(N__43271),
            .I(N__43265));
    LocalMux I__8896 (
            .O(N__43268),
            .I(N__43262));
    Span4Mux_v I__8895 (
            .O(N__43265),
            .I(N__43259));
    Span4Mux_v I__8894 (
            .O(N__43262),
            .I(N__43256));
    Span4Mux_h I__8893 (
            .O(N__43259),
            .I(N__43253));
    Odrv4 I__8892 (
            .O(N__43256),
            .I(side_order_5));
    Odrv4 I__8891 (
            .O(N__43253),
            .I(side_order_5));
    InMux I__8890 (
            .O(N__43248),
            .I(N__43244));
    InMux I__8889 (
            .O(N__43247),
            .I(N__43241));
    LocalMux I__8888 (
            .O(N__43244),
            .I(N__43236));
    LocalMux I__8887 (
            .O(N__43241),
            .I(N__43236));
    Span4Mux_v I__8886 (
            .O(N__43236),
            .I(N__43233));
    Span4Mux_h I__8885 (
            .O(N__43233),
            .I(N__43230));
    Odrv4 I__8884 (
            .O(N__43230),
            .I(side_order_4));
    InMux I__8883 (
            .O(N__43227),
            .I(N__43224));
    LocalMux I__8882 (
            .O(N__43224),
            .I(N__43220));
    InMux I__8881 (
            .O(N__43223),
            .I(N__43217));
    Span4Mux_v I__8880 (
            .O(N__43220),
            .I(N__43211));
    LocalMux I__8879 (
            .O(N__43217),
            .I(N__43211));
    InMux I__8878 (
            .O(N__43216),
            .I(N__43208));
    Span4Mux_h I__8877 (
            .O(N__43211),
            .I(N__43205));
    LocalMux I__8876 (
            .O(N__43208),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv4 I__8875 (
            .O(N__43205),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    InMux I__8874 (
            .O(N__43200),
            .I(N__43196));
    CascadeMux I__8873 (
            .O(N__43199),
            .I(N__43193));
    LocalMux I__8872 (
            .O(N__43196),
            .I(N__43190));
    InMux I__8871 (
            .O(N__43193),
            .I(N__43186));
    Span4Mux_v I__8870 (
            .O(N__43190),
            .I(N__43183));
    InMux I__8869 (
            .O(N__43189),
            .I(N__43180));
    LocalMux I__8868 (
            .O(N__43186),
            .I(N__43173));
    Span4Mux_h I__8867 (
            .O(N__43183),
            .I(N__43173));
    LocalMux I__8866 (
            .O(N__43180),
            .I(N__43173));
    Odrv4 I__8865 (
            .O(N__43173),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    CascadeMux I__8864 (
            .O(N__43170),
            .I(N__43167));
    InMux I__8863 (
            .O(N__43167),
            .I(N__43164));
    LocalMux I__8862 (
            .O(N__43164),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    CascadeMux I__8861 (
            .O(N__43161),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ));
    InMux I__8860 (
            .O(N__43158),
            .I(N__43153));
    InMux I__8859 (
            .O(N__43157),
            .I(N__43148));
    InMux I__8858 (
            .O(N__43156),
            .I(N__43148));
    LocalMux I__8857 (
            .O(N__43153),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__8856 (
            .O(N__43148),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    InMux I__8855 (
            .O(N__43143),
            .I(N__43138));
    InMux I__8854 (
            .O(N__43142),
            .I(N__43133));
    InMux I__8853 (
            .O(N__43141),
            .I(N__43133));
    LocalMux I__8852 (
            .O(N__43138),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__8851 (
            .O(N__43133),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    CascadeMux I__8850 (
            .O(N__43128),
            .I(N__43125));
    InMux I__8849 (
            .O(N__43125),
            .I(N__43121));
    InMux I__8848 (
            .O(N__43124),
            .I(N__43117));
    LocalMux I__8847 (
            .O(N__43121),
            .I(N__43114));
    InMux I__8846 (
            .O(N__43120),
            .I(N__43111));
    LocalMux I__8845 (
            .O(N__43117),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__8844 (
            .O(N__43114),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__8843 (
            .O(N__43111),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    InMux I__8842 (
            .O(N__43104),
            .I(N__43099));
    InMux I__8841 (
            .O(N__43103),
            .I(N__43096));
    InMux I__8840 (
            .O(N__43102),
            .I(N__43093));
    LocalMux I__8839 (
            .O(N__43099),
            .I(N__43090));
    LocalMux I__8838 (
            .O(N__43096),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__8837 (
            .O(N__43093),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    Odrv4 I__8836 (
            .O(N__43090),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    CascadeMux I__8835 (
            .O(N__43083),
            .I(N__43079));
    InMux I__8834 (
            .O(N__43082),
            .I(N__43074));
    InMux I__8833 (
            .O(N__43079),
            .I(N__43074));
    LocalMux I__8832 (
            .O(N__43074),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    InMux I__8831 (
            .O(N__43071),
            .I(N__43068));
    LocalMux I__8830 (
            .O(N__43068),
            .I(N__43065));
    Span4Mux_v I__8829 (
            .O(N__43065),
            .I(N__43062));
    Odrv4 I__8828 (
            .O(N__43062),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    CascadeMux I__8827 (
            .O(N__43059),
            .I(N__43056));
    InMux I__8826 (
            .O(N__43056),
            .I(N__43050));
    InMux I__8825 (
            .O(N__43055),
            .I(N__43050));
    LocalMux I__8824 (
            .O(N__43050),
            .I(N__43047));
    Odrv4 I__8823 (
            .O(N__43047),
            .I(\pid_front.error_d_reg_prevZ0Z_20 ));
    InMux I__8822 (
            .O(N__43044),
            .I(N__43040));
    InMux I__8821 (
            .O(N__43043),
            .I(N__43037));
    LocalMux I__8820 (
            .O(N__43040),
            .I(N__43034));
    LocalMux I__8819 (
            .O(N__43037),
            .I(N__43028));
    Span4Mux_v I__8818 (
            .O(N__43034),
            .I(N__43028));
    CascadeMux I__8817 (
            .O(N__43033),
            .I(N__43025));
    Span4Mux_v I__8816 (
            .O(N__43028),
            .I(N__43022));
    InMux I__8815 (
            .O(N__43025),
            .I(N__43019));
    Span4Mux_h I__8814 (
            .O(N__43022),
            .I(N__43016));
    LocalMux I__8813 (
            .O(N__43019),
            .I(side_order_10));
    Odrv4 I__8812 (
            .O(N__43016),
            .I(side_order_10));
    InMux I__8811 (
            .O(N__43011),
            .I(N__43007));
    CascadeMux I__8810 (
            .O(N__43010),
            .I(N__43003));
    LocalMux I__8809 (
            .O(N__43007),
            .I(N__43000));
    CascadeMux I__8808 (
            .O(N__43006),
            .I(N__42997));
    InMux I__8807 (
            .O(N__43003),
            .I(N__42994));
    Span4Mux_v I__8806 (
            .O(N__43000),
            .I(N__42991));
    InMux I__8805 (
            .O(N__42997),
            .I(N__42988));
    LocalMux I__8804 (
            .O(N__42994),
            .I(N__42983));
    Span4Mux_h I__8803 (
            .O(N__42991),
            .I(N__42983));
    LocalMux I__8802 (
            .O(N__42988),
            .I(N__42978));
    Span4Mux_v I__8801 (
            .O(N__42983),
            .I(N__42978));
    Odrv4 I__8800 (
            .O(N__42978),
            .I(side_order_11));
    CascadeMux I__8799 (
            .O(N__42975),
            .I(N__42971));
    CascadeMux I__8798 (
            .O(N__42974),
            .I(N__42968));
    InMux I__8797 (
            .O(N__42971),
            .I(N__42965));
    InMux I__8796 (
            .O(N__42968),
            .I(N__42962));
    LocalMux I__8795 (
            .O(N__42965),
            .I(N__42958));
    LocalMux I__8794 (
            .O(N__42962),
            .I(N__42955));
    CascadeMux I__8793 (
            .O(N__42961),
            .I(N__42952));
    Span4Mux_v I__8792 (
            .O(N__42958),
            .I(N__42949));
    Span4Mux_v I__8791 (
            .O(N__42955),
            .I(N__42946));
    InMux I__8790 (
            .O(N__42952),
            .I(N__42943));
    Span4Mux_v I__8789 (
            .O(N__42949),
            .I(N__42940));
    Span4Mux_h I__8788 (
            .O(N__42946),
            .I(N__42937));
    LocalMux I__8787 (
            .O(N__42943),
            .I(side_order_6));
    Odrv4 I__8786 (
            .O(N__42940),
            .I(side_order_6));
    Odrv4 I__8785 (
            .O(N__42937),
            .I(side_order_6));
    CascadeMux I__8784 (
            .O(N__42930),
            .I(N__42926));
    CascadeMux I__8783 (
            .O(N__42929),
            .I(N__42923));
    InMux I__8782 (
            .O(N__42926),
            .I(N__42920));
    InMux I__8781 (
            .O(N__42923),
            .I(N__42917));
    LocalMux I__8780 (
            .O(N__42920),
            .I(N__42913));
    LocalMux I__8779 (
            .O(N__42917),
            .I(N__42910));
    CascadeMux I__8778 (
            .O(N__42916),
            .I(N__42907));
    Span4Mux_h I__8777 (
            .O(N__42913),
            .I(N__42904));
    Span4Mux_v I__8776 (
            .O(N__42910),
            .I(N__42901));
    InMux I__8775 (
            .O(N__42907),
            .I(N__42898));
    Sp12to4 I__8774 (
            .O(N__42904),
            .I(N__42895));
    Span4Mux_h I__8773 (
            .O(N__42901),
            .I(N__42892));
    LocalMux I__8772 (
            .O(N__42898),
            .I(side_order_7));
    Odrv12 I__8771 (
            .O(N__42895),
            .I(side_order_7));
    Odrv4 I__8770 (
            .O(N__42892),
            .I(side_order_7));
    InMux I__8769 (
            .O(N__42885),
            .I(N__42881));
    InMux I__8768 (
            .O(N__42884),
            .I(N__42878));
    LocalMux I__8767 (
            .O(N__42881),
            .I(N__42875));
    LocalMux I__8766 (
            .O(N__42878),
            .I(N__42872));
    Span4Mux_v I__8765 (
            .O(N__42875),
            .I(N__42866));
    Span4Mux_v I__8764 (
            .O(N__42872),
            .I(N__42866));
    CascadeMux I__8763 (
            .O(N__42871),
            .I(N__42863));
    Span4Mux_h I__8762 (
            .O(N__42866),
            .I(N__42860));
    InMux I__8761 (
            .O(N__42863),
            .I(N__42857));
    Span4Mux_v I__8760 (
            .O(N__42860),
            .I(N__42854));
    LocalMux I__8759 (
            .O(N__42857),
            .I(side_order_8));
    Odrv4 I__8758 (
            .O(N__42854),
            .I(side_order_8));
    InMux I__8757 (
            .O(N__42849),
            .I(N__42845));
    InMux I__8756 (
            .O(N__42848),
            .I(N__42842));
    LocalMux I__8755 (
            .O(N__42845),
            .I(N__42839));
    LocalMux I__8754 (
            .O(N__42842),
            .I(N__42836));
    Span4Mux_v I__8753 (
            .O(N__42839),
            .I(N__42832));
    Span4Mux_h I__8752 (
            .O(N__42836),
            .I(N__42829));
    CascadeMux I__8751 (
            .O(N__42835),
            .I(N__42826));
    Span4Mux_h I__8750 (
            .O(N__42832),
            .I(N__42821));
    Span4Mux_v I__8749 (
            .O(N__42829),
            .I(N__42821));
    InMux I__8748 (
            .O(N__42826),
            .I(N__42818));
    Span4Mux_v I__8747 (
            .O(N__42821),
            .I(N__42815));
    LocalMux I__8746 (
            .O(N__42818),
            .I(side_order_9));
    Odrv4 I__8745 (
            .O(N__42815),
            .I(side_order_9));
    InMux I__8744 (
            .O(N__42810),
            .I(N__42805));
    InMux I__8743 (
            .O(N__42809),
            .I(N__42802));
    InMux I__8742 (
            .O(N__42808),
            .I(N__42799));
    LocalMux I__8741 (
            .O(N__42805),
            .I(N__42796));
    LocalMux I__8740 (
            .O(N__42802),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__8739 (
            .O(N__42799),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    Odrv4 I__8738 (
            .O(N__42796),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__8737 (
            .O(N__42789),
            .I(N__42784));
    InMux I__8736 (
            .O(N__42788),
            .I(N__42781));
    InMux I__8735 (
            .O(N__42787),
            .I(N__42778));
    LocalMux I__8734 (
            .O(N__42784),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__8733 (
            .O(N__42781),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__8732 (
            .O(N__42778),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    CascadeMux I__8731 (
            .O(N__42771),
            .I(N__42766));
    InMux I__8730 (
            .O(N__42770),
            .I(N__42763));
    InMux I__8729 (
            .O(N__42769),
            .I(N__42760));
    InMux I__8728 (
            .O(N__42766),
            .I(N__42757));
    LocalMux I__8727 (
            .O(N__42763),
            .I(N__42754));
    LocalMux I__8726 (
            .O(N__42760),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__8725 (
            .O(N__42757),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    Odrv4 I__8724 (
            .O(N__42754),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    CascadeMux I__8723 (
            .O(N__42747),
            .I(N__42742));
    InMux I__8722 (
            .O(N__42746),
            .I(N__42739));
    InMux I__8721 (
            .O(N__42745),
            .I(N__42736));
    InMux I__8720 (
            .O(N__42742),
            .I(N__42733));
    LocalMux I__8719 (
            .O(N__42739),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__8718 (
            .O(N__42736),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__8717 (
            .O(N__42733),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__8716 (
            .O(N__42726),
            .I(N__42723));
    LocalMux I__8715 (
            .O(N__42723),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ));
    InMux I__8714 (
            .O(N__42720),
            .I(N__42715));
    InMux I__8713 (
            .O(N__42719),
            .I(N__42712));
    InMux I__8712 (
            .O(N__42718),
            .I(N__42709));
    LocalMux I__8711 (
            .O(N__42715),
            .I(N__42706));
    LocalMux I__8710 (
            .O(N__42712),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__8709 (
            .O(N__42709),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__8708 (
            .O(N__42706),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    CascadeMux I__8707 (
            .O(N__42699),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ));
    CascadeMux I__8706 (
            .O(N__42696),
            .I(N__42693));
    InMux I__8705 (
            .O(N__42693),
            .I(N__42688));
    InMux I__8704 (
            .O(N__42692),
            .I(N__42685));
    InMux I__8703 (
            .O(N__42691),
            .I(N__42682));
    LocalMux I__8702 (
            .O(N__42688),
            .I(N__42679));
    LocalMux I__8701 (
            .O(N__42685),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__8700 (
            .O(N__42682),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv4 I__8699 (
            .O(N__42679),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__8698 (
            .O(N__42672),
            .I(N__42669));
    LocalMux I__8697 (
            .O(N__42669),
            .I(\ppm_encoder_1.N_139_17 ));
    InMux I__8696 (
            .O(N__42666),
            .I(N__42663));
    LocalMux I__8695 (
            .O(N__42663),
            .I(N__42660));
    Odrv4 I__8694 (
            .O(N__42660),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ));
    CascadeMux I__8693 (
            .O(N__42657),
            .I(\ppm_encoder_1.N_139_17_cascade_ ));
    InMux I__8692 (
            .O(N__42654),
            .I(N__42651));
    LocalMux I__8691 (
            .O(N__42651),
            .I(N__42648));
    Span4Mux_h I__8690 (
            .O(N__42648),
            .I(N__42645));
    Span4Mux_v I__8689 (
            .O(N__42645),
            .I(N__42642));
    Span4Mux_v I__8688 (
            .O(N__42642),
            .I(N__42639));
    Odrv4 I__8687 (
            .O(N__42639),
            .I(\ppm_encoder_1.N_139 ));
    CascadeMux I__8686 (
            .O(N__42636),
            .I(N__42629));
    InMux I__8685 (
            .O(N__42635),
            .I(N__42622));
    InMux I__8684 (
            .O(N__42634),
            .I(N__42622));
    InMux I__8683 (
            .O(N__42633),
            .I(N__42617));
    InMux I__8682 (
            .O(N__42632),
            .I(N__42617));
    InMux I__8681 (
            .O(N__42629),
            .I(N__42614));
    InMux I__8680 (
            .O(N__42628),
            .I(N__42611));
    InMux I__8679 (
            .O(N__42627),
            .I(N__42606));
    LocalMux I__8678 (
            .O(N__42622),
            .I(N__42603));
    LocalMux I__8677 (
            .O(N__42617),
            .I(N__42598));
    LocalMux I__8676 (
            .O(N__42614),
            .I(N__42598));
    LocalMux I__8675 (
            .O(N__42611),
            .I(N__42595));
    InMux I__8674 (
            .O(N__42610),
            .I(N__42590));
    InMux I__8673 (
            .O(N__42609),
            .I(N__42590));
    LocalMux I__8672 (
            .O(N__42606),
            .I(N__42587));
    Span4Mux_h I__8671 (
            .O(N__42603),
            .I(N__42582));
    Span4Mux_h I__8670 (
            .O(N__42598),
            .I(N__42582));
    Span4Mux_h I__8669 (
            .O(N__42595),
            .I(N__42579));
    LocalMux I__8668 (
            .O(N__42590),
            .I(N__42572));
    Span4Mux_v I__8667 (
            .O(N__42587),
            .I(N__42572));
    Span4Mux_v I__8666 (
            .O(N__42582),
            .I(N__42572));
    Odrv4 I__8665 (
            .O(N__42579),
            .I(\pid_front.un1_pid_prereg_92 ));
    Odrv4 I__8664 (
            .O(N__42572),
            .I(\pid_front.un1_pid_prereg_92 ));
    CascadeMux I__8663 (
            .O(N__42567),
            .I(N__42563));
    InMux I__8662 (
            .O(N__42566),
            .I(N__42556));
    InMux I__8661 (
            .O(N__42563),
            .I(N__42556));
    InMux I__8660 (
            .O(N__42562),
            .I(N__42553));
    InMux I__8659 (
            .O(N__42561),
            .I(N__42549));
    LocalMux I__8658 (
            .O(N__42556),
            .I(N__42546));
    LocalMux I__8657 (
            .O(N__42553),
            .I(N__42543));
    CascadeMux I__8656 (
            .O(N__42552),
            .I(N__42540));
    LocalMux I__8655 (
            .O(N__42549),
            .I(N__42536));
    Span4Mux_h I__8654 (
            .O(N__42546),
            .I(N__42531));
    Span4Mux_h I__8653 (
            .O(N__42543),
            .I(N__42531));
    InMux I__8652 (
            .O(N__42540),
            .I(N__42526));
    InMux I__8651 (
            .O(N__42539),
            .I(N__42526));
    Span4Mux_v I__8650 (
            .O(N__42536),
            .I(N__42521));
    Span4Mux_v I__8649 (
            .O(N__42531),
            .I(N__42521));
    LocalMux I__8648 (
            .O(N__42526),
            .I(\pid_front.un1_pid_prereg_93 ));
    Odrv4 I__8647 (
            .O(N__42521),
            .I(\pid_front.un1_pid_prereg_93 ));
    CascadeMux I__8646 (
            .O(N__42516),
            .I(N__42513));
    InMux I__8645 (
            .O(N__42513),
            .I(N__42510));
    LocalMux I__8644 (
            .O(N__42510),
            .I(N__42507));
    Odrv4 I__8643 (
            .O(N__42507),
            .I(\pid_front.error_p_reg_esr_RNIGKTC2Z0Z_20 ));
    InMux I__8642 (
            .O(N__42504),
            .I(N__42501));
    LocalMux I__8641 (
            .O(N__42501),
            .I(N__42498));
    Odrv4 I__8640 (
            .O(N__42498),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    CascadeMux I__8639 (
            .O(N__42495),
            .I(N__42492));
    InMux I__8638 (
            .O(N__42492),
            .I(N__42488));
    InMux I__8637 (
            .O(N__42491),
            .I(N__42485));
    LocalMux I__8636 (
            .O(N__42488),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    LocalMux I__8635 (
            .O(N__42485),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    CascadeMux I__8634 (
            .O(N__42480),
            .I(N__42477));
    InMux I__8633 (
            .O(N__42477),
            .I(N__42471));
    InMux I__8632 (
            .O(N__42476),
            .I(N__42471));
    LocalMux I__8631 (
            .O(N__42471),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__8630 (
            .O(N__42468),
            .I(N__42465));
    LocalMux I__8629 (
            .O(N__42465),
            .I(N__42462));
    Odrv4 I__8628 (
            .O(N__42462),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__8627 (
            .O(N__42459),
            .I(N__42454));
    InMux I__8626 (
            .O(N__42458),
            .I(N__42451));
    IoInMux I__8625 (
            .O(N__42457),
            .I(N__42443));
    LocalMux I__8624 (
            .O(N__42454),
            .I(N__42436));
    LocalMux I__8623 (
            .O(N__42451),
            .I(N__42433));
    CascadeMux I__8622 (
            .O(N__42450),
            .I(N__42429));
    CascadeMux I__8621 (
            .O(N__42449),
            .I(N__42426));
    CascadeMux I__8620 (
            .O(N__42448),
            .I(N__42423));
    CascadeMux I__8619 (
            .O(N__42447),
            .I(N__42420));
    CascadeMux I__8618 (
            .O(N__42446),
            .I(N__42417));
    LocalMux I__8617 (
            .O(N__42443),
            .I(N__42414));
    CascadeMux I__8616 (
            .O(N__42442),
            .I(N__42411));
    CascadeMux I__8615 (
            .O(N__42441),
            .I(N__42408));
    CascadeMux I__8614 (
            .O(N__42440),
            .I(N__42405));
    CascadeMux I__8613 (
            .O(N__42439),
            .I(N__42402));
    Span4Mux_v I__8612 (
            .O(N__42436),
            .I(N__42399));
    Span4Mux_v I__8611 (
            .O(N__42433),
            .I(N__42396));
    InMux I__8610 (
            .O(N__42432),
            .I(N__42393));
    InMux I__8609 (
            .O(N__42429),
            .I(N__42389));
    InMux I__8608 (
            .O(N__42426),
            .I(N__42380));
    InMux I__8607 (
            .O(N__42423),
            .I(N__42380));
    InMux I__8606 (
            .O(N__42420),
            .I(N__42380));
    InMux I__8605 (
            .O(N__42417),
            .I(N__42380));
    Span4Mux_s2_v I__8604 (
            .O(N__42414),
            .I(N__42377));
    InMux I__8603 (
            .O(N__42411),
            .I(N__42374));
    InMux I__8602 (
            .O(N__42408),
            .I(N__42367));
    InMux I__8601 (
            .O(N__42405),
            .I(N__42367));
    InMux I__8600 (
            .O(N__42402),
            .I(N__42367));
    Span4Mux_v I__8599 (
            .O(N__42399),
            .I(N__42356));
    Span4Mux_v I__8598 (
            .O(N__42396),
            .I(N__42356));
    LocalMux I__8597 (
            .O(N__42393),
            .I(N__42356));
    InMux I__8596 (
            .O(N__42392),
            .I(N__42353));
    LocalMux I__8595 (
            .O(N__42389),
            .I(N__42347));
    LocalMux I__8594 (
            .O(N__42380),
            .I(N__42347));
    Span4Mux_v I__8593 (
            .O(N__42377),
            .I(N__42340));
    LocalMux I__8592 (
            .O(N__42374),
            .I(N__42340));
    LocalMux I__8591 (
            .O(N__42367),
            .I(N__42340));
    CascadeMux I__8590 (
            .O(N__42366),
            .I(N__42337));
    CascadeMux I__8589 (
            .O(N__42365),
            .I(N__42333));
    CascadeMux I__8588 (
            .O(N__42364),
            .I(N__42330));
    InMux I__8587 (
            .O(N__42363),
            .I(N__42327));
    Span4Mux_v I__8586 (
            .O(N__42356),
            .I(N__42321));
    LocalMux I__8585 (
            .O(N__42353),
            .I(N__42321));
    CascadeMux I__8584 (
            .O(N__42352),
            .I(N__42318));
    Span4Mux_v I__8583 (
            .O(N__42347),
            .I(N__42310));
    Span4Mux_v I__8582 (
            .O(N__42340),
            .I(N__42310));
    InMux I__8581 (
            .O(N__42337),
            .I(N__42307));
    InMux I__8580 (
            .O(N__42336),
            .I(N__42300));
    InMux I__8579 (
            .O(N__42333),
            .I(N__42300));
    InMux I__8578 (
            .O(N__42330),
            .I(N__42300));
    LocalMux I__8577 (
            .O(N__42327),
            .I(N__42292));
    InMux I__8576 (
            .O(N__42326),
            .I(N__42289));
    Span4Mux_v I__8575 (
            .O(N__42321),
            .I(N__42282));
    InMux I__8574 (
            .O(N__42318),
            .I(N__42279));
    CascadeMux I__8573 (
            .O(N__42317),
            .I(N__42275));
    CascadeMux I__8572 (
            .O(N__42316),
            .I(N__42272));
    CascadeMux I__8571 (
            .O(N__42315),
            .I(N__42269));
    Span4Mux_h I__8570 (
            .O(N__42310),
            .I(N__42262));
    LocalMux I__8569 (
            .O(N__42307),
            .I(N__42262));
    LocalMux I__8568 (
            .O(N__42300),
            .I(N__42262));
    InMux I__8567 (
            .O(N__42299),
            .I(N__42259));
    CascadeMux I__8566 (
            .O(N__42298),
            .I(N__42255));
    CascadeMux I__8565 (
            .O(N__42297),
            .I(N__42252));
    CascadeMux I__8564 (
            .O(N__42296),
            .I(N__42249));
    CascadeMux I__8563 (
            .O(N__42295),
            .I(N__42246));
    Span4Mux_v I__8562 (
            .O(N__42292),
            .I(N__42241));
    LocalMux I__8561 (
            .O(N__42289),
            .I(N__42241));
    InMux I__8560 (
            .O(N__42288),
            .I(N__42238));
    InMux I__8559 (
            .O(N__42287),
            .I(N__42234));
    InMux I__8558 (
            .O(N__42286),
            .I(N__42231));
    InMux I__8557 (
            .O(N__42285),
            .I(N__42225));
    Span4Mux_h I__8556 (
            .O(N__42282),
            .I(N__42222));
    LocalMux I__8555 (
            .O(N__42279),
            .I(N__42219));
    InMux I__8554 (
            .O(N__42278),
            .I(N__42212));
    InMux I__8553 (
            .O(N__42275),
            .I(N__42212));
    InMux I__8552 (
            .O(N__42272),
            .I(N__42212));
    InMux I__8551 (
            .O(N__42269),
            .I(N__42209));
    Span4Mux_v I__8550 (
            .O(N__42262),
            .I(N__42206));
    LocalMux I__8549 (
            .O(N__42259),
            .I(N__42203));
    InMux I__8548 (
            .O(N__42258),
            .I(N__42200));
    InMux I__8547 (
            .O(N__42255),
            .I(N__42197));
    InMux I__8546 (
            .O(N__42252),
            .I(N__42194));
    InMux I__8545 (
            .O(N__42249),
            .I(N__42189));
    InMux I__8544 (
            .O(N__42246),
            .I(N__42189));
    Span4Mux_v I__8543 (
            .O(N__42241),
            .I(N__42184));
    LocalMux I__8542 (
            .O(N__42238),
            .I(N__42184));
    InMux I__8541 (
            .O(N__42237),
            .I(N__42181));
    LocalMux I__8540 (
            .O(N__42234),
            .I(N__42176));
    LocalMux I__8539 (
            .O(N__42231),
            .I(N__42176));
    InMux I__8538 (
            .O(N__42230),
            .I(N__42173));
    InMux I__8537 (
            .O(N__42229),
            .I(N__42170));
    InMux I__8536 (
            .O(N__42228),
            .I(N__42167));
    LocalMux I__8535 (
            .O(N__42225),
            .I(N__42164));
    Span4Mux_h I__8534 (
            .O(N__42222),
            .I(N__42161));
    Span4Mux_v I__8533 (
            .O(N__42219),
            .I(N__42156));
    LocalMux I__8532 (
            .O(N__42212),
            .I(N__42156));
    LocalMux I__8531 (
            .O(N__42209),
            .I(N__42153));
    Span4Mux_h I__8530 (
            .O(N__42206),
            .I(N__42148));
    Span4Mux_v I__8529 (
            .O(N__42203),
            .I(N__42148));
    LocalMux I__8528 (
            .O(N__42200),
            .I(N__42139));
    LocalMux I__8527 (
            .O(N__42197),
            .I(N__42139));
    LocalMux I__8526 (
            .O(N__42194),
            .I(N__42139));
    LocalMux I__8525 (
            .O(N__42189),
            .I(N__42139));
    Span4Mux_v I__8524 (
            .O(N__42184),
            .I(N__42134));
    LocalMux I__8523 (
            .O(N__42181),
            .I(N__42134));
    Span4Mux_v I__8522 (
            .O(N__42176),
            .I(N__42127));
    LocalMux I__8521 (
            .O(N__42173),
            .I(N__42127));
    LocalMux I__8520 (
            .O(N__42170),
            .I(N__42127));
    LocalMux I__8519 (
            .O(N__42167),
            .I(N__42124));
    Span12Mux_s8_h I__8518 (
            .O(N__42164),
            .I(N__42119));
    Sp12to4 I__8517 (
            .O(N__42161),
            .I(N__42119));
    Span4Mux_v I__8516 (
            .O(N__42156),
            .I(N__42114));
    Span4Mux_v I__8515 (
            .O(N__42153),
            .I(N__42114));
    Span4Mux_v I__8514 (
            .O(N__42148),
            .I(N__42109));
    Span4Mux_v I__8513 (
            .O(N__42139),
            .I(N__42109));
    Span4Mux_v I__8512 (
            .O(N__42134),
            .I(N__42104));
    Span4Mux_v I__8511 (
            .O(N__42127),
            .I(N__42104));
    Span12Mux_s8_h I__8510 (
            .O(N__42124),
            .I(N__42095));
    Span12Mux_v I__8509 (
            .O(N__42119),
            .I(N__42095));
    Sp12to4 I__8508 (
            .O(N__42114),
            .I(N__42095));
    Sp12to4 I__8507 (
            .O(N__42109),
            .I(N__42095));
    Span4Mux_h I__8506 (
            .O(N__42104),
            .I(N__42092));
    Odrv12 I__8505 (
            .O(N__42095),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8504 (
            .O(N__42092),
            .I(CONSTANT_ONE_NET));
    InMux I__8503 (
            .O(N__42087),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__8502 (
            .O(N__42084),
            .I(N__42081));
    LocalMux I__8501 (
            .O(N__42081),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    InMux I__8500 (
            .O(N__42078),
            .I(N__42072));
    InMux I__8499 (
            .O(N__42077),
            .I(N__42069));
    InMux I__8498 (
            .O(N__42076),
            .I(N__42064));
    InMux I__8497 (
            .O(N__42075),
            .I(N__42064));
    LocalMux I__8496 (
            .O(N__42072),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__8495 (
            .O(N__42069),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__8494 (
            .O(N__42064),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    CascadeMux I__8493 (
            .O(N__42057),
            .I(N__42053));
    InMux I__8492 (
            .O(N__42056),
            .I(N__42048));
    InMux I__8491 (
            .O(N__42053),
            .I(N__42045));
    InMux I__8490 (
            .O(N__42052),
            .I(N__42040));
    InMux I__8489 (
            .O(N__42051),
            .I(N__42040));
    LocalMux I__8488 (
            .O(N__42048),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__8487 (
            .O(N__42045),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__8486 (
            .O(N__42040),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__8485 (
            .O(N__42033),
            .I(N__42030));
    LocalMux I__8484 (
            .O(N__42030),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    CascadeMux I__8483 (
            .O(N__42027),
            .I(N__42022));
    InMux I__8482 (
            .O(N__42026),
            .I(N__42018));
    InMux I__8481 (
            .O(N__42025),
            .I(N__42015));
    InMux I__8480 (
            .O(N__42022),
            .I(N__42010));
    InMux I__8479 (
            .O(N__42021),
            .I(N__42010));
    LocalMux I__8478 (
            .O(N__42018),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__8477 (
            .O(N__42015),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__8476 (
            .O(N__42010),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__8475 (
            .O(N__42003),
            .I(N__42000));
    LocalMux I__8474 (
            .O(N__42000),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__8473 (
            .O(N__41997),
            .I(N__41994));
    LocalMux I__8472 (
            .O(N__41994),
            .I(N__41991));
    Odrv4 I__8471 (
            .O(N__41991),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    InMux I__8470 (
            .O(N__41988),
            .I(N__41985));
    LocalMux I__8469 (
            .O(N__41985),
            .I(N__41982));
    Odrv4 I__8468 (
            .O(N__41982),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__8467 (
            .O(N__41979),
            .I(N__41976));
    LocalMux I__8466 (
            .O(N__41976),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__8465 (
            .O(N__41973),
            .I(N__41970));
    LocalMux I__8464 (
            .O(N__41970),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ));
    CascadeMux I__8463 (
            .O(N__41967),
            .I(\ppm_encoder_1.N_232_cascade_ ));
    IoInMux I__8462 (
            .O(N__41964),
            .I(N__41961));
    LocalMux I__8461 (
            .O(N__41961),
            .I(N__41958));
    Span4Mux_s1_v I__8460 (
            .O(N__41958),
            .I(N__41955));
    Span4Mux_h I__8459 (
            .O(N__41955),
            .I(N__41952));
    Span4Mux_v I__8458 (
            .O(N__41952),
            .I(N__41949));
    Odrv4 I__8457 (
            .O(N__41949),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__8456 (
            .O(N__41946),
            .I(N__41941));
    InMux I__8455 (
            .O(N__41945),
            .I(N__41938));
    InMux I__8454 (
            .O(N__41944),
            .I(N__41935));
    LocalMux I__8453 (
            .O(N__41941),
            .I(N__41932));
    LocalMux I__8452 (
            .O(N__41938),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__8451 (
            .O(N__41935),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    Odrv4 I__8450 (
            .O(N__41932),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    CascadeMux I__8449 (
            .O(N__41925),
            .I(N__41922));
    InMux I__8448 (
            .O(N__41922),
            .I(N__41917));
    InMux I__8447 (
            .O(N__41921),
            .I(N__41914));
    InMux I__8446 (
            .O(N__41920),
            .I(N__41911));
    LocalMux I__8445 (
            .O(N__41917),
            .I(N__41908));
    LocalMux I__8444 (
            .O(N__41914),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__8443 (
            .O(N__41911),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__8442 (
            .O(N__41908),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__8441 (
            .O(N__41901),
            .I(N__41898));
    LocalMux I__8440 (
            .O(N__41898),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__8439 (
            .O(N__41895),
            .I(N__41892));
    LocalMux I__8438 (
            .O(N__41892),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__8437 (
            .O(N__41889),
            .I(N__41886));
    LocalMux I__8436 (
            .O(N__41886),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__8435 (
            .O(N__41883),
            .I(N__41880));
    LocalMux I__8434 (
            .O(N__41880),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__8433 (
            .O(N__41877),
            .I(N__41874));
    LocalMux I__8432 (
            .O(N__41874),
            .I(N__41869));
    InMux I__8431 (
            .O(N__41873),
            .I(N__41866));
    InMux I__8430 (
            .O(N__41872),
            .I(N__41863));
    Span4Mux_v I__8429 (
            .O(N__41869),
            .I(N__41858));
    LocalMux I__8428 (
            .O(N__41866),
            .I(N__41858));
    LocalMux I__8427 (
            .O(N__41863),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__8426 (
            .O(N__41858),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    InMux I__8425 (
            .O(N__41853),
            .I(N__41849));
    InMux I__8424 (
            .O(N__41852),
            .I(N__41845));
    LocalMux I__8423 (
            .O(N__41849),
            .I(N__41842));
    InMux I__8422 (
            .O(N__41848),
            .I(N__41839));
    LocalMux I__8421 (
            .O(N__41845),
            .I(N__41832));
    Span4Mux_v I__8420 (
            .O(N__41842),
            .I(N__41832));
    LocalMux I__8419 (
            .O(N__41839),
            .I(N__41832));
    Odrv4 I__8418 (
            .O(N__41832),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    InMux I__8417 (
            .O(N__41829),
            .I(N__41826));
    LocalMux I__8416 (
            .O(N__41826),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ));
    InMux I__8415 (
            .O(N__41823),
            .I(N__41820));
    LocalMux I__8414 (
            .O(N__41820),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    InMux I__8413 (
            .O(N__41817),
            .I(N__41814));
    LocalMux I__8412 (
            .O(N__41814),
            .I(N__41811));
    Span4Mux_v I__8411 (
            .O(N__41811),
            .I(N__41808));
    Odrv4 I__8410 (
            .O(N__41808),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    InMux I__8409 (
            .O(N__41805),
            .I(N__41802));
    LocalMux I__8408 (
            .O(N__41802),
            .I(N__41799));
    Span12Mux_v I__8407 (
            .O(N__41799),
            .I(N__41796));
    Odrv12 I__8406 (
            .O(N__41796),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ));
    CascadeMux I__8405 (
            .O(N__41793),
            .I(N__41790));
    InMux I__8404 (
            .O(N__41790),
            .I(N__41787));
    LocalMux I__8403 (
            .O(N__41787),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__8402 (
            .O(N__41784),
            .I(N__41781));
    LocalMux I__8401 (
            .O(N__41781),
            .I(N__41778));
    Span4Mux_v I__8400 (
            .O(N__41778),
            .I(N__41775));
    Span4Mux_v I__8399 (
            .O(N__41775),
            .I(N__41772));
    Odrv4 I__8398 (
            .O(N__41772),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ));
    InMux I__8397 (
            .O(N__41769),
            .I(N__41766));
    LocalMux I__8396 (
            .O(N__41766),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    InMux I__8395 (
            .O(N__41763),
            .I(N__41760));
    LocalMux I__8394 (
            .O(N__41760),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    CascadeMux I__8393 (
            .O(N__41757),
            .I(N__41754));
    InMux I__8392 (
            .O(N__41754),
            .I(N__41751));
    LocalMux I__8391 (
            .O(N__41751),
            .I(N__41748));
    Span4Mux_v I__8390 (
            .O(N__41748),
            .I(N__41745));
    Odrv4 I__8389 (
            .O(N__41745),
            .I(\ppm_encoder_1.elevator_RNIH72D6Z0Z_12 ));
    InMux I__8388 (
            .O(N__41742),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    CascadeMux I__8387 (
            .O(N__41739),
            .I(N__41736));
    InMux I__8386 (
            .O(N__41736),
            .I(N__41733));
    LocalMux I__8385 (
            .O(N__41733),
            .I(N__41730));
    Odrv4 I__8384 (
            .O(N__41730),
            .I(\ppm_encoder_1.elevator_RNIMC2D6Z0Z_13 ));
    InMux I__8383 (
            .O(N__41727),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    CascadeMux I__8382 (
            .O(N__41724),
            .I(N__41721));
    InMux I__8381 (
            .O(N__41721),
            .I(N__41718));
    LocalMux I__8380 (
            .O(N__41718),
            .I(\ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14 ));
    InMux I__8379 (
            .O(N__41715),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__8378 (
            .O(N__41712),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__8377 (
            .O(N__41709),
            .I(bfn_15_19_0_));
    InMux I__8376 (
            .O(N__41706),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__8375 (
            .O(N__41703),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    InMux I__8374 (
            .O(N__41700),
            .I(N__41697));
    LocalMux I__8373 (
            .O(N__41697),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_18 ));
    InMux I__8372 (
            .O(N__41694),
            .I(N__41691));
    LocalMux I__8371 (
            .O(N__41691),
            .I(N__41688));
    Odrv12 I__8370 (
            .O(N__41688),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0 ));
    InMux I__8369 (
            .O(N__41685),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    CascadeMux I__8368 (
            .O(N__41682),
            .I(N__41679));
    InMux I__8367 (
            .O(N__41679),
            .I(N__41676));
    LocalMux I__8366 (
            .O(N__41676),
            .I(N__41673));
    Odrv4 I__8365 (
            .O(N__41673),
            .I(\ppm_encoder_1.elevator_RNIFISN6Z0Z_4 ));
    InMux I__8364 (
            .O(N__41670),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    CascadeMux I__8363 (
            .O(N__41667),
            .I(N__41664));
    InMux I__8362 (
            .O(N__41664),
            .I(N__41661));
    LocalMux I__8361 (
            .O(N__41661),
            .I(N__41658));
    Odrv4 I__8360 (
            .O(N__41658),
            .I(\ppm_encoder_1.elevator_RNIKNSN6Z0Z_5 ));
    InMux I__8359 (
            .O(N__41655),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    CascadeMux I__8358 (
            .O(N__41652),
            .I(N__41649));
    InMux I__8357 (
            .O(N__41649),
            .I(N__41646));
    LocalMux I__8356 (
            .O(N__41646),
            .I(N__41643));
    Odrv4 I__8355 (
            .O(N__41643),
            .I(\ppm_encoder_1.throttle_RNIGQOO6Z0Z_6 ));
    InMux I__8354 (
            .O(N__41640),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    CascadeMux I__8353 (
            .O(N__41637),
            .I(N__41634));
    InMux I__8352 (
            .O(N__41634),
            .I(N__41631));
    LocalMux I__8351 (
            .O(N__41631),
            .I(\ppm_encoder_1.throttle_RNILVOO6Z0Z_7 ));
    InMux I__8350 (
            .O(N__41628),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    CascadeMux I__8349 (
            .O(N__41625),
            .I(N__41622));
    InMux I__8348 (
            .O(N__41622),
            .I(N__41619));
    LocalMux I__8347 (
            .O(N__41619),
            .I(\ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8 ));
    InMux I__8346 (
            .O(N__41616),
            .I(bfn_15_18_0_));
    CascadeMux I__8345 (
            .O(N__41613),
            .I(N__41610));
    InMux I__8344 (
            .O(N__41610),
            .I(N__41607));
    LocalMux I__8343 (
            .O(N__41607),
            .I(N__41604));
    Span4Mux_v I__8342 (
            .O(N__41604),
            .I(N__41601));
    Odrv4 I__8341 (
            .O(N__41601),
            .I(\ppm_encoder_1.throttle_RNIV9PO6Z0Z_9 ));
    InMux I__8340 (
            .O(N__41598),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    CascadeMux I__8339 (
            .O(N__41595),
            .I(N__41592));
    InMux I__8338 (
            .O(N__41592),
            .I(N__41589));
    LocalMux I__8337 (
            .O(N__41589),
            .I(\ppm_encoder_1.elevator_RNI7T1D6Z0Z_10 ));
    InMux I__8336 (
            .O(N__41586),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    CascadeMux I__8335 (
            .O(N__41583),
            .I(N__41580));
    InMux I__8334 (
            .O(N__41580),
            .I(N__41577));
    LocalMux I__8333 (
            .O(N__41577),
            .I(N__41574));
    Span4Mux_v I__8332 (
            .O(N__41574),
            .I(N__41571));
    Odrv4 I__8331 (
            .O(N__41571),
            .I(\ppm_encoder_1.elevator_RNIC22D6Z0Z_11 ));
    InMux I__8330 (
            .O(N__41568),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    CascadeMux I__8329 (
            .O(N__41565),
            .I(\ppm_encoder_1.N_287_cascade_ ));
    CascadeMux I__8328 (
            .O(N__41562),
            .I(N__41559));
    InMux I__8327 (
            .O(N__41559),
            .I(N__41556));
    LocalMux I__8326 (
            .O(N__41556),
            .I(N__41553));
    Span4Mux_v I__8325 (
            .O(N__41553),
            .I(N__41550));
    Odrv4 I__8324 (
            .O(N__41550),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ));
    InMux I__8323 (
            .O(N__41547),
            .I(N__41543));
    InMux I__8322 (
            .O(N__41546),
            .I(N__41540));
    LocalMux I__8321 (
            .O(N__41543),
            .I(N__41537));
    LocalMux I__8320 (
            .O(N__41540),
            .I(N__41534));
    Span12Mux_v I__8319 (
            .O(N__41537),
            .I(N__41531));
    Odrv4 I__8318 (
            .O(N__41534),
            .I(side_order_1));
    Odrv12 I__8317 (
            .O(N__41531),
            .I(side_order_1));
    CascadeMux I__8316 (
            .O(N__41526),
            .I(N__41523));
    InMux I__8315 (
            .O(N__41523),
            .I(N__41520));
    LocalMux I__8314 (
            .O(N__41520),
            .I(N__41517));
    Span4Mux_v I__8313 (
            .O(N__41517),
            .I(N__41514));
    Odrv4 I__8312 (
            .O(N__41514),
            .I(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ));
    InMux I__8311 (
            .O(N__41511),
            .I(N__41506));
    InMux I__8310 (
            .O(N__41510),
            .I(N__41501));
    InMux I__8309 (
            .O(N__41509),
            .I(N__41501));
    LocalMux I__8308 (
            .O(N__41506),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    LocalMux I__8307 (
            .O(N__41501),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    InMux I__8306 (
            .O(N__41496),
            .I(N__41493));
    LocalMux I__8305 (
            .O(N__41493),
            .I(N__41490));
    Odrv4 I__8304 (
            .O(N__41490),
            .I(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ));
    CascadeMux I__8303 (
            .O(N__41487),
            .I(N__41484));
    InMux I__8302 (
            .O(N__41484),
            .I(N__41481));
    LocalMux I__8301 (
            .O(N__41481),
            .I(N__41477));
    InMux I__8300 (
            .O(N__41480),
            .I(N__41474));
    Span4Mux_h I__8299 (
            .O(N__41477),
            .I(N__41469));
    LocalMux I__8298 (
            .O(N__41474),
            .I(N__41469));
    Span4Mux_h I__8297 (
            .O(N__41469),
            .I(N__41466));
    Odrv4 I__8296 (
            .O(N__41466),
            .I(front_order_1));
    InMux I__8295 (
            .O(N__41463),
            .I(N__41454));
    InMux I__8294 (
            .O(N__41462),
            .I(N__41454));
    InMux I__8293 (
            .O(N__41461),
            .I(N__41454));
    LocalMux I__8292 (
            .O(N__41454),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    InMux I__8291 (
            .O(N__41451),
            .I(N__41448));
    LocalMux I__8290 (
            .O(N__41448),
            .I(N__41445));
    Span4Mux_h I__8289 (
            .O(N__41445),
            .I(N__41442));
    Odrv4 I__8288 (
            .O(N__41442),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    InMux I__8287 (
            .O(N__41439),
            .I(N__41436));
    LocalMux I__8286 (
            .O(N__41436),
            .I(N__41432));
    InMux I__8285 (
            .O(N__41435),
            .I(N__41429));
    Span4Mux_v I__8284 (
            .O(N__41432),
            .I(N__41426));
    LocalMux I__8283 (
            .O(N__41429),
            .I(N__41423));
    Span4Mux_h I__8282 (
            .O(N__41426),
            .I(N__41418));
    Span4Mux_v I__8281 (
            .O(N__41423),
            .I(N__41418));
    Span4Mux_h I__8280 (
            .O(N__41418),
            .I(N__41415));
    Odrv4 I__8279 (
            .O(N__41415),
            .I(throttle_order_1));
    InMux I__8278 (
            .O(N__41412),
            .I(N__41403));
    InMux I__8277 (
            .O(N__41411),
            .I(N__41403));
    InMux I__8276 (
            .O(N__41410),
            .I(N__41403));
    LocalMux I__8275 (
            .O(N__41403),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    CascadeMux I__8274 (
            .O(N__41400),
            .I(N__41397));
    InMux I__8273 (
            .O(N__41397),
            .I(N__41394));
    LocalMux I__8272 (
            .O(N__41394),
            .I(\ppm_encoder_1.throttle_RNIUINC6Z0Z_1 ));
    InMux I__8271 (
            .O(N__41391),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__8270 (
            .O(N__41388),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    CascadeMux I__8269 (
            .O(N__41385),
            .I(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ));
    InMux I__8268 (
            .O(N__41382),
            .I(N__41379));
    LocalMux I__8267 (
            .O(N__41379),
            .I(\ppm_encoder_1.un2_throttle_iv_1_4 ));
    CascadeMux I__8266 (
            .O(N__41376),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ));
    CascadeMux I__8265 (
            .O(N__41373),
            .I(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ));
    InMux I__8264 (
            .O(N__41370),
            .I(N__41367));
    LocalMux I__8263 (
            .O(N__41367),
            .I(\ppm_encoder_1.un2_throttle_iv_1_5 ));
    CascadeMux I__8262 (
            .O(N__41364),
            .I(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ));
    CascadeMux I__8261 (
            .O(N__41361),
            .I(N__41358));
    InMux I__8260 (
            .O(N__41358),
            .I(N__41349));
    InMux I__8259 (
            .O(N__41357),
            .I(N__41345));
    CascadeMux I__8258 (
            .O(N__41356),
            .I(N__41342));
    CascadeMux I__8257 (
            .O(N__41355),
            .I(N__41339));
    CascadeMux I__8256 (
            .O(N__41354),
            .I(N__41336));
    CascadeMux I__8255 (
            .O(N__41353),
            .I(N__41333));
    CascadeMux I__8254 (
            .O(N__41352),
            .I(N__41329));
    LocalMux I__8253 (
            .O(N__41349),
            .I(N__41324));
    InMux I__8252 (
            .O(N__41348),
            .I(N__41321));
    LocalMux I__8251 (
            .O(N__41345),
            .I(N__41318));
    InMux I__8250 (
            .O(N__41342),
            .I(N__41313));
    InMux I__8249 (
            .O(N__41339),
            .I(N__41313));
    InMux I__8248 (
            .O(N__41336),
            .I(N__41310));
    InMux I__8247 (
            .O(N__41333),
            .I(N__41307));
    InMux I__8246 (
            .O(N__41332),
            .I(N__41304));
    InMux I__8245 (
            .O(N__41329),
            .I(N__41301));
    InMux I__8244 (
            .O(N__41328),
            .I(N__41298));
    InMux I__8243 (
            .O(N__41327),
            .I(N__41295));
    Span4Mux_h I__8242 (
            .O(N__41324),
            .I(N__41286));
    LocalMux I__8241 (
            .O(N__41321),
            .I(N__41286));
    Span4Mux_v I__8240 (
            .O(N__41318),
            .I(N__41286));
    LocalMux I__8239 (
            .O(N__41313),
            .I(N__41286));
    LocalMux I__8238 (
            .O(N__41310),
            .I(N__41281));
    LocalMux I__8237 (
            .O(N__41307),
            .I(N__41281));
    LocalMux I__8236 (
            .O(N__41304),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__8235 (
            .O(N__41301),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__8234 (
            .O(N__41298),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__8233 (
            .O(N__41295),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__8232 (
            .O(N__41286),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__8231 (
            .O(N__41281),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    InMux I__8230 (
            .O(N__41268),
            .I(N__41265));
    LocalMux I__8229 (
            .O(N__41265),
            .I(\ppm_encoder_1.throttle_m_1 ));
    CascadeMux I__8228 (
            .O(N__41262),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ));
    InMux I__8227 (
            .O(N__41259),
            .I(N__41255));
    InMux I__8226 (
            .O(N__41258),
            .I(N__41252));
    LocalMux I__8225 (
            .O(N__41255),
            .I(N__41249));
    LocalMux I__8224 (
            .O(N__41252),
            .I(N__41246));
    Span4Mux_h I__8223 (
            .O(N__41249),
            .I(N__41242));
    Span4Mux_v I__8222 (
            .O(N__41246),
            .I(N__41239));
    CascadeMux I__8221 (
            .O(N__41245),
            .I(N__41236));
    Span4Mux_v I__8220 (
            .O(N__41242),
            .I(N__41232));
    Span4Mux_h I__8219 (
            .O(N__41239),
            .I(N__41229));
    InMux I__8218 (
            .O(N__41236),
            .I(N__41224));
    InMux I__8217 (
            .O(N__41235),
            .I(N__41224));
    Odrv4 I__8216 (
            .O(N__41232),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv4 I__8215 (
            .O(N__41229),
            .I(\scaler_4.un2_source_data_0 ));
    LocalMux I__8214 (
            .O(N__41224),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__8213 (
            .O(N__41217),
            .I(N__41214));
    LocalMux I__8212 (
            .O(N__41214),
            .I(N__41210));
    InMux I__8211 (
            .O(N__41213),
            .I(N__41207));
    Span4Mux_v I__8210 (
            .O(N__41210),
            .I(N__41201));
    LocalMux I__8209 (
            .O(N__41207),
            .I(N__41201));
    CascadeMux I__8208 (
            .O(N__41206),
            .I(N__41198));
    Span4Mux_h I__8207 (
            .O(N__41201),
            .I(N__41194));
    InMux I__8206 (
            .O(N__41198),
            .I(N__41191));
    InMux I__8205 (
            .O(N__41197),
            .I(N__41188));
    Span4Mux_h I__8204 (
            .O(N__41194),
            .I(N__41185));
    LocalMux I__8203 (
            .O(N__41191),
            .I(N__41182));
    LocalMux I__8202 (
            .O(N__41188),
            .I(frame_decoder_OFF4data_0));
    Odrv4 I__8201 (
            .O(N__41185),
            .I(frame_decoder_OFF4data_0));
    Odrv12 I__8200 (
            .O(N__41182),
            .I(frame_decoder_OFF4data_0));
    InMux I__8199 (
            .O(N__41175),
            .I(N__41170));
    InMux I__8198 (
            .O(N__41174),
            .I(N__41167));
    InMux I__8197 (
            .O(N__41173),
            .I(N__41164));
    LocalMux I__8196 (
            .O(N__41170),
            .I(N__41161));
    LocalMux I__8195 (
            .O(N__41167),
            .I(N__41157));
    LocalMux I__8194 (
            .O(N__41164),
            .I(N__41154));
    Span4Mux_h I__8193 (
            .O(N__41161),
            .I(N__41151));
    InMux I__8192 (
            .O(N__41160),
            .I(N__41148));
    Odrv12 I__8191 (
            .O(N__41157),
            .I(frame_decoder_CH4data_0));
    Odrv4 I__8190 (
            .O(N__41154),
            .I(frame_decoder_CH4data_0));
    Odrv4 I__8189 (
            .O(N__41151),
            .I(frame_decoder_CH4data_0));
    LocalMux I__8188 (
            .O(N__41148),
            .I(frame_decoder_CH4data_0));
    CascadeMux I__8187 (
            .O(N__41139),
            .I(N__41136));
    InMux I__8186 (
            .O(N__41136),
            .I(N__41133));
    LocalMux I__8185 (
            .O(N__41133),
            .I(N__41130));
    Span4Mux_h I__8184 (
            .O(N__41130),
            .I(N__41127));
    Odrv4 I__8183 (
            .O(N__41127),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ));
    InMux I__8182 (
            .O(N__41124),
            .I(N__41120));
    InMux I__8181 (
            .O(N__41123),
            .I(N__41117));
    LocalMux I__8180 (
            .O(N__41120),
            .I(N__41114));
    LocalMux I__8179 (
            .O(N__41117),
            .I(N__41109));
    Span4Mux_v I__8178 (
            .O(N__41114),
            .I(N__41109));
    Span4Mux_h I__8177 (
            .O(N__41109),
            .I(N__41106));
    Odrv4 I__8176 (
            .O(N__41106),
            .I(side_order_2));
    InMux I__8175 (
            .O(N__41103),
            .I(N__41099));
    InMux I__8174 (
            .O(N__41102),
            .I(N__41096));
    LocalMux I__8173 (
            .O(N__41099),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__8172 (
            .O(N__41096),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    CascadeMux I__8171 (
            .O(N__41091),
            .I(\ppm_encoder_1.N_221_cascade_ ));
    CascadeMux I__8170 (
            .O(N__41088),
            .I(\ppm_encoder_1.N_313_cascade_ ));
    InMux I__8169 (
            .O(N__41085),
            .I(N__41082));
    LocalMux I__8168 (
            .O(N__41082),
            .I(\ppm_encoder_1.un2_throttle_iv_0_12 ));
    InMux I__8167 (
            .O(N__41079),
            .I(N__41076));
    LocalMux I__8166 (
            .O(N__41076),
            .I(\ppm_encoder_1.un2_throttle_iv_1_12 ));
    CascadeMux I__8165 (
            .O(N__41073),
            .I(N__41069));
    InMux I__8164 (
            .O(N__41072),
            .I(N__41066));
    InMux I__8163 (
            .O(N__41069),
            .I(N__41063));
    LocalMux I__8162 (
            .O(N__41066),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    LocalMux I__8161 (
            .O(N__41063),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    InMux I__8160 (
            .O(N__41058),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__8159 (
            .O(N__41055),
            .I(bfn_14_25_0_));
    InMux I__8158 (
            .O(N__41052),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__8157 (
            .O(N__41049),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    SRMux I__8156 (
            .O(N__41046),
            .I(N__41037));
    SRMux I__8155 (
            .O(N__41045),
            .I(N__41037));
    SRMux I__8154 (
            .O(N__41044),
            .I(N__41037));
    GlobalMux I__8153 (
            .O(N__41037),
            .I(N__41034));
    gio2CtrlBuf I__8152 (
            .O(N__41034),
            .I(\ppm_encoder_1.N_419_g ));
    IoInMux I__8151 (
            .O(N__41031),
            .I(N__41028));
    LocalMux I__8150 (
            .O(N__41028),
            .I(N__41025));
    Span4Mux_s2_v I__8149 (
            .O(N__41025),
            .I(N__41022));
    Span4Mux_v I__8148 (
            .O(N__41022),
            .I(N__41018));
    InMux I__8147 (
            .O(N__41021),
            .I(N__41015));
    Span4Mux_v I__8146 (
            .O(N__41018),
            .I(N__41010));
    LocalMux I__8145 (
            .O(N__41015),
            .I(N__41010));
    Span4Mux_h I__8144 (
            .O(N__41010),
            .I(N__41005));
    CascadeMux I__8143 (
            .O(N__41009),
            .I(N__41002));
    InMux I__8142 (
            .O(N__41008),
            .I(N__40999));
    Span4Mux_h I__8141 (
            .O(N__41005),
            .I(N__40996));
    InMux I__8140 (
            .O(N__41002),
            .I(N__40993));
    LocalMux I__8139 (
            .O(N__40999),
            .I(N__40990));
    Odrv4 I__8138 (
            .O(N__40996),
            .I(debug_CH3_20A_c));
    LocalMux I__8137 (
            .O(N__40993),
            .I(debug_CH3_20A_c));
    Odrv4 I__8136 (
            .O(N__40990),
            .I(debug_CH3_20A_c));
    InMux I__8135 (
            .O(N__40983),
            .I(N__40976));
    InMux I__8134 (
            .O(N__40982),
            .I(N__40971));
    InMux I__8133 (
            .O(N__40981),
            .I(N__40965));
    InMux I__8132 (
            .O(N__40980),
            .I(N__40961));
    InMux I__8131 (
            .O(N__40979),
            .I(N__40958));
    LocalMux I__8130 (
            .O(N__40976),
            .I(N__40955));
    InMux I__8129 (
            .O(N__40975),
            .I(N__40952));
    InMux I__8128 (
            .O(N__40974),
            .I(N__40949));
    LocalMux I__8127 (
            .O(N__40971),
            .I(N__40946));
    InMux I__8126 (
            .O(N__40970),
            .I(N__40938));
    InMux I__8125 (
            .O(N__40969),
            .I(N__40938));
    InMux I__8124 (
            .O(N__40968),
            .I(N__40935));
    LocalMux I__8123 (
            .O(N__40965),
            .I(N__40932));
    InMux I__8122 (
            .O(N__40964),
            .I(N__40929));
    LocalMux I__8121 (
            .O(N__40961),
            .I(N__40924));
    LocalMux I__8120 (
            .O(N__40958),
            .I(N__40924));
    Span4Mux_h I__8119 (
            .O(N__40955),
            .I(N__40919));
    LocalMux I__8118 (
            .O(N__40952),
            .I(N__40919));
    LocalMux I__8117 (
            .O(N__40949),
            .I(N__40914));
    Span4Mux_h I__8116 (
            .O(N__40946),
            .I(N__40914));
    InMux I__8115 (
            .O(N__40945),
            .I(N__40909));
    InMux I__8114 (
            .O(N__40944),
            .I(N__40909));
    InMux I__8113 (
            .O(N__40943),
            .I(N__40906));
    LocalMux I__8112 (
            .O(N__40938),
            .I(N__40897));
    LocalMux I__8111 (
            .O(N__40935),
            .I(N__40897));
    Span4Mux_v I__8110 (
            .O(N__40932),
            .I(N__40897));
    LocalMux I__8109 (
            .O(N__40929),
            .I(N__40897));
    Span4Mux_v I__8108 (
            .O(N__40924),
            .I(N__40894));
    Span4Mux_v I__8107 (
            .O(N__40919),
            .I(N__40891));
    Span4Mux_h I__8106 (
            .O(N__40914),
            .I(N__40882));
    LocalMux I__8105 (
            .O(N__40909),
            .I(N__40882));
    LocalMux I__8104 (
            .O(N__40906),
            .I(N__40882));
    Span4Mux_v I__8103 (
            .O(N__40897),
            .I(N__40882));
    Odrv4 I__8102 (
            .O(N__40894),
            .I(uart_drone_data_rdy));
    Odrv4 I__8101 (
            .O(N__40891),
            .I(uart_drone_data_rdy));
    Odrv4 I__8100 (
            .O(N__40882),
            .I(uart_drone_data_rdy));
    SRMux I__8099 (
            .O(N__40875),
            .I(N__40872));
    LocalMux I__8098 (
            .O(N__40872),
            .I(N__40868));
    SRMux I__8097 (
            .O(N__40871),
            .I(N__40865));
    Span4Mux_v I__8096 (
            .O(N__40868),
            .I(N__40860));
    LocalMux I__8095 (
            .O(N__40865),
            .I(N__40860));
    Span4Mux_v I__8094 (
            .O(N__40860),
            .I(N__40857));
    Span4Mux_h I__8093 (
            .O(N__40857),
            .I(N__40854));
    Odrv4 I__8092 (
            .O(N__40854),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    InMux I__8091 (
            .O(N__40851),
            .I(N__40846));
    InMux I__8090 (
            .O(N__40850),
            .I(N__40843));
    InMux I__8089 (
            .O(N__40849),
            .I(N__40840));
    LocalMux I__8088 (
            .O(N__40846),
            .I(N__40837));
    LocalMux I__8087 (
            .O(N__40843),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    LocalMux I__8086 (
            .O(N__40840),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__8085 (
            .O(N__40837),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    InMux I__8084 (
            .O(N__40830),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__8083 (
            .O(N__40827),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    InMux I__8082 (
            .O(N__40824),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__8081 (
            .O(N__40821),
            .I(bfn_14_24_0_));
    InMux I__8080 (
            .O(N__40818),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__8079 (
            .O(N__40815),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__8078 (
            .O(N__40812),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__8077 (
            .O(N__40809),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__8076 (
            .O(N__40806),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__8075 (
            .O(N__40803),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__8074 (
            .O(N__40800),
            .I(N__40797));
    LocalMux I__8073 (
            .O(N__40797),
            .I(N__40794));
    Odrv4 I__8072 (
            .O(N__40794),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ));
    InMux I__8071 (
            .O(N__40791),
            .I(N__40788));
    LocalMux I__8070 (
            .O(N__40788),
            .I(N__40785));
    Span12Mux_s9_v I__8069 (
            .O(N__40785),
            .I(N__40782));
    Odrv12 I__8068 (
            .O(N__40782),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ));
    InMux I__8067 (
            .O(N__40779),
            .I(N__40776));
    LocalMux I__8066 (
            .O(N__40776),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    CascadeMux I__8065 (
            .O(N__40773),
            .I(N__40770));
    InMux I__8064 (
            .O(N__40770),
            .I(N__40767));
    LocalMux I__8063 (
            .O(N__40767),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    CascadeMux I__8062 (
            .O(N__40764),
            .I(N__40760));
    InMux I__8061 (
            .O(N__40763),
            .I(N__40757));
    InMux I__8060 (
            .O(N__40760),
            .I(N__40754));
    LocalMux I__8059 (
            .O(N__40757),
            .I(N__40749));
    LocalMux I__8058 (
            .O(N__40754),
            .I(N__40749));
    Span4Mux_v I__8057 (
            .O(N__40749),
            .I(N__40746));
    Odrv4 I__8056 (
            .O(N__40746),
            .I(\ppm_encoder_1.N_2150_i ));
    InMux I__8055 (
            .O(N__40743),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    InMux I__8054 (
            .O(N__40740),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__8053 (
            .O(N__40737),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__8052 (
            .O(N__40734),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    CascadeMux I__8051 (
            .O(N__40731),
            .I(N__40728));
    InMux I__8050 (
            .O(N__40728),
            .I(N__40725));
    LocalMux I__8049 (
            .O(N__40725),
            .I(N__40722));
    Span4Mux_v I__8048 (
            .O(N__40722),
            .I(N__40718));
    InMux I__8047 (
            .O(N__40721),
            .I(N__40715));
    Odrv4 I__8046 (
            .O(N__40718),
            .I(drone_H_disp_front_13));
    LocalMux I__8045 (
            .O(N__40715),
            .I(drone_H_disp_front_13));
    InMux I__8044 (
            .O(N__40710),
            .I(N__40707));
    LocalMux I__8043 (
            .O(N__40707),
            .I(N__40704));
    Span4Mux_v I__8042 (
            .O(N__40704),
            .I(N__40701));
    Odrv4 I__8041 (
            .O(N__40701),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ));
    InMux I__8040 (
            .O(N__40698),
            .I(N__40695));
    LocalMux I__8039 (
            .O(N__40695),
            .I(N__40692));
    Odrv4 I__8038 (
            .O(N__40692),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ));
    InMux I__8037 (
            .O(N__40689),
            .I(N__40686));
    LocalMux I__8036 (
            .O(N__40686),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__8035 (
            .O(N__40683),
            .I(N__40680));
    LocalMux I__8034 (
            .O(N__40680),
            .I(N__40677));
    Odrv4 I__8033 (
            .O(N__40677),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ));
    InMux I__8032 (
            .O(N__40674),
            .I(N__40671));
    LocalMux I__8031 (
            .O(N__40671),
            .I(N__40668));
    Span4Mux_v I__8030 (
            .O(N__40668),
            .I(N__40665));
    Odrv4 I__8029 (
            .O(N__40665),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ));
    CascadeMux I__8028 (
            .O(N__40662),
            .I(N__40659));
    InMux I__8027 (
            .O(N__40659),
            .I(N__40656));
    LocalMux I__8026 (
            .O(N__40656),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__8025 (
            .O(N__40653),
            .I(N__40650));
    LocalMux I__8024 (
            .O(N__40650),
            .I(N__40647));
    Odrv4 I__8023 (
            .O(N__40647),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ));
    InMux I__8022 (
            .O(N__40644),
            .I(N__40641));
    LocalMux I__8021 (
            .O(N__40641),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__8020 (
            .O(N__40638),
            .I(N__40635));
    LocalMux I__8019 (
            .O(N__40635),
            .I(N__40632));
    Span4Mux_v I__8018 (
            .O(N__40632),
            .I(N__40629));
    Odrv4 I__8017 (
            .O(N__40629),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ));
    InMux I__8016 (
            .O(N__40626),
            .I(N__40623));
    LocalMux I__8015 (
            .O(N__40623),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    InMux I__8014 (
            .O(N__40620),
            .I(N__40617));
    LocalMux I__8013 (
            .O(N__40617),
            .I(N__40614));
    Odrv12 I__8012 (
            .O(N__40614),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__8011 (
            .O(N__40611),
            .I(N__40607));
    InMux I__8010 (
            .O(N__40610),
            .I(N__40603));
    LocalMux I__8009 (
            .O(N__40607),
            .I(N__40600));
    InMux I__8008 (
            .O(N__40606),
            .I(N__40597));
    LocalMux I__8007 (
            .O(N__40603),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__8006 (
            .O(N__40600),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    LocalMux I__8005 (
            .O(N__40597),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    CascadeMux I__8004 (
            .O(N__40590),
            .I(\ppm_encoder_1.un2_throttle_iv_1_10_cascade_ ));
    InMux I__8003 (
            .O(N__40587),
            .I(N__40584));
    LocalMux I__8002 (
            .O(N__40584),
            .I(\ppm_encoder_1.un2_throttle_iv_0_10 ));
    InMux I__8001 (
            .O(N__40581),
            .I(N__40578));
    LocalMux I__8000 (
            .O(N__40578),
            .I(N__40573));
    InMux I__7999 (
            .O(N__40577),
            .I(N__40570));
    InMux I__7998 (
            .O(N__40576),
            .I(N__40567));
    Span4Mux_v I__7997 (
            .O(N__40573),
            .I(N__40562));
    LocalMux I__7996 (
            .O(N__40570),
            .I(N__40562));
    LocalMux I__7995 (
            .O(N__40567),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__7994 (
            .O(N__40562),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    InMux I__7993 (
            .O(N__40557),
            .I(N__40554));
    LocalMux I__7992 (
            .O(N__40554),
            .I(N__40549));
    InMux I__7991 (
            .O(N__40553),
            .I(N__40546));
    CascadeMux I__7990 (
            .O(N__40552),
            .I(N__40543));
    Span4Mux_v I__7989 (
            .O(N__40549),
            .I(N__40538));
    LocalMux I__7988 (
            .O(N__40546),
            .I(N__40538));
    InMux I__7987 (
            .O(N__40543),
            .I(N__40535));
    Span4Mux_h I__7986 (
            .O(N__40538),
            .I(N__40532));
    LocalMux I__7985 (
            .O(N__40535),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__7984 (
            .O(N__40532),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__7983 (
            .O(N__40527),
            .I(N__40521));
    InMux I__7982 (
            .O(N__40526),
            .I(N__40521));
    LocalMux I__7981 (
            .O(N__40521),
            .I(N__40517));
    InMux I__7980 (
            .O(N__40520),
            .I(N__40514));
    Span4Mux_h I__7979 (
            .O(N__40517),
            .I(N__40511));
    LocalMux I__7978 (
            .O(N__40514),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__7977 (
            .O(N__40511),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    CascadeMux I__7976 (
            .O(N__40506),
            .I(\ppm_encoder_1.N_296_cascade_ ));
    InMux I__7975 (
            .O(N__40503),
            .I(N__40497));
    InMux I__7974 (
            .O(N__40502),
            .I(N__40497));
    LocalMux I__7973 (
            .O(N__40497),
            .I(N__40493));
    InMux I__7972 (
            .O(N__40496),
            .I(N__40490));
    Span4Mux_h I__7971 (
            .O(N__40493),
            .I(N__40487));
    LocalMux I__7970 (
            .O(N__40490),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    Odrv4 I__7969 (
            .O(N__40487),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__7968 (
            .O(N__40482),
            .I(N__40479));
    LocalMux I__7967 (
            .O(N__40479),
            .I(\ppm_encoder_1.un2_throttle_iv_1_8 ));
    InMux I__7966 (
            .O(N__40476),
            .I(N__40470));
    InMux I__7965 (
            .O(N__40475),
            .I(N__40470));
    LocalMux I__7964 (
            .O(N__40470),
            .I(N__40466));
    InMux I__7963 (
            .O(N__40469),
            .I(N__40463));
    Span4Mux_h I__7962 (
            .O(N__40466),
            .I(N__40460));
    LocalMux I__7961 (
            .O(N__40463),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    Odrv4 I__7960 (
            .O(N__40460),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    InMux I__7959 (
            .O(N__40455),
            .I(N__40450));
    InMux I__7958 (
            .O(N__40454),
            .I(N__40445));
    InMux I__7957 (
            .O(N__40453),
            .I(N__40445));
    LocalMux I__7956 (
            .O(N__40450),
            .I(N__40442));
    LocalMux I__7955 (
            .O(N__40445),
            .I(N__40439));
    Odrv4 I__7954 (
            .O(N__40442),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    Odrv4 I__7953 (
            .O(N__40439),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    CascadeMux I__7952 (
            .O(N__40434),
            .I(\ppm_encoder_1.N_294_cascade_ ));
    InMux I__7951 (
            .O(N__40431),
            .I(N__40428));
    LocalMux I__7950 (
            .O(N__40428),
            .I(N__40425));
    Span4Mux_v I__7949 (
            .O(N__40425),
            .I(N__40422));
    Odrv4 I__7948 (
            .O(N__40422),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__7947 (
            .O(N__40419),
            .I(N__40410));
    InMux I__7946 (
            .O(N__40418),
            .I(N__40410));
    InMux I__7945 (
            .O(N__40417),
            .I(N__40410));
    LocalMux I__7944 (
            .O(N__40410),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    CascadeMux I__7943 (
            .O(N__40407),
            .I(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ));
    InMux I__7942 (
            .O(N__40404),
            .I(N__40401));
    LocalMux I__7941 (
            .O(N__40401),
            .I(\ppm_encoder_1.un2_throttle_iv_1_14 ));
    InMux I__7940 (
            .O(N__40398),
            .I(N__40392));
    InMux I__7939 (
            .O(N__40397),
            .I(N__40392));
    LocalMux I__7938 (
            .O(N__40392),
            .I(N__40389));
    Odrv4 I__7937 (
            .O(N__40389),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    InMux I__7936 (
            .O(N__40386),
            .I(N__40382));
    InMux I__7935 (
            .O(N__40385),
            .I(N__40379));
    LocalMux I__7934 (
            .O(N__40382),
            .I(N__40374));
    LocalMux I__7933 (
            .O(N__40379),
            .I(N__40374));
    Span4Mux_h I__7932 (
            .O(N__40374),
            .I(N__40371));
    Odrv4 I__7931 (
            .O(N__40371),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    CascadeMux I__7930 (
            .O(N__40368),
            .I(\ppm_encoder_1.N_300_cascade_ ));
    InMux I__7929 (
            .O(N__40365),
            .I(N__40359));
    InMux I__7928 (
            .O(N__40364),
            .I(N__40359));
    LocalMux I__7927 (
            .O(N__40359),
            .I(N__40356));
    Odrv12 I__7926 (
            .O(N__40356),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    CascadeMux I__7925 (
            .O(N__40353),
            .I(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ));
    InMux I__7924 (
            .O(N__40350),
            .I(N__40347));
    LocalMux I__7923 (
            .O(N__40347),
            .I(\ppm_encoder_1.un2_throttle_iv_1_7 ));
    InMux I__7922 (
            .O(N__40344),
            .I(N__40337));
    InMux I__7921 (
            .O(N__40343),
            .I(N__40337));
    InMux I__7920 (
            .O(N__40342),
            .I(N__40334));
    LocalMux I__7919 (
            .O(N__40337),
            .I(N__40331));
    LocalMux I__7918 (
            .O(N__40334),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    Odrv12 I__7917 (
            .O(N__40331),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    CascadeMux I__7916 (
            .O(N__40326),
            .I(\ppm_encoder_1.N_293_cascade_ ));
    InMux I__7915 (
            .O(N__40323),
            .I(N__40320));
    LocalMux I__7914 (
            .O(N__40320),
            .I(N__40317));
    Span4Mux_h I__7913 (
            .O(N__40317),
            .I(N__40314));
    Odrv4 I__7912 (
            .O(N__40314),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__7911 (
            .O(N__40311),
            .I(N__40302));
    InMux I__7910 (
            .O(N__40310),
            .I(N__40302));
    InMux I__7909 (
            .O(N__40309),
            .I(N__40302));
    LocalMux I__7908 (
            .O(N__40302),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    InMux I__7907 (
            .O(N__40299),
            .I(N__40296));
    LocalMux I__7906 (
            .O(N__40296),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__7905 (
            .O(N__40293),
            .I(N__40288));
    InMux I__7904 (
            .O(N__40292),
            .I(N__40285));
    CascadeMux I__7903 (
            .O(N__40291),
            .I(N__40282));
    LocalMux I__7902 (
            .O(N__40288),
            .I(N__40277));
    LocalMux I__7901 (
            .O(N__40285),
            .I(N__40277));
    InMux I__7900 (
            .O(N__40282),
            .I(N__40274));
    Span4Mux_v I__7899 (
            .O(N__40277),
            .I(N__40271));
    LocalMux I__7898 (
            .O(N__40274),
            .I(front_order_7));
    Odrv4 I__7897 (
            .O(N__40271),
            .I(front_order_7));
    InMux I__7896 (
            .O(N__40266),
            .I(N__40257));
    InMux I__7895 (
            .O(N__40265),
            .I(N__40257));
    InMux I__7894 (
            .O(N__40264),
            .I(N__40257));
    LocalMux I__7893 (
            .O(N__40257),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    CascadeMux I__7892 (
            .O(N__40254),
            .I(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ));
    CascadeMux I__7891 (
            .O(N__40251),
            .I(N__40246));
    InMux I__7890 (
            .O(N__40250),
            .I(N__40241));
    InMux I__7889 (
            .O(N__40249),
            .I(N__40241));
    InMux I__7888 (
            .O(N__40246),
            .I(N__40238));
    LocalMux I__7887 (
            .O(N__40241),
            .I(N__40235));
    LocalMux I__7886 (
            .O(N__40238),
            .I(N__40230));
    Span4Mux_v I__7885 (
            .O(N__40235),
            .I(N__40230));
    Odrv4 I__7884 (
            .O(N__40230),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__7883 (
            .O(N__40227),
            .I(N__40222));
    InMux I__7882 (
            .O(N__40226),
            .I(N__40217));
    InMux I__7881 (
            .O(N__40225),
            .I(N__40217));
    LocalMux I__7880 (
            .O(N__40222),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    LocalMux I__7879 (
            .O(N__40217),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__7878 (
            .O(N__40212),
            .I(N__40209));
    LocalMux I__7877 (
            .O(N__40209),
            .I(\ppm_encoder_1.N_295 ));
    InMux I__7876 (
            .O(N__40206),
            .I(N__40199));
    InMux I__7875 (
            .O(N__40205),
            .I(N__40199));
    InMux I__7874 (
            .O(N__40204),
            .I(N__40196));
    LocalMux I__7873 (
            .O(N__40199),
            .I(N__40193));
    LocalMux I__7872 (
            .O(N__40196),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv12 I__7871 (
            .O(N__40193),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__7870 (
            .O(N__40188),
            .I(N__40185));
    LocalMux I__7869 (
            .O(N__40185),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ));
    CascadeMux I__7868 (
            .O(N__40182),
            .I(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ));
    InMux I__7867 (
            .O(N__40179),
            .I(N__40176));
    LocalMux I__7866 (
            .O(N__40176),
            .I(\ppm_encoder_1.un2_throttle_iv_1_6 ));
    InMux I__7865 (
            .O(N__40173),
            .I(N__40166));
    InMux I__7864 (
            .O(N__40172),
            .I(N__40166));
    CascadeMux I__7863 (
            .O(N__40171),
            .I(N__40163));
    LocalMux I__7862 (
            .O(N__40166),
            .I(N__40160));
    InMux I__7861 (
            .O(N__40163),
            .I(N__40157));
    Span4Mux_h I__7860 (
            .O(N__40160),
            .I(N__40154));
    LocalMux I__7859 (
            .O(N__40157),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv4 I__7858 (
            .O(N__40154),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    CascadeMux I__7857 (
            .O(N__40149),
            .I(N__40145));
    CascadeMux I__7856 (
            .O(N__40148),
            .I(N__40141));
    InMux I__7855 (
            .O(N__40145),
            .I(N__40138));
    InMux I__7854 (
            .O(N__40144),
            .I(N__40133));
    InMux I__7853 (
            .O(N__40141),
            .I(N__40133));
    LocalMux I__7852 (
            .O(N__40138),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    LocalMux I__7851 (
            .O(N__40133),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    CascadeMux I__7850 (
            .O(N__40128),
            .I(\ppm_encoder_1.N_292_cascade_ ));
    InMux I__7849 (
            .O(N__40125),
            .I(N__40122));
    LocalMux I__7848 (
            .O(N__40122),
            .I(N__40119));
    Span4Mux_h I__7847 (
            .O(N__40119),
            .I(N__40116));
    Odrv4 I__7846 (
            .O(N__40116),
            .I(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ));
    InMux I__7845 (
            .O(N__40113),
            .I(N__40104));
    InMux I__7844 (
            .O(N__40112),
            .I(N__40104));
    InMux I__7843 (
            .O(N__40111),
            .I(N__40104));
    LocalMux I__7842 (
            .O(N__40104),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    InMux I__7841 (
            .O(N__40101),
            .I(N__40094));
    InMux I__7840 (
            .O(N__40100),
            .I(N__40094));
    InMux I__7839 (
            .O(N__40099),
            .I(N__40091));
    LocalMux I__7838 (
            .O(N__40094),
            .I(N__40088));
    LocalMux I__7837 (
            .O(N__40091),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    Odrv4 I__7836 (
            .O(N__40088),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    CascadeMux I__7835 (
            .O(N__40083),
            .I(\ppm_encoder_1.N_297_cascade_ ));
    InMux I__7834 (
            .O(N__40080),
            .I(N__40077));
    LocalMux I__7833 (
            .O(N__40077),
            .I(N__40074));
    Span4Mux_h I__7832 (
            .O(N__40074),
            .I(N__40071));
    Span4Mux_v I__7831 (
            .O(N__40071),
            .I(N__40068));
    Odrv4 I__7830 (
            .O(N__40068),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__7829 (
            .O(N__40065),
            .I(N__40056));
    InMux I__7828 (
            .O(N__40064),
            .I(N__40056));
    InMux I__7827 (
            .O(N__40063),
            .I(N__40056));
    LocalMux I__7826 (
            .O(N__40056),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    InMux I__7825 (
            .O(N__40053),
            .I(N__40050));
    LocalMux I__7824 (
            .O(N__40050),
            .I(N__40047));
    Span4Mux_v I__7823 (
            .O(N__40047),
            .I(N__40042));
    InMux I__7822 (
            .O(N__40046),
            .I(N__40039));
    CascadeMux I__7821 (
            .O(N__40045),
            .I(N__40036));
    Span4Mux_h I__7820 (
            .O(N__40042),
            .I(N__40033));
    LocalMux I__7819 (
            .O(N__40039),
            .I(N__40030));
    InMux I__7818 (
            .O(N__40036),
            .I(N__40027));
    Sp12to4 I__7817 (
            .O(N__40033),
            .I(N__40022));
    Span12Mux_v I__7816 (
            .O(N__40030),
            .I(N__40022));
    LocalMux I__7815 (
            .O(N__40027),
            .I(throttle_order_11));
    Odrv12 I__7814 (
            .O(N__40022),
            .I(throttle_order_11));
    InMux I__7813 (
            .O(N__40017),
            .I(N__40014));
    LocalMux I__7812 (
            .O(N__40014),
            .I(N__40011));
    Span4Mux_v I__7811 (
            .O(N__40011),
            .I(N__40008));
    Odrv4 I__7810 (
            .O(N__40008),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    CascadeMux I__7809 (
            .O(N__40005),
            .I(N__40002));
    InMux I__7808 (
            .O(N__40002),
            .I(N__39997));
    InMux I__7807 (
            .O(N__40001),
            .I(N__39992));
    InMux I__7806 (
            .O(N__40000),
            .I(N__39992));
    LocalMux I__7805 (
            .O(N__39997),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    LocalMux I__7804 (
            .O(N__39992),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    CascadeMux I__7803 (
            .O(N__39987),
            .I(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ));
    CascadeMux I__7802 (
            .O(N__39984),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ));
    InMux I__7801 (
            .O(N__39981),
            .I(N__39975));
    InMux I__7800 (
            .O(N__39980),
            .I(N__39975));
    LocalMux I__7799 (
            .O(N__39975),
            .I(N__39971));
    InMux I__7798 (
            .O(N__39974),
            .I(N__39968));
    Span4Mux_h I__7797 (
            .O(N__39971),
            .I(N__39965));
    LocalMux I__7796 (
            .O(N__39968),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    Odrv4 I__7795 (
            .O(N__39965),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    InMux I__7794 (
            .O(N__39960),
            .I(N__39957));
    LocalMux I__7793 (
            .O(N__39957),
            .I(\ppm_encoder_1.un2_throttle_iv_1_9 ));
    InMux I__7792 (
            .O(N__39954),
            .I(N__39947));
    InMux I__7791 (
            .O(N__39953),
            .I(N__39947));
    CascadeMux I__7790 (
            .O(N__39952),
            .I(N__39944));
    LocalMux I__7789 (
            .O(N__39947),
            .I(N__39941));
    InMux I__7788 (
            .O(N__39944),
            .I(N__39938));
    Span4Mux_h I__7787 (
            .O(N__39941),
            .I(N__39935));
    LocalMux I__7786 (
            .O(N__39938),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    Odrv4 I__7785 (
            .O(N__39935),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    CascadeMux I__7784 (
            .O(N__39930),
            .I(\ppm_encoder_1.N_298_cascade_ ));
    CascadeMux I__7783 (
            .O(N__39927),
            .I(N__39924));
    InMux I__7782 (
            .O(N__39924),
            .I(N__39921));
    LocalMux I__7781 (
            .O(N__39921),
            .I(N__39918));
    Span4Mux_h I__7780 (
            .O(N__39918),
            .I(N__39915));
    Span4Mux_v I__7779 (
            .O(N__39915),
            .I(N__39912));
    Odrv4 I__7778 (
            .O(N__39912),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__7777 (
            .O(N__39909),
            .I(N__39900));
    InMux I__7776 (
            .O(N__39908),
            .I(N__39900));
    InMux I__7775 (
            .O(N__39907),
            .I(N__39900));
    LocalMux I__7774 (
            .O(N__39900),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    InMux I__7773 (
            .O(N__39897),
            .I(N__39894));
    LocalMux I__7772 (
            .O(N__39894),
            .I(N__39891));
    Span4Mux_h I__7771 (
            .O(N__39891),
            .I(N__39887));
    InMux I__7770 (
            .O(N__39890),
            .I(N__39884));
    Sp12to4 I__7769 (
            .O(N__39887),
            .I(N__39879));
    LocalMux I__7768 (
            .O(N__39884),
            .I(N__39879));
    Span12Mux_v I__7767 (
            .O(N__39879),
            .I(N__39876));
    Odrv12 I__7766 (
            .O(N__39876),
            .I(front_order_12));
    InMux I__7765 (
            .O(N__39873),
            .I(N__39870));
    LocalMux I__7764 (
            .O(N__39870),
            .I(N__39867));
    Span4Mux_v I__7763 (
            .O(N__39867),
            .I(N__39864));
    Odrv4 I__7762 (
            .O(N__39864),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__7761 (
            .O(N__39861),
            .I(N__39852));
    InMux I__7760 (
            .O(N__39860),
            .I(N__39852));
    InMux I__7759 (
            .O(N__39859),
            .I(N__39852));
    LocalMux I__7758 (
            .O(N__39852),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    CascadeMux I__7757 (
            .O(N__39849),
            .I(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ));
    InMux I__7756 (
            .O(N__39846),
            .I(N__39843));
    LocalMux I__7755 (
            .O(N__39843),
            .I(\ppm_encoder_1.un2_throttle_iv_1_11 ));
    CEMux I__7754 (
            .O(N__39840),
            .I(N__39837));
    LocalMux I__7753 (
            .O(N__39837),
            .I(N__39834));
    Odrv4 I__7752 (
            .O(N__39834),
            .I(\pid_alt.state_1_0_0 ));
    InMux I__7751 (
            .O(N__39831),
            .I(N__39827));
    InMux I__7750 (
            .O(N__39830),
            .I(N__39824));
    LocalMux I__7749 (
            .O(N__39827),
            .I(N__39821));
    LocalMux I__7748 (
            .O(N__39824),
            .I(N__39818));
    Odrv4 I__7747 (
            .O(N__39821),
            .I(scaler_4_data_9));
    Odrv4 I__7746 (
            .O(N__39818),
            .I(scaler_4_data_9));
    InMux I__7745 (
            .O(N__39813),
            .I(N__39810));
    LocalMux I__7744 (
            .O(N__39810),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__7743 (
            .O(N__39807),
            .I(N__39804));
    LocalMux I__7742 (
            .O(N__39804),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__7741 (
            .O(N__39801),
            .I(N__39797));
    InMux I__7740 (
            .O(N__39800),
            .I(N__39794));
    LocalMux I__7739 (
            .O(N__39797),
            .I(N__39791));
    LocalMux I__7738 (
            .O(N__39794),
            .I(N__39788));
    Odrv4 I__7737 (
            .O(N__39791),
            .I(scaler_4_data_8));
    Odrv4 I__7736 (
            .O(N__39788),
            .I(scaler_4_data_8));
    InMux I__7735 (
            .O(N__39783),
            .I(N__39779));
    InMux I__7734 (
            .O(N__39782),
            .I(N__39776));
    LocalMux I__7733 (
            .O(N__39779),
            .I(N__39771));
    LocalMux I__7732 (
            .O(N__39776),
            .I(N__39771));
    Odrv4 I__7731 (
            .O(N__39771),
            .I(scaler_4_data_10));
    InMux I__7730 (
            .O(N__39768),
            .I(N__39765));
    LocalMux I__7729 (
            .O(N__39765),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    InMux I__7728 (
            .O(N__39762),
            .I(N__39758));
    InMux I__7727 (
            .O(N__39761),
            .I(N__39755));
    LocalMux I__7726 (
            .O(N__39758),
            .I(N__39752));
    LocalMux I__7725 (
            .O(N__39755),
            .I(N__39749));
    Odrv4 I__7724 (
            .O(N__39752),
            .I(scaler_4_data_13));
    Odrv4 I__7723 (
            .O(N__39749),
            .I(scaler_4_data_13));
    InMux I__7722 (
            .O(N__39744),
            .I(N__39741));
    LocalMux I__7721 (
            .O(N__39741),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    CascadeMux I__7720 (
            .O(N__39738),
            .I(N__39732));
    InMux I__7719 (
            .O(N__39737),
            .I(N__39706));
    InMux I__7718 (
            .O(N__39736),
            .I(N__39706));
    InMux I__7717 (
            .O(N__39735),
            .I(N__39706));
    InMux I__7716 (
            .O(N__39732),
            .I(N__39706));
    InMux I__7715 (
            .O(N__39731),
            .I(N__39706));
    InMux I__7714 (
            .O(N__39730),
            .I(N__39701));
    InMux I__7713 (
            .O(N__39729),
            .I(N__39701));
    InMux I__7712 (
            .O(N__39728),
            .I(N__39686));
    InMux I__7711 (
            .O(N__39727),
            .I(N__39686));
    InMux I__7710 (
            .O(N__39726),
            .I(N__39686));
    InMux I__7709 (
            .O(N__39725),
            .I(N__39686));
    InMux I__7708 (
            .O(N__39724),
            .I(N__39686));
    InMux I__7707 (
            .O(N__39723),
            .I(N__39686));
    InMux I__7706 (
            .O(N__39722),
            .I(N__39686));
    InMux I__7705 (
            .O(N__39721),
            .I(N__39679));
    InMux I__7704 (
            .O(N__39720),
            .I(N__39679));
    InMux I__7703 (
            .O(N__39719),
            .I(N__39679));
    InMux I__7702 (
            .O(N__39718),
            .I(N__39672));
    InMux I__7701 (
            .O(N__39717),
            .I(N__39669));
    LocalMux I__7700 (
            .O(N__39706),
            .I(N__39666));
    LocalMux I__7699 (
            .O(N__39701),
            .I(N__39659));
    LocalMux I__7698 (
            .O(N__39686),
            .I(N__39659));
    LocalMux I__7697 (
            .O(N__39679),
            .I(N__39659));
    InMux I__7696 (
            .O(N__39678),
            .I(N__39656));
    InMux I__7695 (
            .O(N__39677),
            .I(N__39653));
    InMux I__7694 (
            .O(N__39676),
            .I(N__39650));
    InMux I__7693 (
            .O(N__39675),
            .I(N__39647));
    LocalMux I__7692 (
            .O(N__39672),
            .I(N__39642));
    LocalMux I__7691 (
            .O(N__39669),
            .I(N__39642));
    Span4Mux_v I__7690 (
            .O(N__39666),
            .I(N__39635));
    Span4Mux_v I__7689 (
            .O(N__39659),
            .I(N__39635));
    LocalMux I__7688 (
            .O(N__39656),
            .I(N__39635));
    LocalMux I__7687 (
            .O(N__39653),
            .I(N__39632));
    LocalMux I__7686 (
            .O(N__39650),
            .I(N__39629));
    LocalMux I__7685 (
            .O(N__39647),
            .I(N__39626));
    Span4Mux_v I__7684 (
            .O(N__39642),
            .I(N__39623));
    Span4Mux_h I__7683 (
            .O(N__39635),
            .I(N__39618));
    Span4Mux_h I__7682 (
            .O(N__39632),
            .I(N__39618));
    Span4Mux_v I__7681 (
            .O(N__39629),
            .I(N__39615));
    Span12Mux_h I__7680 (
            .O(N__39626),
            .I(N__39612));
    Span4Mux_v I__7679 (
            .O(N__39623),
            .I(N__39607));
    Span4Mux_h I__7678 (
            .O(N__39618),
            .I(N__39607));
    Odrv4 I__7677 (
            .O(N__39615),
            .I(\pid_alt.N_72_i ));
    Odrv12 I__7676 (
            .O(N__39612),
            .I(\pid_alt.N_72_i ));
    Odrv4 I__7675 (
            .O(N__39607),
            .I(\pid_alt.N_72_i ));
    InMux I__7674 (
            .O(N__39600),
            .I(N__39596));
    InMux I__7673 (
            .O(N__39599),
            .I(N__39592));
    LocalMux I__7672 (
            .O(N__39596),
            .I(N__39589));
    CascadeMux I__7671 (
            .O(N__39595),
            .I(N__39585));
    LocalMux I__7670 (
            .O(N__39592),
            .I(N__39581));
    Sp12to4 I__7669 (
            .O(N__39589),
            .I(N__39578));
    InMux I__7668 (
            .O(N__39588),
            .I(N__39575));
    InMux I__7667 (
            .O(N__39585),
            .I(N__39572));
    InMux I__7666 (
            .O(N__39584),
            .I(N__39569));
    Sp12to4 I__7665 (
            .O(N__39581),
            .I(N__39564));
    Span12Mux_s9_v I__7664 (
            .O(N__39578),
            .I(N__39564));
    LocalMux I__7663 (
            .O(N__39575),
            .I(N__39559));
    LocalMux I__7662 (
            .O(N__39572),
            .I(N__39559));
    LocalMux I__7661 (
            .O(N__39569),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv12 I__7660 (
            .O(N__39564),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__7659 (
            .O(N__39559),
            .I(\pid_alt.stateZ0Z_0 ));
    CascadeMux I__7658 (
            .O(N__39552),
            .I(N__39548));
    InMux I__7657 (
            .O(N__39551),
            .I(N__39545));
    InMux I__7656 (
            .O(N__39548),
            .I(N__39542));
    LocalMux I__7655 (
            .O(N__39545),
            .I(N__39537));
    LocalMux I__7654 (
            .O(N__39542),
            .I(N__39537));
    Odrv4 I__7653 (
            .O(N__39537),
            .I(scaler_4_data_11));
    InMux I__7652 (
            .O(N__39534),
            .I(N__39531));
    LocalMux I__7651 (
            .O(N__39531),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__7650 (
            .O(N__39528),
            .I(N__39524));
    InMux I__7649 (
            .O(N__39527),
            .I(N__39521));
    LocalMux I__7648 (
            .O(N__39524),
            .I(N__39518));
    LocalMux I__7647 (
            .O(N__39521),
            .I(scaler_4_data_12));
    Odrv4 I__7646 (
            .O(N__39518),
            .I(scaler_4_data_12));
    InMux I__7645 (
            .O(N__39513),
            .I(N__39510));
    LocalMux I__7644 (
            .O(N__39510),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__7643 (
            .O(N__39507),
            .I(N__39504));
    LocalMux I__7642 (
            .O(N__39504),
            .I(N__39501));
    Odrv12 I__7641 (
            .O(N__39501),
            .I(drone_H_disp_front_i_13));
    InMux I__7640 (
            .O(N__39498),
            .I(N__39495));
    LocalMux I__7639 (
            .O(N__39495),
            .I(N__39491));
    InMux I__7638 (
            .O(N__39494),
            .I(N__39488));
    Span4Mux_s2_h I__7637 (
            .O(N__39491),
            .I(N__39485));
    LocalMux I__7636 (
            .O(N__39488),
            .I(N__39482));
    Span4Mux_v I__7635 (
            .O(N__39485),
            .I(N__39479));
    Span4Mux_s3_h I__7634 (
            .O(N__39482),
            .I(N__39476));
    Span4Mux_h I__7633 (
            .O(N__39479),
            .I(N__39473));
    Span4Mux_h I__7632 (
            .O(N__39476),
            .I(N__39470));
    Span4Mux_h I__7631 (
            .O(N__39473),
            .I(N__39467));
    Span4Mux_h I__7630 (
            .O(N__39470),
            .I(N__39462));
    Span4Mux_h I__7629 (
            .O(N__39467),
            .I(N__39462));
    Odrv4 I__7628 (
            .O(N__39462),
            .I(\pid_front.error_14 ));
    InMux I__7627 (
            .O(N__39459),
            .I(\pid_front.error_cry_9 ));
    InMux I__7626 (
            .O(N__39456),
            .I(\pid_front.error_cry_10 ));
    InMux I__7625 (
            .O(N__39453),
            .I(N__39449));
    InMux I__7624 (
            .O(N__39452),
            .I(N__39446));
    LocalMux I__7623 (
            .O(N__39449),
            .I(N__39443));
    LocalMux I__7622 (
            .O(N__39446),
            .I(N__39440));
    Span4Mux_s2_h I__7621 (
            .O(N__39443),
            .I(N__39437));
    Span4Mux_s3_h I__7620 (
            .O(N__39440),
            .I(N__39434));
    Sp12to4 I__7619 (
            .O(N__39437),
            .I(N__39431));
    Span4Mux_h I__7618 (
            .O(N__39434),
            .I(N__39428));
    Span12Mux_v I__7617 (
            .O(N__39431),
            .I(N__39425));
    Span4Mux_h I__7616 (
            .O(N__39428),
            .I(N__39422));
    Odrv12 I__7615 (
            .O(N__39425),
            .I(\pid_front.error_15 ));
    Odrv4 I__7614 (
            .O(N__39422),
            .I(\pid_front.error_15 ));
    InMux I__7613 (
            .O(N__39417),
            .I(N__39414));
    LocalMux I__7612 (
            .O(N__39414),
            .I(\dron_frame_decoder_1.drone_H_disp_front_10 ));
    InMux I__7611 (
            .O(N__39411),
            .I(N__39405));
    InMux I__7610 (
            .O(N__39410),
            .I(N__39405));
    LocalMux I__7609 (
            .O(N__39405),
            .I(drone_H_disp_front_11));
    CascadeMux I__7608 (
            .O(N__39402),
            .I(N__39399));
    InMux I__7607 (
            .O(N__39399),
            .I(N__39394));
    InMux I__7606 (
            .O(N__39398),
            .I(N__39389));
    InMux I__7605 (
            .O(N__39397),
            .I(N__39389));
    LocalMux I__7604 (
            .O(N__39394),
            .I(drone_H_disp_front_12));
    LocalMux I__7603 (
            .O(N__39389),
            .I(drone_H_disp_front_12));
    CascadeMux I__7602 (
            .O(N__39384),
            .I(N__39380));
    InMux I__7601 (
            .O(N__39383),
            .I(N__39375));
    InMux I__7600 (
            .O(N__39380),
            .I(N__39375));
    LocalMux I__7599 (
            .O(N__39375),
            .I(N__39372));
    Odrv4 I__7598 (
            .O(N__39372),
            .I(drone_H_disp_front_14));
    InMux I__7597 (
            .O(N__39369),
            .I(N__39366));
    LocalMux I__7596 (
            .O(N__39366),
            .I(N__39363));
    Odrv4 I__7595 (
            .O(N__39363),
            .I(drone_H_disp_front_15));
    InMux I__7594 (
            .O(N__39360),
            .I(N__39357));
    LocalMux I__7593 (
            .O(N__39357),
            .I(N__39354));
    Odrv12 I__7592 (
            .O(N__39354),
            .I(\dron_frame_decoder_1.drone_H_disp_front_8 ));
    IoInMux I__7591 (
            .O(N__39351),
            .I(N__39348));
    LocalMux I__7590 (
            .O(N__39348),
            .I(N__39345));
    Odrv4 I__7589 (
            .O(N__39345),
            .I(\pid_alt.state_0_0 ));
    InMux I__7588 (
            .O(N__39342),
            .I(N__39339));
    LocalMux I__7587 (
            .O(N__39339),
            .I(drone_H_disp_front_i_6));
    CascadeMux I__7586 (
            .O(N__39336),
            .I(N__39333));
    InMux I__7585 (
            .O(N__39333),
            .I(N__39330));
    LocalMux I__7584 (
            .O(N__39330),
            .I(front_command_2));
    InMux I__7583 (
            .O(N__39327),
            .I(N__39323));
    InMux I__7582 (
            .O(N__39326),
            .I(N__39320));
    LocalMux I__7581 (
            .O(N__39323),
            .I(N__39317));
    LocalMux I__7580 (
            .O(N__39320),
            .I(N__39314));
    Span4Mux_s3_h I__7579 (
            .O(N__39317),
            .I(N__39311));
    Span12Mux_s1_h I__7578 (
            .O(N__39314),
            .I(N__39308));
    Span4Mux_h I__7577 (
            .O(N__39311),
            .I(N__39305));
    Span12Mux_h I__7576 (
            .O(N__39308),
            .I(N__39302));
    Span4Mux_h I__7575 (
            .O(N__39305),
            .I(N__39299));
    Odrv12 I__7574 (
            .O(N__39302),
            .I(\pid_front.error_6 ));
    Odrv4 I__7573 (
            .O(N__39299),
            .I(\pid_front.error_6 ));
    InMux I__7572 (
            .O(N__39294),
            .I(\pid_front.error_cry_1_0 ));
    InMux I__7571 (
            .O(N__39291),
            .I(N__39288));
    LocalMux I__7570 (
            .O(N__39288),
            .I(N__39285));
    Span4Mux_v I__7569 (
            .O(N__39285),
            .I(N__39282));
    Odrv4 I__7568 (
            .O(N__39282),
            .I(drone_H_disp_front_i_7));
    CascadeMux I__7567 (
            .O(N__39279),
            .I(N__39276));
    InMux I__7566 (
            .O(N__39276),
            .I(N__39273));
    LocalMux I__7565 (
            .O(N__39273),
            .I(front_command_3));
    InMux I__7564 (
            .O(N__39270),
            .I(N__39267));
    LocalMux I__7563 (
            .O(N__39267),
            .I(N__39263));
    InMux I__7562 (
            .O(N__39266),
            .I(N__39260));
    Span4Mux_v I__7561 (
            .O(N__39263),
            .I(N__39257));
    LocalMux I__7560 (
            .O(N__39260),
            .I(N__39254));
    Span4Mux_h I__7559 (
            .O(N__39257),
            .I(N__39251));
    Span4Mux_s3_h I__7558 (
            .O(N__39254),
            .I(N__39248));
    Span4Mux_h I__7557 (
            .O(N__39251),
            .I(N__39245));
    Span4Mux_h I__7556 (
            .O(N__39248),
            .I(N__39242));
    Span4Mux_h I__7555 (
            .O(N__39245),
            .I(N__39239));
    Span4Mux_h I__7554 (
            .O(N__39242),
            .I(N__39236));
    Odrv4 I__7553 (
            .O(N__39239),
            .I(\pid_front.error_7 ));
    Odrv4 I__7552 (
            .O(N__39236),
            .I(\pid_front.error_7 ));
    InMux I__7551 (
            .O(N__39231),
            .I(\pid_front.error_cry_2_0 ));
    InMux I__7550 (
            .O(N__39228),
            .I(N__39225));
    LocalMux I__7549 (
            .O(N__39225),
            .I(N__39222));
    Odrv4 I__7548 (
            .O(N__39222),
            .I(drone_H_disp_front_i_8));
    CascadeMux I__7547 (
            .O(N__39219),
            .I(N__39216));
    InMux I__7546 (
            .O(N__39216),
            .I(N__39213));
    LocalMux I__7545 (
            .O(N__39213),
            .I(front_command_4));
    InMux I__7544 (
            .O(N__39210),
            .I(N__39207));
    LocalMux I__7543 (
            .O(N__39207),
            .I(N__39203));
    InMux I__7542 (
            .O(N__39206),
            .I(N__39200));
    Span4Mux_v I__7541 (
            .O(N__39203),
            .I(N__39197));
    LocalMux I__7540 (
            .O(N__39200),
            .I(N__39194));
    Span4Mux_h I__7539 (
            .O(N__39197),
            .I(N__39191));
    Span4Mux_s3_h I__7538 (
            .O(N__39194),
            .I(N__39188));
    Span4Mux_h I__7537 (
            .O(N__39191),
            .I(N__39185));
    Span4Mux_h I__7536 (
            .O(N__39188),
            .I(N__39182));
    Span4Mux_h I__7535 (
            .O(N__39185),
            .I(N__39179));
    Span4Mux_h I__7534 (
            .O(N__39182),
            .I(N__39176));
    Odrv4 I__7533 (
            .O(N__39179),
            .I(\pid_front.error_8 ));
    Odrv4 I__7532 (
            .O(N__39176),
            .I(\pid_front.error_8 ));
    InMux I__7531 (
            .O(N__39171),
            .I(bfn_13_24_0_));
    CascadeMux I__7530 (
            .O(N__39168),
            .I(N__39165));
    InMux I__7529 (
            .O(N__39165),
            .I(N__39162));
    LocalMux I__7528 (
            .O(N__39162),
            .I(front_command_5));
    InMux I__7527 (
            .O(N__39159),
            .I(N__39156));
    LocalMux I__7526 (
            .O(N__39156),
            .I(N__39152));
    InMux I__7525 (
            .O(N__39155),
            .I(N__39149));
    Span4Mux_v I__7524 (
            .O(N__39152),
            .I(N__39146));
    LocalMux I__7523 (
            .O(N__39149),
            .I(N__39143));
    Span4Mux_h I__7522 (
            .O(N__39146),
            .I(N__39140));
    Span4Mux_s3_h I__7521 (
            .O(N__39143),
            .I(N__39137));
    Span4Mux_h I__7520 (
            .O(N__39140),
            .I(N__39134));
    Span4Mux_h I__7519 (
            .O(N__39137),
            .I(N__39131));
    Span4Mux_h I__7518 (
            .O(N__39134),
            .I(N__39128));
    Span4Mux_h I__7517 (
            .O(N__39131),
            .I(N__39125));
    Odrv4 I__7516 (
            .O(N__39128),
            .I(\pid_front.error_9 ));
    Odrv4 I__7515 (
            .O(N__39125),
            .I(\pid_front.error_9 ));
    InMux I__7514 (
            .O(N__39120),
            .I(\pid_front.error_cry_4 ));
    InMux I__7513 (
            .O(N__39117),
            .I(N__39114));
    LocalMux I__7512 (
            .O(N__39114),
            .I(drone_H_disp_front_i_10));
    CascadeMux I__7511 (
            .O(N__39111),
            .I(N__39108));
    InMux I__7510 (
            .O(N__39108),
            .I(N__39105));
    LocalMux I__7509 (
            .O(N__39105),
            .I(N__39102));
    Odrv4 I__7508 (
            .O(N__39102),
            .I(front_command_6));
    InMux I__7507 (
            .O(N__39099),
            .I(N__39096));
    LocalMux I__7506 (
            .O(N__39096),
            .I(N__39092));
    InMux I__7505 (
            .O(N__39095),
            .I(N__39089));
    Span4Mux_v I__7504 (
            .O(N__39092),
            .I(N__39086));
    LocalMux I__7503 (
            .O(N__39089),
            .I(N__39083));
    Span4Mux_h I__7502 (
            .O(N__39086),
            .I(N__39080));
    Span4Mux_s3_h I__7501 (
            .O(N__39083),
            .I(N__39077));
    Span4Mux_h I__7500 (
            .O(N__39080),
            .I(N__39074));
    Span4Mux_h I__7499 (
            .O(N__39077),
            .I(N__39071));
    Span4Mux_h I__7498 (
            .O(N__39074),
            .I(N__39068));
    Span4Mux_h I__7497 (
            .O(N__39071),
            .I(N__39065));
    Odrv4 I__7496 (
            .O(N__39068),
            .I(\pid_front.error_10 ));
    Odrv4 I__7495 (
            .O(N__39065),
            .I(\pid_front.error_10 ));
    InMux I__7494 (
            .O(N__39060),
            .I(\pid_front.error_cry_5 ));
    InMux I__7493 (
            .O(N__39057),
            .I(N__39054));
    LocalMux I__7492 (
            .O(N__39054),
            .I(\pid_front.error_axbZ0Z_7 ));
    InMux I__7491 (
            .O(N__39051),
            .I(N__39048));
    LocalMux I__7490 (
            .O(N__39048),
            .I(N__39044));
    InMux I__7489 (
            .O(N__39047),
            .I(N__39041));
    Span4Mux_v I__7488 (
            .O(N__39044),
            .I(N__39038));
    LocalMux I__7487 (
            .O(N__39041),
            .I(N__39035));
    Span4Mux_h I__7486 (
            .O(N__39038),
            .I(N__39032));
    Span4Mux_s3_h I__7485 (
            .O(N__39035),
            .I(N__39029));
    Span4Mux_h I__7484 (
            .O(N__39032),
            .I(N__39026));
    Span4Mux_h I__7483 (
            .O(N__39029),
            .I(N__39023));
    Span4Mux_h I__7482 (
            .O(N__39026),
            .I(N__39020));
    Span4Mux_h I__7481 (
            .O(N__39023),
            .I(N__39017));
    Odrv4 I__7480 (
            .O(N__39020),
            .I(\pid_front.error_11 ));
    Odrv4 I__7479 (
            .O(N__39017),
            .I(\pid_front.error_11 ));
    InMux I__7478 (
            .O(N__39012),
            .I(\pid_front.error_cry_6 ));
    InMux I__7477 (
            .O(N__39009),
            .I(N__39006));
    LocalMux I__7476 (
            .O(N__39006),
            .I(\pid_front.error_axb_8_l_ofx_0 ));
    InMux I__7475 (
            .O(N__39003),
            .I(N__39000));
    LocalMux I__7474 (
            .O(N__39000),
            .I(N__38997));
    Span4Mux_v I__7473 (
            .O(N__38997),
            .I(N__38994));
    Span4Mux_h I__7472 (
            .O(N__38994),
            .I(N__38990));
    InMux I__7471 (
            .O(N__38993),
            .I(N__38987));
    Span4Mux_h I__7470 (
            .O(N__38990),
            .I(N__38984));
    LocalMux I__7469 (
            .O(N__38987),
            .I(N__38981));
    Span4Mux_h I__7468 (
            .O(N__38984),
            .I(N__38978));
    Span12Mux_s6_v I__7467 (
            .O(N__38981),
            .I(N__38975));
    Odrv4 I__7466 (
            .O(N__38978),
            .I(\pid_front.error_12 ));
    Odrv12 I__7465 (
            .O(N__38975),
            .I(\pid_front.error_12 ));
    InMux I__7464 (
            .O(N__38970),
            .I(\pid_front.error_cry_7 ));
    InMux I__7463 (
            .O(N__38967),
            .I(N__38964));
    LocalMux I__7462 (
            .O(N__38964),
            .I(drone_H_disp_front_i_12));
    InMux I__7461 (
            .O(N__38961),
            .I(N__38957));
    InMux I__7460 (
            .O(N__38960),
            .I(N__38954));
    LocalMux I__7459 (
            .O(N__38957),
            .I(N__38951));
    LocalMux I__7458 (
            .O(N__38954),
            .I(N__38948));
    Span4Mux_v I__7457 (
            .O(N__38951),
            .I(N__38945));
    Span12Mux_s1_h I__7456 (
            .O(N__38948),
            .I(N__38942));
    Span4Mux_h I__7455 (
            .O(N__38945),
            .I(N__38939));
    Span12Mux_h I__7454 (
            .O(N__38942),
            .I(N__38936));
    Span4Mux_h I__7453 (
            .O(N__38939),
            .I(N__38933));
    Odrv12 I__7452 (
            .O(N__38936),
            .I(\pid_front.error_13 ));
    Odrv4 I__7451 (
            .O(N__38933),
            .I(\pid_front.error_13 ));
    InMux I__7450 (
            .O(N__38928),
            .I(\pid_front.error_cry_8 ));
    InMux I__7449 (
            .O(N__38925),
            .I(N__38922));
    LocalMux I__7448 (
            .O(N__38922),
            .I(N__38919));
    Odrv4 I__7447 (
            .O(N__38919),
            .I(drone_H_disp_front_2));
    InMux I__7446 (
            .O(N__38916),
            .I(N__38913));
    LocalMux I__7445 (
            .O(N__38913),
            .I(N__38909));
    InMux I__7444 (
            .O(N__38912),
            .I(N__38906));
    Span4Mux_v I__7443 (
            .O(N__38909),
            .I(N__38903));
    LocalMux I__7442 (
            .O(N__38906),
            .I(N__38899));
    Span4Mux_h I__7441 (
            .O(N__38903),
            .I(N__38896));
    InMux I__7440 (
            .O(N__38902),
            .I(N__38893));
    Span12Mux_v I__7439 (
            .O(N__38899),
            .I(N__38890));
    Span4Mux_h I__7438 (
            .O(N__38896),
            .I(N__38887));
    LocalMux I__7437 (
            .O(N__38893),
            .I(N__38884));
    Span12Mux_h I__7436 (
            .O(N__38890),
            .I(N__38881));
    Span4Mux_h I__7435 (
            .O(N__38887),
            .I(N__38876));
    Span4Mux_v I__7434 (
            .O(N__38884),
            .I(N__38876));
    Odrv12 I__7433 (
            .O(N__38881),
            .I(drone_H_disp_front_0));
    Odrv4 I__7432 (
            .O(N__38876),
            .I(drone_H_disp_front_0));
    InMux I__7431 (
            .O(N__38871),
            .I(N__38868));
    LocalMux I__7430 (
            .O(N__38868),
            .I(\pid_front.error_axb_0 ));
    InMux I__7429 (
            .O(N__38865),
            .I(N__38862));
    LocalMux I__7428 (
            .O(N__38862),
            .I(N__38859));
    Span4Mux_v I__7427 (
            .O(N__38859),
            .I(N__38856));
    Odrv4 I__7426 (
            .O(N__38856),
            .I(\pid_front.error_axbZ0Z_1 ));
    InMux I__7425 (
            .O(N__38853),
            .I(N__38850));
    LocalMux I__7424 (
            .O(N__38850),
            .I(N__38846));
    InMux I__7423 (
            .O(N__38849),
            .I(N__38843));
    Span4Mux_s1_h I__7422 (
            .O(N__38846),
            .I(N__38840));
    LocalMux I__7421 (
            .O(N__38843),
            .I(N__38837));
    Span4Mux_v I__7420 (
            .O(N__38840),
            .I(N__38834));
    Span4Mux_s0_h I__7419 (
            .O(N__38837),
            .I(N__38831));
    Span4Mux_h I__7418 (
            .O(N__38834),
            .I(N__38828));
    Span4Mux_h I__7417 (
            .O(N__38831),
            .I(N__38825));
    Span4Mux_h I__7416 (
            .O(N__38828),
            .I(N__38822));
    Span4Mux_h I__7415 (
            .O(N__38825),
            .I(N__38819));
    Span4Mux_h I__7414 (
            .O(N__38822),
            .I(N__38814));
    Span4Mux_h I__7413 (
            .O(N__38819),
            .I(N__38814));
    Odrv4 I__7412 (
            .O(N__38814),
            .I(\pid_front.error_1 ));
    InMux I__7411 (
            .O(N__38811),
            .I(\pid_front.error_cry_0 ));
    InMux I__7410 (
            .O(N__38808),
            .I(N__38805));
    LocalMux I__7409 (
            .O(N__38805),
            .I(\pid_front.error_axbZ0Z_2 ));
    InMux I__7408 (
            .O(N__38802),
            .I(N__38799));
    LocalMux I__7407 (
            .O(N__38799),
            .I(N__38796));
    Span4Mux_v I__7406 (
            .O(N__38796),
            .I(N__38792));
    InMux I__7405 (
            .O(N__38795),
            .I(N__38789));
    Span4Mux_v I__7404 (
            .O(N__38792),
            .I(N__38786));
    LocalMux I__7403 (
            .O(N__38789),
            .I(N__38783));
    Span4Mux_h I__7402 (
            .O(N__38786),
            .I(N__38780));
    Span4Mux_v I__7401 (
            .O(N__38783),
            .I(N__38777));
    Span4Mux_h I__7400 (
            .O(N__38780),
            .I(N__38774));
    Span4Mux_h I__7399 (
            .O(N__38777),
            .I(N__38771));
    Span4Mux_h I__7398 (
            .O(N__38774),
            .I(N__38766));
    Span4Mux_h I__7397 (
            .O(N__38771),
            .I(N__38766));
    Odrv4 I__7396 (
            .O(N__38766),
            .I(\pid_front.error_2 ));
    InMux I__7395 (
            .O(N__38763),
            .I(\pid_front.error_cry_1 ));
    InMux I__7394 (
            .O(N__38760),
            .I(N__38757));
    LocalMux I__7393 (
            .O(N__38757),
            .I(N__38754));
    Odrv4 I__7392 (
            .O(N__38754),
            .I(\pid_front.error_axbZ0Z_3 ));
    InMux I__7391 (
            .O(N__38751),
            .I(N__38748));
    LocalMux I__7390 (
            .O(N__38748),
            .I(N__38744));
    InMux I__7389 (
            .O(N__38747),
            .I(N__38741));
    Span4Mux_v I__7388 (
            .O(N__38744),
            .I(N__38738));
    LocalMux I__7387 (
            .O(N__38741),
            .I(N__38735));
    Span4Mux_h I__7386 (
            .O(N__38738),
            .I(N__38732));
    Span4Mux_v I__7385 (
            .O(N__38735),
            .I(N__38729));
    Span4Mux_h I__7384 (
            .O(N__38732),
            .I(N__38726));
    Span4Mux_h I__7383 (
            .O(N__38729),
            .I(N__38723));
    Span4Mux_h I__7382 (
            .O(N__38726),
            .I(N__38720));
    Span4Mux_h I__7381 (
            .O(N__38723),
            .I(N__38717));
    Odrv4 I__7380 (
            .O(N__38720),
            .I(\pid_front.error_3 ));
    Odrv4 I__7379 (
            .O(N__38717),
            .I(\pid_front.error_3 ));
    InMux I__7378 (
            .O(N__38712),
            .I(\pid_front.error_cry_2 ));
    InMux I__7377 (
            .O(N__38709),
            .I(N__38706));
    LocalMux I__7376 (
            .O(N__38706),
            .I(drone_H_disp_front_i_4));
    CascadeMux I__7375 (
            .O(N__38703),
            .I(N__38700));
    InMux I__7374 (
            .O(N__38700),
            .I(N__38697));
    LocalMux I__7373 (
            .O(N__38697),
            .I(N__38694));
    Odrv4 I__7372 (
            .O(N__38694),
            .I(front_command_0));
    InMux I__7371 (
            .O(N__38691),
            .I(N__38688));
    LocalMux I__7370 (
            .O(N__38688),
            .I(N__38685));
    Span4Mux_s2_h I__7369 (
            .O(N__38685),
            .I(N__38681));
    InMux I__7368 (
            .O(N__38684),
            .I(N__38678));
    Span4Mux_v I__7367 (
            .O(N__38681),
            .I(N__38675));
    LocalMux I__7366 (
            .O(N__38678),
            .I(N__38672));
    Span4Mux_h I__7365 (
            .O(N__38675),
            .I(N__38669));
    Span4Mux_s3_h I__7364 (
            .O(N__38672),
            .I(N__38666));
    Span4Mux_h I__7363 (
            .O(N__38669),
            .I(N__38663));
    Span4Mux_h I__7362 (
            .O(N__38666),
            .I(N__38660));
    Span4Mux_h I__7361 (
            .O(N__38663),
            .I(N__38655));
    Span4Mux_h I__7360 (
            .O(N__38660),
            .I(N__38655));
    Odrv4 I__7359 (
            .O(N__38655),
            .I(\pid_front.error_4 ));
    InMux I__7358 (
            .O(N__38652),
            .I(\pid_front.error_cry_3 ));
    InMux I__7357 (
            .O(N__38649),
            .I(N__38646));
    LocalMux I__7356 (
            .O(N__38646),
            .I(drone_H_disp_front_i_5));
    CascadeMux I__7355 (
            .O(N__38643),
            .I(N__38640));
    InMux I__7354 (
            .O(N__38640),
            .I(N__38637));
    LocalMux I__7353 (
            .O(N__38637),
            .I(front_command_1));
    InMux I__7352 (
            .O(N__38634),
            .I(N__38631));
    LocalMux I__7351 (
            .O(N__38631),
            .I(N__38627));
    InMux I__7350 (
            .O(N__38630),
            .I(N__38624));
    Span4Mux_v I__7349 (
            .O(N__38627),
            .I(N__38621));
    LocalMux I__7348 (
            .O(N__38624),
            .I(N__38618));
    Span4Mux_h I__7347 (
            .O(N__38621),
            .I(N__38615));
    Span4Mux_v I__7346 (
            .O(N__38618),
            .I(N__38612));
    Span4Mux_h I__7345 (
            .O(N__38615),
            .I(N__38609));
    Span4Mux_h I__7344 (
            .O(N__38612),
            .I(N__38606));
    Span4Mux_h I__7343 (
            .O(N__38609),
            .I(N__38603));
    Span4Mux_h I__7342 (
            .O(N__38606),
            .I(N__38600));
    Odrv4 I__7341 (
            .O(N__38603),
            .I(\pid_front.error_5 ));
    Odrv4 I__7340 (
            .O(N__38600),
            .I(\pid_front.error_5 ));
    InMux I__7339 (
            .O(N__38595),
            .I(\pid_front.error_cry_0_0 ));
    CascadeMux I__7338 (
            .O(N__38592),
            .I(\pid_front.error_p_reg_esr_RNI6MF7Z0Z_1_cascade_ ));
    CascadeMux I__7337 (
            .O(N__38589),
            .I(N__38585));
    InMux I__7336 (
            .O(N__38588),
            .I(N__38582));
    InMux I__7335 (
            .O(N__38585),
            .I(N__38579));
    LocalMux I__7334 (
            .O(N__38582),
            .I(\pid_front.un1_pid_prereg ));
    LocalMux I__7333 (
            .O(N__38579),
            .I(\pid_front.un1_pid_prereg ));
    InMux I__7332 (
            .O(N__38574),
            .I(N__38571));
    LocalMux I__7331 (
            .O(N__38571),
            .I(drone_H_disp_front_3));
    InMux I__7330 (
            .O(N__38568),
            .I(N__38565));
    LocalMux I__7329 (
            .O(N__38565),
            .I(N__38561));
    InMux I__7328 (
            .O(N__38564),
            .I(N__38558));
    Odrv4 I__7327 (
            .O(N__38561),
            .I(\pid_front.error_p_reg_esr_RNI6MF7Z0Z_1 ));
    LocalMux I__7326 (
            .O(N__38558),
            .I(\pid_front.error_p_reg_esr_RNI6MF7Z0Z_1 ));
    InMux I__7325 (
            .O(N__38553),
            .I(N__38546));
    InMux I__7324 (
            .O(N__38552),
            .I(N__38546));
    InMux I__7323 (
            .O(N__38551),
            .I(N__38543));
    LocalMux I__7322 (
            .O(N__38546),
            .I(N__38540));
    LocalMux I__7321 (
            .O(N__38543),
            .I(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ));
    Odrv4 I__7320 (
            .O(N__38540),
            .I(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ));
    InMux I__7319 (
            .O(N__38535),
            .I(N__38532));
    LocalMux I__7318 (
            .O(N__38532),
            .I(\pid_front.error_p_reg_esr_RNIUQTFZ0Z_1 ));
    InMux I__7317 (
            .O(N__38529),
            .I(N__38524));
    InMux I__7316 (
            .O(N__38528),
            .I(N__38521));
    InMux I__7315 (
            .O(N__38527),
            .I(N__38518));
    LocalMux I__7314 (
            .O(N__38524),
            .I(N__38515));
    LocalMux I__7313 (
            .O(N__38521),
            .I(N__38512));
    LocalMux I__7312 (
            .O(N__38518),
            .I(N__38507));
    Span4Mux_v I__7311 (
            .O(N__38515),
            .I(N__38507));
    Span12Mux_v I__7310 (
            .O(N__38512),
            .I(N__38504));
    Span4Mux_v I__7309 (
            .O(N__38507),
            .I(N__38501));
    Span12Mux_h I__7308 (
            .O(N__38504),
            .I(N__38498));
    Span4Mux_v I__7307 (
            .O(N__38501),
            .I(N__38495));
    Odrv12 I__7306 (
            .O(N__38498),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    Odrv4 I__7305 (
            .O(N__38495),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    InMux I__7304 (
            .O(N__38490),
            .I(N__38487));
    LocalMux I__7303 (
            .O(N__38487),
            .I(N__38483));
    InMux I__7302 (
            .O(N__38486),
            .I(N__38480));
    Span4Mux_v I__7301 (
            .O(N__38483),
            .I(N__38477));
    LocalMux I__7300 (
            .O(N__38480),
            .I(N__38474));
    Span4Mux_h I__7299 (
            .O(N__38477),
            .I(N__38471));
    Span4Mux_v I__7298 (
            .O(N__38474),
            .I(N__38468));
    Span4Mux_h I__7297 (
            .O(N__38471),
            .I(N__38465));
    Span4Mux_v I__7296 (
            .O(N__38468),
            .I(N__38462));
    Odrv4 I__7295 (
            .O(N__38465),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    Odrv4 I__7294 (
            .O(N__38462),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    InMux I__7293 (
            .O(N__38457),
            .I(N__38454));
    LocalMux I__7292 (
            .O(N__38454),
            .I(N__38450));
    InMux I__7291 (
            .O(N__38453),
            .I(N__38447));
    Span12Mux_h I__7290 (
            .O(N__38450),
            .I(N__38444));
    LocalMux I__7289 (
            .O(N__38447),
            .I(N__38441));
    Span12Mux_v I__7288 (
            .O(N__38444),
            .I(N__38438));
    Span4Mux_v I__7287 (
            .O(N__38441),
            .I(N__38435));
    Odrv12 I__7286 (
            .O(N__38438),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    Odrv4 I__7285 (
            .O(N__38435),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    InMux I__7284 (
            .O(N__38430),
            .I(N__38424));
    InMux I__7283 (
            .O(N__38429),
            .I(N__38424));
    LocalMux I__7282 (
            .O(N__38424),
            .I(N__38421));
    Span12Mux_h I__7281 (
            .O(N__38421),
            .I(N__38418));
    Odrv12 I__7280 (
            .O(N__38418),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ));
    InMux I__7279 (
            .O(N__38415),
            .I(N__38412));
    LocalMux I__7278 (
            .O(N__38412),
            .I(N__38409));
    Odrv4 I__7277 (
            .O(N__38409),
            .I(\dron_frame_decoder_1.drone_H_disp_front_5 ));
    InMux I__7276 (
            .O(N__38406),
            .I(N__38403));
    LocalMux I__7275 (
            .O(N__38403),
            .I(N__38400));
    Odrv4 I__7274 (
            .O(N__38400),
            .I(\dron_frame_decoder_1.drone_H_disp_front_4 ));
    InMux I__7273 (
            .O(N__38397),
            .I(N__38393));
    InMux I__7272 (
            .O(N__38396),
            .I(N__38390));
    LocalMux I__7271 (
            .O(N__38393),
            .I(N__38387));
    LocalMux I__7270 (
            .O(N__38390),
            .I(N__38383));
    Span4Mux_h I__7269 (
            .O(N__38387),
            .I(N__38380));
    InMux I__7268 (
            .O(N__38386),
            .I(N__38377));
    Span4Mux_h I__7267 (
            .O(N__38383),
            .I(N__38374));
    Span4Mux_h I__7266 (
            .O(N__38380),
            .I(N__38371));
    LocalMux I__7265 (
            .O(N__38377),
            .I(N__38368));
    Span4Mux_h I__7264 (
            .O(N__38374),
            .I(N__38365));
    Span4Mux_v I__7263 (
            .O(N__38371),
            .I(N__38362));
    Span4Mux_h I__7262 (
            .O(N__38368),
            .I(N__38357));
    Span4Mux_v I__7261 (
            .O(N__38365),
            .I(N__38357));
    Odrv4 I__7260 (
            .O(N__38362),
            .I(\pid_front.error_p_regZ0Z_0 ));
    Odrv4 I__7259 (
            .O(N__38357),
            .I(\pid_front.error_p_regZ0Z_0 ));
    InMux I__7258 (
            .O(N__38352),
            .I(N__38349));
    LocalMux I__7257 (
            .O(N__38349),
            .I(N__38344));
    InMux I__7256 (
            .O(N__38348),
            .I(N__38341));
    InMux I__7255 (
            .O(N__38347),
            .I(N__38338));
    Span4Mux_h I__7254 (
            .O(N__38344),
            .I(N__38335));
    LocalMux I__7253 (
            .O(N__38341),
            .I(N__38332));
    LocalMux I__7252 (
            .O(N__38338),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    Odrv4 I__7251 (
            .O(N__38335),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    Odrv4 I__7250 (
            .O(N__38332),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    InMux I__7249 (
            .O(N__38325),
            .I(N__38321));
    InMux I__7248 (
            .O(N__38324),
            .I(N__38318));
    LocalMux I__7247 (
            .O(N__38321),
            .I(\pid_front.N_1427_i ));
    LocalMux I__7246 (
            .O(N__38318),
            .I(\pid_front.N_1427_i ));
    InMux I__7245 (
            .O(N__38313),
            .I(N__38310));
    LocalMux I__7244 (
            .O(N__38310),
            .I(N__38307));
    Odrv4 I__7243 (
            .O(N__38307),
            .I(\dron_frame_decoder_1.drone_H_disp_front_6 ));
    InMux I__7242 (
            .O(N__38304),
            .I(N__38298));
    InMux I__7241 (
            .O(N__38303),
            .I(N__38298));
    LocalMux I__7240 (
            .O(N__38298),
            .I(N__38295));
    Span4Mux_v I__7239 (
            .O(N__38295),
            .I(N__38290));
    InMux I__7238 (
            .O(N__38294),
            .I(N__38285));
    InMux I__7237 (
            .O(N__38293),
            .I(N__38285));
    Odrv4 I__7236 (
            .O(N__38290),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    LocalMux I__7235 (
            .O(N__38285),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    InMux I__7234 (
            .O(N__38280),
            .I(N__38274));
    InMux I__7233 (
            .O(N__38279),
            .I(N__38274));
    LocalMux I__7232 (
            .O(N__38274),
            .I(N__38271));
    Span4Mux_h I__7231 (
            .O(N__38271),
            .I(N__38268));
    Span4Mux_h I__7230 (
            .O(N__38268),
            .I(N__38265));
    Span4Mux_h I__7229 (
            .O(N__38265),
            .I(N__38262));
    Odrv4 I__7228 (
            .O(N__38262),
            .I(\pid_front.error_p_regZ0Z_4 ));
    InMux I__7227 (
            .O(N__38259),
            .I(N__38253));
    InMux I__7226 (
            .O(N__38258),
            .I(N__38253));
    LocalMux I__7225 (
            .O(N__38253),
            .I(\pid_front.error_d_reg_prevZ0Z_4 ));
    CascadeMux I__7224 (
            .O(N__38250),
            .I(N__38247));
    InMux I__7223 (
            .O(N__38247),
            .I(N__38243));
    InMux I__7222 (
            .O(N__38246),
            .I(N__38240));
    LocalMux I__7221 (
            .O(N__38243),
            .I(\pid_front.un1_pid_prereg_17 ));
    LocalMux I__7220 (
            .O(N__38240),
            .I(\pid_front.un1_pid_prereg_17 ));
    CascadeMux I__7219 (
            .O(N__38235),
            .I(\pid_front.un1_pid_prereg_17_cascade_ ));
    InMux I__7218 (
            .O(N__38232),
            .I(N__38225));
    InMux I__7217 (
            .O(N__38231),
            .I(N__38225));
    InMux I__7216 (
            .O(N__38230),
            .I(N__38222));
    LocalMux I__7215 (
            .O(N__38225),
            .I(\pid_front.un1_pid_prereg_3 ));
    LocalMux I__7214 (
            .O(N__38222),
            .I(\pid_front.un1_pid_prereg_3 ));
    InMux I__7213 (
            .O(N__38217),
            .I(N__38214));
    LocalMux I__7212 (
            .O(N__38214),
            .I(\pid_front.error_p_reg_esr_RNIPISGZ0Z_3 ));
    CascadeMux I__7211 (
            .O(N__38211),
            .I(\pid_front.error_p_reg_esr_RNI4KF7Z0Z_0_cascade_ ));
    InMux I__7210 (
            .O(N__38208),
            .I(N__38205));
    LocalMux I__7209 (
            .O(N__38205),
            .I(\pid_front.error_d_reg_esr_RNINGRVZ0Z_1 ));
    InMux I__7208 (
            .O(N__38202),
            .I(N__38196));
    InMux I__7207 (
            .O(N__38201),
            .I(N__38196));
    LocalMux I__7206 (
            .O(N__38196),
            .I(N__38193));
    Span12Mux_v I__7205 (
            .O(N__38193),
            .I(N__38190));
    Odrv12 I__7204 (
            .O(N__38190),
            .I(\pid_front.error_p_regZ0Z_1 ));
    InMux I__7203 (
            .O(N__38187),
            .I(N__38184));
    LocalMux I__7202 (
            .O(N__38184),
            .I(\ppm_encoder_1.un2_throttle_iv_1_13 ));
    InMux I__7201 (
            .O(N__38181),
            .I(N__38178));
    LocalMux I__7200 (
            .O(N__38178),
            .I(\ppm_encoder_1.N_299 ));
    CascadeMux I__7199 (
            .O(N__38175),
            .I(N__38172));
    InMux I__7198 (
            .O(N__38172),
            .I(N__38167));
    InMux I__7197 (
            .O(N__38171),
            .I(N__38162));
    InMux I__7196 (
            .O(N__38170),
            .I(N__38162));
    LocalMux I__7195 (
            .O(N__38167),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    LocalMux I__7194 (
            .O(N__38162),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    InMux I__7193 (
            .O(N__38157),
            .I(N__38154));
    LocalMux I__7192 (
            .O(N__38154),
            .I(N__38150));
    InMux I__7191 (
            .O(N__38153),
            .I(N__38147));
    Span4Mux_h I__7190 (
            .O(N__38150),
            .I(N__38144));
    LocalMux I__7189 (
            .O(N__38147),
            .I(N__38141));
    Span4Mux_v I__7188 (
            .O(N__38144),
            .I(N__38138));
    Span12Mux_h I__7187 (
            .O(N__38141),
            .I(N__38135));
    Odrv4 I__7186 (
            .O(N__38138),
            .I(front_order_13));
    Odrv12 I__7185 (
            .O(N__38135),
            .I(front_order_13));
    InMux I__7184 (
            .O(N__38130),
            .I(N__38127));
    LocalMux I__7183 (
            .O(N__38127),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__7182 (
            .O(N__38124),
            .I(N__38119));
    InMux I__7181 (
            .O(N__38123),
            .I(N__38114));
    InMux I__7180 (
            .O(N__38122),
            .I(N__38114));
    LocalMux I__7179 (
            .O(N__38119),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    LocalMux I__7178 (
            .O(N__38114),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__7177 (
            .O(N__38109),
            .I(N__38106));
    LocalMux I__7176 (
            .O(N__38106),
            .I(\dron_frame_decoder_1.drone_H_disp_front_7 ));
    InMux I__7175 (
            .O(N__38103),
            .I(N__38099));
    InMux I__7174 (
            .O(N__38102),
            .I(N__38096));
    LocalMux I__7173 (
            .O(N__38099),
            .I(N__38091));
    LocalMux I__7172 (
            .O(N__38096),
            .I(N__38091));
    Span4Mux_h I__7171 (
            .O(N__38091),
            .I(N__38088));
    Span4Mux_v I__7170 (
            .O(N__38088),
            .I(N__38085));
    Odrv4 I__7169 (
            .O(N__38085),
            .I(\pid_front.error_p_regZ0Z_2 ));
    InMux I__7168 (
            .O(N__38082),
            .I(N__38078));
    InMux I__7167 (
            .O(N__38081),
            .I(N__38075));
    LocalMux I__7166 (
            .O(N__38078),
            .I(\pid_front.error_d_reg_prevZ0Z_2 ));
    LocalMux I__7165 (
            .O(N__38075),
            .I(\pid_front.error_d_reg_prevZ0Z_2 ));
    CascadeMux I__7164 (
            .O(N__38070),
            .I(N__38067));
    InMux I__7163 (
            .O(N__38067),
            .I(N__38064));
    LocalMux I__7162 (
            .O(N__38064),
            .I(\pid_front.error_d_reg_esr_RNIOBP11Z0Z_5 ));
    InMux I__7161 (
            .O(N__38061),
            .I(N__38058));
    LocalMux I__7160 (
            .O(N__38058),
            .I(\pid_front.un1_pid_prereg_40_0 ));
    InMux I__7159 (
            .O(N__38055),
            .I(N__38052));
    LocalMux I__7158 (
            .O(N__38052),
            .I(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ));
    InMux I__7157 (
            .O(N__38049),
            .I(N__38041));
    InMux I__7156 (
            .O(N__38048),
            .I(N__38041));
    InMux I__7155 (
            .O(N__38047),
            .I(N__38036));
    InMux I__7154 (
            .O(N__38046),
            .I(N__38036));
    LocalMux I__7153 (
            .O(N__38041),
            .I(N__38033));
    LocalMux I__7152 (
            .O(N__38036),
            .I(N__38030));
    Span4Mux_v I__7151 (
            .O(N__38033),
            .I(N__38025));
    Span4Mux_h I__7150 (
            .O(N__38030),
            .I(N__38025));
    Span4Mux_h I__7149 (
            .O(N__38025),
            .I(N__38022));
    Span4Mux_v I__7148 (
            .O(N__38022),
            .I(N__38019));
    Odrv4 I__7147 (
            .O(N__38019),
            .I(\pid_front.error_p_regZ0Z_5 ));
    CascadeMux I__7146 (
            .O(N__38016),
            .I(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ));
    InMux I__7145 (
            .O(N__38013),
            .I(N__38010));
    LocalMux I__7144 (
            .O(N__38010),
            .I(N__38007));
    Span4Mux_h I__7143 (
            .O(N__38007),
            .I(N__38003));
    InMux I__7142 (
            .O(N__38006),
            .I(N__38000));
    Odrv4 I__7141 (
            .O(N__38003),
            .I(\pid_front.error_d_reg_esr_RNIVOSGZ0Z_5 ));
    LocalMux I__7140 (
            .O(N__38000),
            .I(\pid_front.error_d_reg_esr_RNIVOSGZ0Z_5 ));
    InMux I__7139 (
            .O(N__37995),
            .I(N__37990));
    InMux I__7138 (
            .O(N__37994),
            .I(N__37987));
    CascadeMux I__7137 (
            .O(N__37993),
            .I(N__37984));
    LocalMux I__7136 (
            .O(N__37990),
            .I(N__37979));
    LocalMux I__7135 (
            .O(N__37987),
            .I(N__37979));
    InMux I__7134 (
            .O(N__37984),
            .I(N__37976));
    Span4Mux_h I__7133 (
            .O(N__37979),
            .I(N__37973));
    LocalMux I__7132 (
            .O(N__37976),
            .I(front_order_8));
    Odrv4 I__7131 (
            .O(N__37973),
            .I(front_order_8));
    InMux I__7130 (
            .O(N__37968),
            .I(N__37965));
    LocalMux I__7129 (
            .O(N__37965),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__7128 (
            .O(N__37962),
            .I(bfn_13_17_0_));
    InMux I__7127 (
            .O(N__37959),
            .I(N__37956));
    LocalMux I__7126 (
            .O(N__37956),
            .I(N__37951));
    InMux I__7125 (
            .O(N__37955),
            .I(N__37948));
    CascadeMux I__7124 (
            .O(N__37954),
            .I(N__37945));
    Span4Mux_v I__7123 (
            .O(N__37951),
            .I(N__37940));
    LocalMux I__7122 (
            .O(N__37948),
            .I(N__37940));
    InMux I__7121 (
            .O(N__37945),
            .I(N__37937));
    Span4Mux_h I__7120 (
            .O(N__37940),
            .I(N__37934));
    LocalMux I__7119 (
            .O(N__37937),
            .I(front_order_9));
    Odrv4 I__7118 (
            .O(N__37934),
            .I(front_order_9));
    InMux I__7117 (
            .O(N__37929),
            .I(N__37926));
    LocalMux I__7116 (
            .O(N__37926),
            .I(N__37923));
    Odrv4 I__7115 (
            .O(N__37923),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__7114 (
            .O(N__37920),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__7113 (
            .O(N__37917),
            .I(N__37912));
    InMux I__7112 (
            .O(N__37916),
            .I(N__37909));
    CascadeMux I__7111 (
            .O(N__37915),
            .I(N__37906));
    LocalMux I__7110 (
            .O(N__37912),
            .I(N__37903));
    LocalMux I__7109 (
            .O(N__37909),
            .I(N__37900));
    InMux I__7108 (
            .O(N__37906),
            .I(N__37897));
    Span4Mux_v I__7107 (
            .O(N__37903),
            .I(N__37894));
    Span4Mux_h I__7106 (
            .O(N__37900),
            .I(N__37891));
    LocalMux I__7105 (
            .O(N__37897),
            .I(front_order_10));
    Odrv4 I__7104 (
            .O(N__37894),
            .I(front_order_10));
    Odrv4 I__7103 (
            .O(N__37891),
            .I(front_order_10));
    InMux I__7102 (
            .O(N__37884),
            .I(N__37881));
    LocalMux I__7101 (
            .O(N__37881),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__7100 (
            .O(N__37878),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__7099 (
            .O(N__37875),
            .I(N__37870));
    InMux I__7098 (
            .O(N__37874),
            .I(N__37867));
    CascadeMux I__7097 (
            .O(N__37873),
            .I(N__37864));
    LocalMux I__7096 (
            .O(N__37870),
            .I(N__37861));
    LocalMux I__7095 (
            .O(N__37867),
            .I(N__37858));
    InMux I__7094 (
            .O(N__37864),
            .I(N__37855));
    Span4Mux_h I__7093 (
            .O(N__37861),
            .I(N__37852));
    Span4Mux_h I__7092 (
            .O(N__37858),
            .I(N__37849));
    LocalMux I__7091 (
            .O(N__37855),
            .I(front_order_11));
    Odrv4 I__7090 (
            .O(N__37852),
            .I(front_order_11));
    Odrv4 I__7089 (
            .O(N__37849),
            .I(front_order_11));
    InMux I__7088 (
            .O(N__37842),
            .I(N__37839));
    LocalMux I__7087 (
            .O(N__37839),
            .I(N__37836));
    Odrv4 I__7086 (
            .O(N__37836),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__7085 (
            .O(N__37833),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__7084 (
            .O(N__37830),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__7083 (
            .O(N__37827),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__7082 (
            .O(N__37824),
            .I(\ppm_encoder_1.un1_elevator_cry_13 ));
    InMux I__7081 (
            .O(N__37821),
            .I(N__37817));
    InMux I__7080 (
            .O(N__37820),
            .I(N__37814));
    LocalMux I__7079 (
            .O(N__37817),
            .I(N__37808));
    LocalMux I__7078 (
            .O(N__37814),
            .I(N__37808));
    InMux I__7077 (
            .O(N__37813),
            .I(N__37805));
    Span4Mux_h I__7076 (
            .O(N__37808),
            .I(N__37802));
    LocalMux I__7075 (
            .O(N__37805),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    Odrv4 I__7074 (
            .O(N__37802),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    CascadeMux I__7073 (
            .O(N__37797),
            .I(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ));
    InMux I__7072 (
            .O(N__37794),
            .I(\ppm_encoder_1.un1_elevator_cry_0 ));
    InMux I__7071 (
            .O(N__37791),
            .I(N__37787));
    InMux I__7070 (
            .O(N__37790),
            .I(N__37784));
    LocalMux I__7069 (
            .O(N__37787),
            .I(N__37779));
    LocalMux I__7068 (
            .O(N__37784),
            .I(N__37779));
    Span4Mux_h I__7067 (
            .O(N__37779),
            .I(N__37776));
    Odrv4 I__7066 (
            .O(N__37776),
            .I(front_order_2));
    InMux I__7065 (
            .O(N__37773),
            .I(N__37770));
    LocalMux I__7064 (
            .O(N__37770),
            .I(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ));
    InMux I__7063 (
            .O(N__37767),
            .I(\ppm_encoder_1.un1_elevator_cry_1 ));
    InMux I__7062 (
            .O(N__37764),
            .I(\ppm_encoder_1.un1_elevator_cry_2 ));
    InMux I__7061 (
            .O(N__37761),
            .I(N__37757));
    InMux I__7060 (
            .O(N__37760),
            .I(N__37754));
    LocalMux I__7059 (
            .O(N__37757),
            .I(N__37751));
    LocalMux I__7058 (
            .O(N__37754),
            .I(N__37748));
    Span4Mux_v I__7057 (
            .O(N__37751),
            .I(N__37743));
    Span4Mux_h I__7056 (
            .O(N__37748),
            .I(N__37743));
    Span4Mux_v I__7055 (
            .O(N__37743),
            .I(N__37740));
    Odrv4 I__7054 (
            .O(N__37740),
            .I(front_order_4));
    InMux I__7053 (
            .O(N__37737),
            .I(N__37734));
    LocalMux I__7052 (
            .O(N__37734),
            .I(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ));
    InMux I__7051 (
            .O(N__37731),
            .I(\ppm_encoder_1.un1_elevator_cry_3 ));
    InMux I__7050 (
            .O(N__37728),
            .I(N__37724));
    InMux I__7049 (
            .O(N__37727),
            .I(N__37721));
    LocalMux I__7048 (
            .O(N__37724),
            .I(N__37718));
    LocalMux I__7047 (
            .O(N__37721),
            .I(N__37715));
    Span4Mux_h I__7046 (
            .O(N__37718),
            .I(N__37712));
    Span4Mux_h I__7045 (
            .O(N__37715),
            .I(N__37709));
    Span4Mux_v I__7044 (
            .O(N__37712),
            .I(N__37706));
    Span4Mux_v I__7043 (
            .O(N__37709),
            .I(N__37703));
    Odrv4 I__7042 (
            .O(N__37706),
            .I(front_order_5));
    Odrv4 I__7041 (
            .O(N__37703),
            .I(front_order_5));
    InMux I__7040 (
            .O(N__37698),
            .I(N__37695));
    LocalMux I__7039 (
            .O(N__37695),
            .I(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ));
    InMux I__7038 (
            .O(N__37692),
            .I(\ppm_encoder_1.un1_elevator_cry_4 ));
    InMux I__7037 (
            .O(N__37689),
            .I(N__37685));
    CascadeMux I__7036 (
            .O(N__37688),
            .I(N__37682));
    LocalMux I__7035 (
            .O(N__37685),
            .I(N__37678));
    InMux I__7034 (
            .O(N__37682),
            .I(N__37675));
    CascadeMux I__7033 (
            .O(N__37681),
            .I(N__37672));
    Span4Mux_v I__7032 (
            .O(N__37678),
            .I(N__37667));
    LocalMux I__7031 (
            .O(N__37675),
            .I(N__37667));
    InMux I__7030 (
            .O(N__37672),
            .I(N__37664));
    Span4Mux_h I__7029 (
            .O(N__37667),
            .I(N__37661));
    LocalMux I__7028 (
            .O(N__37664),
            .I(front_order_6));
    Odrv4 I__7027 (
            .O(N__37661),
            .I(front_order_6));
    InMux I__7026 (
            .O(N__37656),
            .I(N__37653));
    LocalMux I__7025 (
            .O(N__37653),
            .I(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ));
    InMux I__7024 (
            .O(N__37650),
            .I(\ppm_encoder_1.un1_elevator_cry_5 ));
    InMux I__7023 (
            .O(N__37647),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    CascadeMux I__7022 (
            .O(N__37644),
            .I(\ppm_encoder_1.N_134_0_cascade_ ));
    IoInMux I__7021 (
            .O(N__37641),
            .I(N__37638));
    LocalMux I__7020 (
            .O(N__37638),
            .I(N__37635));
    Span12Mux_s11_v I__7019 (
            .O(N__37635),
            .I(N__37631));
    InMux I__7018 (
            .O(N__37634),
            .I(N__37628));
    Odrv12 I__7017 (
            .O(N__37631),
            .I(ppm_output_c));
    LocalMux I__7016 (
            .O(N__37628),
            .I(ppm_output_c));
    InMux I__7015 (
            .O(N__37623),
            .I(N__37620));
    LocalMux I__7014 (
            .O(N__37620),
            .I(N__37617));
    Odrv12 I__7013 (
            .O(N__37617),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    InMux I__7012 (
            .O(N__37614),
            .I(N__37610));
    InMux I__7011 (
            .O(N__37613),
            .I(N__37607));
    LocalMux I__7010 (
            .O(N__37610),
            .I(N__37602));
    LocalMux I__7009 (
            .O(N__37607),
            .I(N__37602));
    Span12Mux_h I__7008 (
            .O(N__37602),
            .I(N__37599));
    Odrv12 I__7007 (
            .O(N__37599),
            .I(throttle_order_2));
    InMux I__7006 (
            .O(N__37596),
            .I(N__37592));
    InMux I__7005 (
            .O(N__37595),
            .I(N__37589));
    LocalMux I__7004 (
            .O(N__37592),
            .I(N__37586));
    LocalMux I__7003 (
            .O(N__37589),
            .I(N__37583));
    Odrv12 I__7002 (
            .O(N__37586),
            .I(scaler_4_data_6));
    Odrv4 I__7001 (
            .O(N__37583),
            .I(scaler_4_data_6));
    InMux I__7000 (
            .O(N__37578),
            .I(N__37575));
    LocalMux I__6999 (
            .O(N__37575),
            .I(N__37572));
    Span4Mux_h I__6998 (
            .O(N__37572),
            .I(N__37569));
    Span4Mux_h I__6997 (
            .O(N__37569),
            .I(N__37566));
    Odrv4 I__6996 (
            .O(N__37566),
            .I(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ));
    CascadeMux I__6995 (
            .O(N__37563),
            .I(N__37560));
    InMux I__6994 (
            .O(N__37560),
            .I(N__37554));
    InMux I__6993 (
            .O(N__37559),
            .I(N__37554));
    LocalMux I__6992 (
            .O(N__37554),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__6991 (
            .O(N__37551),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    CascadeMux I__6990 (
            .O(N__37548),
            .I(N__37545));
    InMux I__6989 (
            .O(N__37545),
            .I(N__37539));
    InMux I__6988 (
            .O(N__37544),
            .I(N__37539));
    LocalMux I__6987 (
            .O(N__37539),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__6986 (
            .O(N__37536),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    CascadeMux I__6985 (
            .O(N__37533),
            .I(N__37530));
    InMux I__6984 (
            .O(N__37530),
            .I(N__37524));
    InMux I__6983 (
            .O(N__37529),
            .I(N__37524));
    LocalMux I__6982 (
            .O(N__37524),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__6981 (
            .O(N__37521),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    CascadeMux I__6980 (
            .O(N__37518),
            .I(N__37515));
    InMux I__6979 (
            .O(N__37515),
            .I(N__37509));
    InMux I__6978 (
            .O(N__37514),
            .I(N__37509));
    LocalMux I__6977 (
            .O(N__37509),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__6976 (
            .O(N__37506),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__6975 (
            .O(N__37503),
            .I(N__37499));
    InMux I__6974 (
            .O(N__37502),
            .I(N__37496));
    LocalMux I__6973 (
            .O(N__37499),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    LocalMux I__6972 (
            .O(N__37496),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    CascadeMux I__6971 (
            .O(N__37491),
            .I(N__37488));
    InMux I__6970 (
            .O(N__37488),
            .I(N__37485));
    LocalMux I__6969 (
            .O(N__37485),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__6968 (
            .O(N__37482),
            .I(bfn_13_13_0_));
    InMux I__6967 (
            .O(N__37479),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    InMux I__6966 (
            .O(N__37476),
            .I(N__37473));
    LocalMux I__6965 (
            .O(N__37473),
            .I(N__37470));
    Odrv4 I__6964 (
            .O(N__37470),
            .I(scaler_4_data_14));
    CEMux I__6963 (
            .O(N__37467),
            .I(N__37463));
    CEMux I__6962 (
            .O(N__37466),
            .I(N__37460));
    LocalMux I__6961 (
            .O(N__37463),
            .I(N__37457));
    LocalMux I__6960 (
            .O(N__37460),
            .I(N__37454));
    Span4Mux_v I__6959 (
            .O(N__37457),
            .I(N__37448));
    Span4Mux_v I__6958 (
            .O(N__37454),
            .I(N__37448));
    CEMux I__6957 (
            .O(N__37453),
            .I(N__37445));
    Sp12to4 I__6956 (
            .O(N__37448),
            .I(N__37440));
    LocalMux I__6955 (
            .O(N__37445),
            .I(N__37440));
    Odrv12 I__6954 (
            .O(N__37440),
            .I(\scaler_4.debug_CH3_20A_c_0 ));
    InMux I__6953 (
            .O(N__37437),
            .I(N__37434));
    LocalMux I__6952 (
            .O(N__37434),
            .I(N__37431));
    Odrv12 I__6951 (
            .O(N__37431),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__6950 (
            .O(N__37428),
            .I(N__37424));
    InMux I__6949 (
            .O(N__37427),
            .I(N__37421));
    LocalMux I__6948 (
            .O(N__37424),
            .I(N__37418));
    LocalMux I__6947 (
            .O(N__37421),
            .I(N__37415));
    Odrv4 I__6946 (
            .O(N__37418),
            .I(scaler_4_data_7));
    Odrv4 I__6945 (
            .O(N__37415),
            .I(scaler_4_data_7));
    InMux I__6944 (
            .O(N__37410),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__6943 (
            .O(N__37407),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__6942 (
            .O(N__37404),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__6941 (
            .O(N__37401),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__6940 (
            .O(N__37398),
            .I(bfn_13_11_0_));
    InMux I__6939 (
            .O(N__37395),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    CascadeMux I__6938 (
            .O(N__37392),
            .I(N__37389));
    InMux I__6937 (
            .O(N__37389),
            .I(N__37383));
    InMux I__6936 (
            .O(N__37388),
            .I(N__37383));
    LocalMux I__6935 (
            .O(N__37383),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__6934 (
            .O(N__37380),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    CascadeMux I__6933 (
            .O(N__37377),
            .I(N__37374));
    InMux I__6932 (
            .O(N__37374),
            .I(N__37368));
    InMux I__6931 (
            .O(N__37373),
            .I(N__37368));
    LocalMux I__6930 (
            .O(N__37368),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    InMux I__6929 (
            .O(N__37365),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    InMux I__6928 (
            .O(N__37362),
            .I(N__37356));
    InMux I__6927 (
            .O(N__37361),
            .I(N__37356));
    LocalMux I__6926 (
            .O(N__37356),
            .I(N__37353));
    Span12Mux_h I__6925 (
            .O(N__37353),
            .I(N__37350));
    Odrv12 I__6924 (
            .O(N__37350),
            .I(\pid_front.error_p_regZ0Z_20 ));
    InMux I__6923 (
            .O(N__37347),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__6922 (
            .O(N__37344),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__6921 (
            .O(N__37341),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    CEMux I__6920 (
            .O(N__37338),
            .I(N__37335));
    LocalMux I__6919 (
            .O(N__37335),
            .I(N__37332));
    Span4Mux_h I__6918 (
            .O(N__37332),
            .I(N__37329));
    Span4Mux_h I__6917 (
            .O(N__37329),
            .I(N__37326));
    Sp12to4 I__6916 (
            .O(N__37326),
            .I(N__37323));
    Odrv12 I__6915 (
            .O(N__37323),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__6914 (
            .O(N__37320),
            .I(N__37317));
    LocalMux I__6913 (
            .O(N__37317),
            .I(N__37314));
    Odrv4 I__6912 (
            .O(N__37314),
            .I(\pid_front.un1_pid_prereg_axb_21 ));
    CascadeMux I__6911 (
            .O(N__37311),
            .I(N__37308));
    InMux I__6910 (
            .O(N__37308),
            .I(N__37302));
    InMux I__6909 (
            .O(N__37307),
            .I(N__37302));
    LocalMux I__6908 (
            .O(N__37302),
            .I(front_command_7));
    InMux I__6907 (
            .O(N__37299),
            .I(N__37296));
    LocalMux I__6906 (
            .O(N__37296),
            .I(N__37293));
    Odrv4 I__6905 (
            .O(N__37293),
            .I(\pid_front.error_p_reg_esr_RNIHGOC2Z0Z_16 ));
    CascadeMux I__6904 (
            .O(N__37290),
            .I(N__37287));
    InMux I__6903 (
            .O(N__37287),
            .I(N__37284));
    LocalMux I__6902 (
            .O(N__37284),
            .I(N__37281));
    Odrv4 I__6901 (
            .O(N__37281),
            .I(\pid_front.error_p_reg_esr_RNI87HP4Z0Z_16 ));
    CascadeMux I__6900 (
            .O(N__37278),
            .I(N__37275));
    InMux I__6899 (
            .O(N__37275),
            .I(N__37272));
    LocalMux I__6898 (
            .O(N__37272),
            .I(\pid_front.pid_preregZ0Z_18 ));
    InMux I__6897 (
            .O(N__37269),
            .I(\pid_front.un1_pid_prereg_cry_15 ));
    InMux I__6896 (
            .O(N__37266),
            .I(N__37263));
    LocalMux I__6895 (
            .O(N__37263),
            .I(N__37260));
    Odrv4 I__6894 (
            .O(N__37260),
            .I(\pid_front.error_p_reg_esr_RNINMOC2Z0Z_17 ));
    CascadeMux I__6893 (
            .O(N__37257),
            .I(N__37254));
    InMux I__6892 (
            .O(N__37254),
            .I(N__37251));
    LocalMux I__6891 (
            .O(N__37251),
            .I(N__37248));
    Odrv4 I__6890 (
            .O(N__37248),
            .I(\pid_front.error_p_reg_esr_RNIKJHP4Z0Z_17 ));
    InMux I__6889 (
            .O(N__37245),
            .I(N__37242));
    LocalMux I__6888 (
            .O(N__37242),
            .I(\pid_front.pid_preregZ0Z_19 ));
    InMux I__6887 (
            .O(N__37239),
            .I(\pid_front.un1_pid_prereg_cry_16 ));
    InMux I__6886 (
            .O(N__37236),
            .I(N__37233));
    LocalMux I__6885 (
            .O(N__37233),
            .I(N__37230));
    Odrv12 I__6884 (
            .O(N__37230),
            .I(\pid_front.error_p_reg_esr_RNITSOC2Z0Z_18 ));
    CascadeMux I__6883 (
            .O(N__37227),
            .I(N__37224));
    InMux I__6882 (
            .O(N__37224),
            .I(N__37221));
    LocalMux I__6881 (
            .O(N__37221),
            .I(N__37218));
    Span4Mux_h I__6880 (
            .O(N__37218),
            .I(N__37215));
    Odrv4 I__6879 (
            .O(N__37215),
            .I(\pid_front.error_p_reg_esr_RNI57KP4Z0Z_18 ));
    InMux I__6878 (
            .O(N__37212),
            .I(N__37209));
    LocalMux I__6877 (
            .O(N__37209),
            .I(\pid_front.pid_preregZ0Z_20 ));
    InMux I__6876 (
            .O(N__37206),
            .I(\pid_front.un1_pid_prereg_cry_17 ));
    InMux I__6875 (
            .O(N__37203),
            .I(N__37200));
    LocalMux I__6874 (
            .O(N__37200),
            .I(N__37197));
    Odrv12 I__6873 (
            .O(N__37197),
            .I(\pid_front.error_p_reg_esr_RNI8ARC2Z0Z_19 ));
    CascadeMux I__6872 (
            .O(N__37194),
            .I(N__37191));
    InMux I__6871 (
            .O(N__37191),
            .I(N__37188));
    LocalMux I__6870 (
            .O(N__37188),
            .I(N__37185));
    Span4Mux_v I__6869 (
            .O(N__37185),
            .I(N__37182));
    Odrv4 I__6868 (
            .O(N__37182),
            .I(\pid_front.error_p_reg_esr_RNIOUOP4Z0Z_19 ));
    InMux I__6867 (
            .O(N__37179),
            .I(N__37176));
    LocalMux I__6866 (
            .O(N__37176),
            .I(\pid_front.pid_preregZ0Z_21 ));
    InMux I__6865 (
            .O(N__37173),
            .I(\pid_front.un1_pid_prereg_cry_18 ));
    InMux I__6864 (
            .O(N__37170),
            .I(N__37167));
    LocalMux I__6863 (
            .O(N__37167),
            .I(N__37164));
    Span4Mux_h I__6862 (
            .O(N__37164),
            .I(N__37161));
    Odrv4 I__6861 (
            .O(N__37161),
            .I(\pid_front.error_p_reg_esr_RNI09RP4Z0Z_20 ));
    InMux I__6860 (
            .O(N__37158),
            .I(N__37155));
    LocalMux I__6859 (
            .O(N__37155),
            .I(\pid_front.pid_preregZ0Z_22 ));
    InMux I__6858 (
            .O(N__37152),
            .I(\pid_front.un1_pid_prereg_cry_19 ));
    InMux I__6857 (
            .O(N__37149),
            .I(\pid_front.un1_pid_prereg_cry_20 ));
    CascadeMux I__6856 (
            .O(N__37146),
            .I(N__37143));
    InMux I__6855 (
            .O(N__37143),
            .I(N__37136));
    InMux I__6854 (
            .O(N__37142),
            .I(N__37131));
    InMux I__6853 (
            .O(N__37141),
            .I(N__37131));
    InMux I__6852 (
            .O(N__37140),
            .I(N__37128));
    CascadeMux I__6851 (
            .O(N__37139),
            .I(N__37125));
    LocalMux I__6850 (
            .O(N__37136),
            .I(N__37121));
    LocalMux I__6849 (
            .O(N__37131),
            .I(N__37118));
    LocalMux I__6848 (
            .O(N__37128),
            .I(N__37115));
    InMux I__6847 (
            .O(N__37125),
            .I(N__37110));
    InMux I__6846 (
            .O(N__37124),
            .I(N__37110));
    Span4Mux_v I__6845 (
            .O(N__37121),
            .I(N__37105));
    Span4Mux_v I__6844 (
            .O(N__37118),
            .I(N__37105));
    Span4Mux_h I__6843 (
            .O(N__37115),
            .I(N__37102));
    LocalMux I__6842 (
            .O(N__37110),
            .I(\pid_front.pid_preregZ0Z_23 ));
    Odrv4 I__6841 (
            .O(N__37105),
            .I(\pid_front.pid_preregZ0Z_23 ));
    Odrv4 I__6840 (
            .O(N__37102),
            .I(\pid_front.pid_preregZ0Z_23 ));
    InMux I__6839 (
            .O(N__37095),
            .I(\pid_front.un1_pid_prereg_cry_7 ));
    InMux I__6838 (
            .O(N__37092),
            .I(N__37089));
    LocalMux I__6837 (
            .O(N__37089),
            .I(N__37086));
    Odrv4 I__6836 (
            .O(N__37086),
            .I(\pid_front.error_d_reg_esr_RNI9NAB3Z0Z_10 ));
    CascadeMux I__6835 (
            .O(N__37083),
            .I(N__37079));
    CascadeMux I__6834 (
            .O(N__37082),
            .I(N__37076));
    InMux I__6833 (
            .O(N__37079),
            .I(N__37073));
    InMux I__6832 (
            .O(N__37076),
            .I(N__37070));
    LocalMux I__6831 (
            .O(N__37073),
            .I(N__37067));
    LocalMux I__6830 (
            .O(N__37070),
            .I(\pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10 ));
    Odrv4 I__6829 (
            .O(N__37067),
            .I(\pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10 ));
    InMux I__6828 (
            .O(N__37062),
            .I(N__37059));
    LocalMux I__6827 (
            .O(N__37059),
            .I(N__37056));
    Span4Mux_h I__6826 (
            .O(N__37056),
            .I(N__37050));
    InMux I__6825 (
            .O(N__37055),
            .I(N__37043));
    InMux I__6824 (
            .O(N__37054),
            .I(N__37043));
    InMux I__6823 (
            .O(N__37053),
            .I(N__37043));
    Odrv4 I__6822 (
            .O(N__37050),
            .I(\pid_front.pid_preregZ0Z_11 ));
    LocalMux I__6821 (
            .O(N__37043),
            .I(\pid_front.pid_preregZ0Z_11 ));
    InMux I__6820 (
            .O(N__37038),
            .I(\pid_front.un1_pid_prereg_cry_8 ));
    InMux I__6819 (
            .O(N__37035),
            .I(N__37032));
    LocalMux I__6818 (
            .O(N__37032),
            .I(N__37029));
    Span4Mux_h I__6817 (
            .O(N__37029),
            .I(N__37026));
    Odrv4 I__6816 (
            .O(N__37026),
            .I(\pid_front.error_p_reg_esr_RNIESET1Z0Z_10 ));
    CascadeMux I__6815 (
            .O(N__37023),
            .I(N__37020));
    InMux I__6814 (
            .O(N__37020),
            .I(N__37017));
    LocalMux I__6813 (
            .O(N__37017),
            .I(N__37014));
    Span4Mux_h I__6812 (
            .O(N__37014),
            .I(N__37011));
    Odrv4 I__6811 (
            .O(N__37011),
            .I(\pid_front.error_p_reg_esr_RNI1E6A4Z0Z_12 ));
    InMux I__6810 (
            .O(N__37008),
            .I(N__37005));
    LocalMux I__6809 (
            .O(N__37005),
            .I(N__36999));
    InMux I__6808 (
            .O(N__37004),
            .I(N__36992));
    InMux I__6807 (
            .O(N__37003),
            .I(N__36992));
    InMux I__6806 (
            .O(N__37002),
            .I(N__36992));
    Odrv4 I__6805 (
            .O(N__36999),
            .I(\pid_front.pid_preregZ0Z_12 ));
    LocalMux I__6804 (
            .O(N__36992),
            .I(\pid_front.pid_preregZ0Z_12 ));
    InMux I__6803 (
            .O(N__36987),
            .I(\pid_front.un1_pid_prereg_cry_9 ));
    InMux I__6802 (
            .O(N__36984),
            .I(N__36980));
    InMux I__6801 (
            .O(N__36983),
            .I(N__36977));
    LocalMux I__6800 (
            .O(N__36980),
            .I(N__36974));
    LocalMux I__6799 (
            .O(N__36977),
            .I(\pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12 ));
    Odrv4 I__6798 (
            .O(N__36974),
            .I(\pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12 ));
    CascadeMux I__6797 (
            .O(N__36969),
            .I(N__36966));
    InMux I__6796 (
            .O(N__36966),
            .I(N__36963));
    LocalMux I__6795 (
            .O(N__36963),
            .I(N__36960));
    Odrv12 I__6794 (
            .O(N__36960),
            .I(\pid_front.error_d_reg_esr_RNIBO6A4Z0Z_12 ));
    InMux I__6793 (
            .O(N__36957),
            .I(N__36953));
    InMux I__6792 (
            .O(N__36956),
            .I(N__36950));
    LocalMux I__6791 (
            .O(N__36953),
            .I(N__36943));
    LocalMux I__6790 (
            .O(N__36950),
            .I(N__36943));
    InMux I__6789 (
            .O(N__36949),
            .I(N__36937));
    InMux I__6788 (
            .O(N__36948),
            .I(N__36937));
    Span4Mux_h I__6787 (
            .O(N__36943),
            .I(N__36934));
    InMux I__6786 (
            .O(N__36942),
            .I(N__36931));
    LocalMux I__6785 (
            .O(N__36937),
            .I(\pid_front.pid_preregZ0Z_13 ));
    Odrv4 I__6784 (
            .O(N__36934),
            .I(\pid_front.pid_preregZ0Z_13 ));
    LocalMux I__6783 (
            .O(N__36931),
            .I(\pid_front.pid_preregZ0Z_13 ));
    InMux I__6782 (
            .O(N__36924),
            .I(\pid_front.un1_pid_prereg_cry_10 ));
    InMux I__6781 (
            .O(N__36921),
            .I(N__36918));
    LocalMux I__6780 (
            .O(N__36918),
            .I(N__36915));
    Odrv12 I__6779 (
            .O(N__36915),
            .I(\pid_front.error_p_reg_esr_RNIO6FT1Z0Z_12 ));
    CascadeMux I__6778 (
            .O(N__36912),
            .I(N__36909));
    InMux I__6777 (
            .O(N__36909),
            .I(N__36906));
    LocalMux I__6776 (
            .O(N__36906),
            .I(N__36903));
    Odrv12 I__6775 (
            .O(N__36903),
            .I(\pid_front.error_p_reg_esr_RNIN47A4Z0Z_12 ));
    InMux I__6774 (
            .O(N__36900),
            .I(N__36897));
    LocalMux I__6773 (
            .O(N__36897),
            .I(\pid_front.pid_preregZ0Z_14 ));
    InMux I__6772 (
            .O(N__36894),
            .I(\pid_front.un1_pid_prereg_cry_11 ));
    InMux I__6771 (
            .O(N__36891),
            .I(N__36888));
    LocalMux I__6770 (
            .O(N__36888),
            .I(N__36885));
    Span4Mux_h I__6769 (
            .O(N__36885),
            .I(N__36882));
    Odrv4 I__6768 (
            .O(N__36882),
            .I(\pid_front.error_p_reg_esr_RNI42GP4Z0Z_13 ));
    CascadeMux I__6767 (
            .O(N__36879),
            .I(N__36876));
    InMux I__6766 (
            .O(N__36876),
            .I(N__36873));
    LocalMux I__6765 (
            .O(N__36873),
            .I(N__36870));
    Span4Mux_h I__6764 (
            .O(N__36870),
            .I(N__36867));
    Odrv4 I__6763 (
            .O(N__36867),
            .I(\pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13 ));
    InMux I__6762 (
            .O(N__36864),
            .I(N__36861));
    LocalMux I__6761 (
            .O(N__36861),
            .I(\pid_front.pid_preregZ0Z_15 ));
    InMux I__6760 (
            .O(N__36858),
            .I(\pid_front.un1_pid_prereg_cry_12 ));
    InMux I__6759 (
            .O(N__36855),
            .I(N__36852));
    LocalMux I__6758 (
            .O(N__36852),
            .I(N__36849));
    Odrv12 I__6757 (
            .O(N__36849),
            .I(\pid_front.error_p_reg_esr_RNI54OC2Z0Z_14 ));
    CascadeMux I__6756 (
            .O(N__36846),
            .I(N__36843));
    InMux I__6755 (
            .O(N__36843),
            .I(N__36840));
    LocalMux I__6754 (
            .O(N__36840),
            .I(N__36837));
    Span4Mux_h I__6753 (
            .O(N__36837),
            .I(N__36834));
    Odrv4 I__6752 (
            .O(N__36834),
            .I(\pid_front.error_p_reg_esr_RNIGEGP4Z0Z_14 ));
    InMux I__6751 (
            .O(N__36831),
            .I(N__36828));
    LocalMux I__6750 (
            .O(N__36828),
            .I(\pid_front.pid_preregZ0Z_16 ));
    InMux I__6749 (
            .O(N__36825),
            .I(bfn_12_23_0_));
    InMux I__6748 (
            .O(N__36822),
            .I(N__36819));
    LocalMux I__6747 (
            .O(N__36819),
            .I(N__36816));
    Odrv12 I__6746 (
            .O(N__36816),
            .I(\pid_front.error_p_reg_esr_RNIBAOC2Z0Z_15 ));
    CascadeMux I__6745 (
            .O(N__36813),
            .I(N__36810));
    InMux I__6744 (
            .O(N__36810),
            .I(N__36807));
    LocalMux I__6743 (
            .O(N__36807),
            .I(N__36804));
    Odrv12 I__6742 (
            .O(N__36804),
            .I(\pid_front.error_p_reg_esr_RNISQGP4Z0Z_15 ));
    InMux I__6741 (
            .O(N__36801),
            .I(N__36798));
    LocalMux I__6740 (
            .O(N__36798),
            .I(\pid_front.pid_preregZ0Z_17 ));
    InMux I__6739 (
            .O(N__36795),
            .I(\pid_front.un1_pid_prereg_cry_14 ));
    CascadeMux I__6738 (
            .O(N__36792),
            .I(N__36789));
    InMux I__6737 (
            .O(N__36789),
            .I(N__36786));
    LocalMux I__6736 (
            .O(N__36786),
            .I(N__36783));
    Odrv4 I__6735 (
            .O(N__36783),
            .I(\pid_front.error_p_reg_esr_RNIH7Q01Z0Z_1 ));
    CascadeMux I__6734 (
            .O(N__36780),
            .I(N__36777));
    InMux I__6733 (
            .O(N__36777),
            .I(N__36773));
    CascadeMux I__6732 (
            .O(N__36776),
            .I(N__36770));
    LocalMux I__6731 (
            .O(N__36773),
            .I(N__36767));
    InMux I__6730 (
            .O(N__36770),
            .I(N__36764));
    Span4Mux_h I__6729 (
            .O(N__36767),
            .I(N__36761));
    LocalMux I__6728 (
            .O(N__36764),
            .I(\pid_front.pid_preregZ0Z_3 ));
    Odrv4 I__6727 (
            .O(N__36761),
            .I(\pid_front.pid_preregZ0Z_3 ));
    InMux I__6726 (
            .O(N__36756),
            .I(\pid_front.un1_pid_prereg_cry_0_0 ));
    InMux I__6725 (
            .O(N__36753),
            .I(N__36750));
    LocalMux I__6724 (
            .O(N__36750),
            .I(N__36747));
    Odrv4 I__6723 (
            .O(N__36747),
            .I(\pid_front.error_p_reg_esr_RNIJCSGZ0Z_2 ));
    CascadeMux I__6722 (
            .O(N__36744),
            .I(N__36741));
    InMux I__6721 (
            .O(N__36741),
            .I(N__36738));
    LocalMux I__6720 (
            .O(N__36738),
            .I(N__36735));
    Odrv4 I__6719 (
            .O(N__36735),
            .I(\pid_front.error_p_reg_esr_RNICVO11Z0Z_2 ));
    InMux I__6718 (
            .O(N__36732),
            .I(N__36728));
    CascadeMux I__6717 (
            .O(N__36731),
            .I(N__36720));
    LocalMux I__6716 (
            .O(N__36728),
            .I(N__36717));
    InMux I__6715 (
            .O(N__36727),
            .I(N__36712));
    InMux I__6714 (
            .O(N__36726),
            .I(N__36712));
    InMux I__6713 (
            .O(N__36725),
            .I(N__36705));
    InMux I__6712 (
            .O(N__36724),
            .I(N__36705));
    InMux I__6711 (
            .O(N__36723),
            .I(N__36705));
    InMux I__6710 (
            .O(N__36720),
            .I(N__36702));
    Span4Mux_v I__6709 (
            .O(N__36717),
            .I(N__36699));
    LocalMux I__6708 (
            .O(N__36712),
            .I(\pid_front.pid_preregZ0Z_4 ));
    LocalMux I__6707 (
            .O(N__36705),
            .I(\pid_front.pid_preregZ0Z_4 ));
    LocalMux I__6706 (
            .O(N__36702),
            .I(\pid_front.pid_preregZ0Z_4 ));
    Odrv4 I__6705 (
            .O(N__36699),
            .I(\pid_front.pid_preregZ0Z_4 ));
    InMux I__6704 (
            .O(N__36690),
            .I(\pid_front.un1_pid_prereg_cry_1_0 ));
    CascadeMux I__6703 (
            .O(N__36687),
            .I(N__36682));
    CascadeMux I__6702 (
            .O(N__36686),
            .I(N__36679));
    CascadeMux I__6701 (
            .O(N__36685),
            .I(N__36675));
    InMux I__6700 (
            .O(N__36682),
            .I(N__36670));
    InMux I__6699 (
            .O(N__36679),
            .I(N__36670));
    InMux I__6698 (
            .O(N__36678),
            .I(N__36667));
    InMux I__6697 (
            .O(N__36675),
            .I(N__36664));
    LocalMux I__6696 (
            .O(N__36670),
            .I(N__36661));
    LocalMux I__6695 (
            .O(N__36667),
            .I(N__36658));
    LocalMux I__6694 (
            .O(N__36664),
            .I(N__36655));
    Span4Mux_v I__6693 (
            .O(N__36661),
            .I(N__36650));
    Span4Mux_h I__6692 (
            .O(N__36658),
            .I(N__36650));
    Odrv4 I__6691 (
            .O(N__36655),
            .I(\pid_front.pid_preregZ0Z_5 ));
    Odrv4 I__6690 (
            .O(N__36650),
            .I(\pid_front.pid_preregZ0Z_5 ));
    InMux I__6689 (
            .O(N__36645),
            .I(\pid_front.un1_pid_prereg_cry_2 ));
    CascadeMux I__6688 (
            .O(N__36642),
            .I(N__36639));
    InMux I__6687 (
            .O(N__36639),
            .I(N__36636));
    LocalMux I__6686 (
            .O(N__36636),
            .I(\pid_front.error_p_reg_esr_RNIH8R01Z0Z_5 ));
    InMux I__6685 (
            .O(N__36633),
            .I(N__36630));
    LocalMux I__6684 (
            .O(N__36630),
            .I(N__36627));
    Span4Mux_h I__6683 (
            .O(N__36627),
            .I(N__36622));
    InMux I__6682 (
            .O(N__36626),
            .I(N__36619));
    InMux I__6681 (
            .O(N__36625),
            .I(N__36616));
    Odrv4 I__6680 (
            .O(N__36622),
            .I(\pid_front.pid_preregZ0Z_6 ));
    LocalMux I__6679 (
            .O(N__36619),
            .I(\pid_front.pid_preregZ0Z_6 ));
    LocalMux I__6678 (
            .O(N__36616),
            .I(\pid_front.pid_preregZ0Z_6 ));
    InMux I__6677 (
            .O(N__36609),
            .I(\pid_front.un1_pid_prereg_cry_3 ));
    InMux I__6676 (
            .O(N__36606),
            .I(N__36602));
    InMux I__6675 (
            .O(N__36605),
            .I(N__36599));
    LocalMux I__6674 (
            .O(N__36602),
            .I(\pid_front.error_d_reg_esr_RNIIFUFZ0Z_6 ));
    LocalMux I__6673 (
            .O(N__36599),
            .I(\pid_front.error_d_reg_esr_RNIIFUFZ0Z_6 ));
    CascadeMux I__6672 (
            .O(N__36594),
            .I(N__36591));
    InMux I__6671 (
            .O(N__36591),
            .I(N__36588));
    LocalMux I__6670 (
            .O(N__36588),
            .I(\pid_front.error_p_reg_esr_RNI94TVZ0Z_6 ));
    InMux I__6669 (
            .O(N__36585),
            .I(N__36582));
    LocalMux I__6668 (
            .O(N__36582),
            .I(N__36577));
    CascadeMux I__6667 (
            .O(N__36581),
            .I(N__36574));
    CascadeMux I__6666 (
            .O(N__36580),
            .I(N__36571));
    Span4Mux_h I__6665 (
            .O(N__36577),
            .I(N__36568));
    InMux I__6664 (
            .O(N__36574),
            .I(N__36565));
    InMux I__6663 (
            .O(N__36571),
            .I(N__36562));
    Odrv4 I__6662 (
            .O(N__36568),
            .I(\pid_front.pid_preregZ0Z_7 ));
    LocalMux I__6661 (
            .O(N__36565),
            .I(\pid_front.pid_preregZ0Z_7 ));
    LocalMux I__6660 (
            .O(N__36562),
            .I(\pid_front.pid_preregZ0Z_7 ));
    InMux I__6659 (
            .O(N__36555),
            .I(\pid_front.un1_pid_prereg_cry_4 ));
    InMux I__6658 (
            .O(N__36552),
            .I(N__36549));
    LocalMux I__6657 (
            .O(N__36549),
            .I(N__36546));
    Span4Mux_h I__6656 (
            .O(N__36546),
            .I(N__36543));
    Odrv4 I__6655 (
            .O(N__36543),
            .I(\pid_front.error_p_reg_esr_RNIJETVZ0Z_7 ));
    CascadeMux I__6654 (
            .O(N__36540),
            .I(N__36537));
    InMux I__6653 (
            .O(N__36537),
            .I(N__36534));
    LocalMux I__6652 (
            .O(N__36534),
            .I(N__36531));
    Span4Mux_h I__6651 (
            .O(N__36531),
            .I(N__36528));
    Odrv4 I__6650 (
            .O(N__36528),
            .I(\pid_front.error_d_reg_esr_RNINKUFZ0Z_7 ));
    InMux I__6649 (
            .O(N__36525),
            .I(N__36521));
    InMux I__6648 (
            .O(N__36524),
            .I(N__36518));
    LocalMux I__6647 (
            .O(N__36521),
            .I(N__36515));
    LocalMux I__6646 (
            .O(N__36518),
            .I(N__36511));
    Span4Mux_h I__6645 (
            .O(N__36515),
            .I(N__36508));
    InMux I__6644 (
            .O(N__36514),
            .I(N__36505));
    Span4Mux_h I__6643 (
            .O(N__36511),
            .I(N__36502));
    Odrv4 I__6642 (
            .O(N__36508),
            .I(\pid_front.pid_preregZ0Z_8 ));
    LocalMux I__6641 (
            .O(N__36505),
            .I(\pid_front.pid_preregZ0Z_8 ));
    Odrv4 I__6640 (
            .O(N__36502),
            .I(\pid_front.pid_preregZ0Z_8 ));
    InMux I__6639 (
            .O(N__36495),
            .I(bfn_12_22_0_));
    InMux I__6638 (
            .O(N__36492),
            .I(N__36489));
    LocalMux I__6637 (
            .O(N__36489),
            .I(N__36485));
    InMux I__6636 (
            .O(N__36488),
            .I(N__36482));
    Span4Mux_v I__6635 (
            .O(N__36485),
            .I(N__36479));
    LocalMux I__6634 (
            .O(N__36482),
            .I(\pid_front.error_d_reg_esr_RNISPUFZ0Z_8 ));
    Odrv4 I__6633 (
            .O(N__36479),
            .I(\pid_front.error_d_reg_esr_RNISPUFZ0Z_8 ));
    CascadeMux I__6632 (
            .O(N__36474),
            .I(N__36471));
    InMux I__6631 (
            .O(N__36471),
            .I(N__36468));
    LocalMux I__6630 (
            .O(N__36468),
            .I(N__36465));
    Span4Mux_h I__6629 (
            .O(N__36465),
            .I(N__36462));
    Odrv4 I__6628 (
            .O(N__36462),
            .I(\pid_front.error_p_reg_esr_RNITOTVZ0Z_8 ));
    InMux I__6627 (
            .O(N__36459),
            .I(N__36456));
    LocalMux I__6626 (
            .O(N__36456),
            .I(N__36453));
    Span4Mux_h I__6625 (
            .O(N__36453),
            .I(N__36448));
    InMux I__6624 (
            .O(N__36452),
            .I(N__36445));
    InMux I__6623 (
            .O(N__36451),
            .I(N__36442));
    Odrv4 I__6622 (
            .O(N__36448),
            .I(\pid_front.pid_preregZ0Z_9 ));
    LocalMux I__6621 (
            .O(N__36445),
            .I(\pid_front.pid_preregZ0Z_9 ));
    LocalMux I__6620 (
            .O(N__36442),
            .I(\pid_front.pid_preregZ0Z_9 ));
    InMux I__6619 (
            .O(N__36435),
            .I(\pid_front.un1_pid_prereg_cry_6 ));
    InMux I__6618 (
            .O(N__36432),
            .I(N__36429));
    LocalMux I__6617 (
            .O(N__36429),
            .I(N__36426));
    Span4Mux_h I__6616 (
            .O(N__36426),
            .I(N__36423));
    Odrv4 I__6615 (
            .O(N__36423),
            .I(\pid_front.error_d_reg_esr_RNISPQT1Z0Z_10 ));
    CascadeMux I__6614 (
            .O(N__36420),
            .I(N__36416));
    CascadeMux I__6613 (
            .O(N__36419),
            .I(N__36413));
    InMux I__6612 (
            .O(N__36416),
            .I(N__36410));
    InMux I__6611 (
            .O(N__36413),
            .I(N__36407));
    LocalMux I__6610 (
            .O(N__36410),
            .I(N__36404));
    LocalMux I__6609 (
            .O(N__36407),
            .I(N__36401));
    Span4Mux_h I__6608 (
            .O(N__36404),
            .I(N__36398));
    Span4Mux_v I__6607 (
            .O(N__36401),
            .I(N__36395));
    Span4Mux_v I__6606 (
            .O(N__36398),
            .I(N__36392));
    Span4Mux_h I__6605 (
            .O(N__36395),
            .I(N__36389));
    Span4Mux_v I__6604 (
            .O(N__36392),
            .I(N__36386));
    Span4Mux_h I__6603 (
            .O(N__36389),
            .I(N__36383));
    Odrv4 I__6602 (
            .O(N__36386),
            .I(\pid_front.error_d_reg_esr_RNI1VUFZ0Z_9 ));
    Odrv4 I__6601 (
            .O(N__36383),
            .I(\pid_front.error_d_reg_esr_RNI1VUFZ0Z_9 ));
    InMux I__6600 (
            .O(N__36378),
            .I(N__36375));
    LocalMux I__6599 (
            .O(N__36375),
            .I(N__36372));
    Span4Mux_h I__6598 (
            .O(N__36372),
            .I(N__36366));
    InMux I__6597 (
            .O(N__36371),
            .I(N__36359));
    InMux I__6596 (
            .O(N__36370),
            .I(N__36359));
    InMux I__6595 (
            .O(N__36369),
            .I(N__36359));
    Odrv4 I__6594 (
            .O(N__36366),
            .I(\pid_front.pid_preregZ0Z_10 ));
    LocalMux I__6593 (
            .O(N__36359),
            .I(\pid_front.pid_preregZ0Z_10 ));
    CEMux I__6592 (
            .O(N__36354),
            .I(N__36351));
    LocalMux I__6591 (
            .O(N__36351),
            .I(N__36348));
    Span4Mux_v I__6590 (
            .O(N__36348),
            .I(N__36345));
    Span4Mux_h I__6589 (
            .O(N__36345),
            .I(N__36342));
    Odrv4 I__6588 (
            .O(N__36342),
            .I(\dron_frame_decoder_1.N_489_0 ));
    InMux I__6587 (
            .O(N__36339),
            .I(\pid_front.un1_pid_prereg_cry_0 ));
    InMux I__6586 (
            .O(N__36336),
            .I(N__36332));
    CascadeMux I__6585 (
            .O(N__36335),
            .I(N__36329));
    LocalMux I__6584 (
            .O(N__36332),
            .I(N__36326));
    InMux I__6583 (
            .O(N__36329),
            .I(N__36323));
    Span4Mux_v I__6582 (
            .O(N__36326),
            .I(N__36320));
    LocalMux I__6581 (
            .O(N__36323),
            .I(\pid_front.pid_preregZ0Z_2 ));
    Odrv4 I__6580 (
            .O(N__36320),
            .I(\pid_front.pid_preregZ0Z_2 ));
    InMux I__6579 (
            .O(N__36315),
            .I(\pid_front.un1_pid_prereg_cry_1 ));
    InMux I__6578 (
            .O(N__36312),
            .I(N__36306));
    InMux I__6577 (
            .O(N__36311),
            .I(N__36306));
    LocalMux I__6576 (
            .O(N__36306),
            .I(N__36303));
    Span4Mux_v I__6575 (
            .O(N__36303),
            .I(N__36300));
    Sp12to4 I__6574 (
            .O(N__36300),
            .I(N__36297));
    Odrv12 I__6573 (
            .O(N__36297),
            .I(\pid_front.error_p_regZ0Z_3 ));
    CascadeMux I__6572 (
            .O(N__36294),
            .I(\pid_front.un1_pid_prereg_2_cascade_ ));
    InMux I__6571 (
            .O(N__36291),
            .I(N__36285));
    InMux I__6570 (
            .O(N__36290),
            .I(N__36285));
    LocalMux I__6569 (
            .O(N__36285),
            .I(\pid_front.un1_pid_prereg_0 ));
    CascadeMux I__6568 (
            .O(N__36282),
            .I(N__36279));
    InMux I__6567 (
            .O(N__36279),
            .I(N__36273));
    InMux I__6566 (
            .O(N__36278),
            .I(N__36273));
    LocalMux I__6565 (
            .O(N__36273),
            .I(\pid_front.un1_pid_prereg_2 ));
    CascadeMux I__6564 (
            .O(N__36270),
            .I(\pid_front.un1_pid_prereg_0_cascade_ ));
    CascadeMux I__6563 (
            .O(N__36267),
            .I(N__36264));
    InMux I__6562 (
            .O(N__36264),
            .I(N__36258));
    InMux I__6561 (
            .O(N__36263),
            .I(N__36258));
    LocalMux I__6560 (
            .O(N__36258),
            .I(\pid_front.error_d_reg_prevZ0Z_3 ));
    InMux I__6559 (
            .O(N__36255),
            .I(N__36252));
    LocalMux I__6558 (
            .O(N__36252),
            .I(drone_H_disp_front_1));
    InMux I__6557 (
            .O(N__36249),
            .I(N__36245));
    InMux I__6556 (
            .O(N__36248),
            .I(N__36242));
    LocalMux I__6555 (
            .O(N__36245),
            .I(N__36237));
    LocalMux I__6554 (
            .O(N__36242),
            .I(N__36237));
    Span4Mux_v I__6553 (
            .O(N__36237),
            .I(N__36234));
    Span4Mux_h I__6552 (
            .O(N__36234),
            .I(N__36231));
    Odrv4 I__6551 (
            .O(N__36231),
            .I(throttle_order_0));
    InMux I__6550 (
            .O(N__36228),
            .I(N__36225));
    LocalMux I__6549 (
            .O(N__36225),
            .I(N__36222));
    Odrv4 I__6548 (
            .O(N__36222),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    InMux I__6547 (
            .O(N__36219),
            .I(N__36216));
    LocalMux I__6546 (
            .O(N__36216),
            .I(N__36211));
    CascadeMux I__6545 (
            .O(N__36215),
            .I(N__36208));
    InMux I__6544 (
            .O(N__36214),
            .I(N__36205));
    Span4Mux_h I__6543 (
            .O(N__36211),
            .I(N__36202));
    InMux I__6542 (
            .O(N__36208),
            .I(N__36199));
    LocalMux I__6541 (
            .O(N__36205),
            .I(N__36196));
    Span4Mux_h I__6540 (
            .O(N__36202),
            .I(N__36193));
    LocalMux I__6539 (
            .O(N__36199),
            .I(throttle_order_7));
    Odrv12 I__6538 (
            .O(N__36196),
            .I(throttle_order_7));
    Odrv4 I__6537 (
            .O(N__36193),
            .I(throttle_order_7));
    InMux I__6536 (
            .O(N__36186),
            .I(N__36183));
    LocalMux I__6535 (
            .O(N__36183),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__6534 (
            .O(N__36180),
            .I(N__36177));
    LocalMux I__6533 (
            .O(N__36177),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__6532 (
            .O(N__36174),
            .I(N__36171));
    LocalMux I__6531 (
            .O(N__36171),
            .I(N__36167));
    InMux I__6530 (
            .O(N__36170),
            .I(N__36164));
    Span4Mux_h I__6529 (
            .O(N__36167),
            .I(N__36161));
    LocalMux I__6528 (
            .O(N__36164),
            .I(N__36158));
    Odrv4 I__6527 (
            .O(N__36161),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    Odrv12 I__6526 (
            .O(N__36158),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    InMux I__6525 (
            .O(N__36153),
            .I(N__36149));
    InMux I__6524 (
            .O(N__36152),
            .I(N__36145));
    LocalMux I__6523 (
            .O(N__36149),
            .I(N__36142));
    InMux I__6522 (
            .O(N__36148),
            .I(N__36139));
    LocalMux I__6521 (
            .O(N__36145),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    Odrv4 I__6520 (
            .O(N__36142),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    LocalMux I__6519 (
            .O(N__36139),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    InMux I__6518 (
            .O(N__36132),
            .I(N__36129));
    LocalMux I__6517 (
            .O(N__36129),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    InMux I__6516 (
            .O(N__36126),
            .I(N__36121));
    InMux I__6515 (
            .O(N__36125),
            .I(N__36118));
    CascadeMux I__6514 (
            .O(N__36124),
            .I(N__36115));
    LocalMux I__6513 (
            .O(N__36121),
            .I(N__36110));
    LocalMux I__6512 (
            .O(N__36118),
            .I(N__36110));
    InMux I__6511 (
            .O(N__36115),
            .I(N__36107));
    Span4Mux_v I__6510 (
            .O(N__36110),
            .I(N__36104));
    LocalMux I__6509 (
            .O(N__36107),
            .I(N__36099));
    Span4Mux_h I__6508 (
            .O(N__36104),
            .I(N__36099));
    Odrv4 I__6507 (
            .O(N__36099),
            .I(throttle_order_6));
    InMux I__6506 (
            .O(N__36096),
            .I(N__36093));
    LocalMux I__6505 (
            .O(N__36093),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    InMux I__6504 (
            .O(N__36090),
            .I(N__36087));
    LocalMux I__6503 (
            .O(N__36087),
            .I(N__36083));
    InMux I__6502 (
            .O(N__36086),
            .I(N__36080));
    Span4Mux_v I__6501 (
            .O(N__36083),
            .I(N__36077));
    LocalMux I__6500 (
            .O(N__36080),
            .I(N__36074));
    Sp12to4 I__6499 (
            .O(N__36077),
            .I(N__36069));
    Span12Mux_v I__6498 (
            .O(N__36074),
            .I(N__36069));
    Odrv12 I__6497 (
            .O(N__36069),
            .I(throttle_order_3));
    InMux I__6496 (
            .O(N__36066),
            .I(N__36062));
    InMux I__6495 (
            .O(N__36065),
            .I(N__36059));
    LocalMux I__6494 (
            .O(N__36062),
            .I(N__36053));
    LocalMux I__6493 (
            .O(N__36059),
            .I(N__36053));
    CascadeMux I__6492 (
            .O(N__36058),
            .I(N__36050));
    Span4Mux_h I__6491 (
            .O(N__36053),
            .I(N__36047));
    InMux I__6490 (
            .O(N__36050),
            .I(N__36044));
    Span4Mux_h I__6489 (
            .O(N__36047),
            .I(N__36041));
    LocalMux I__6488 (
            .O(N__36044),
            .I(throttle_order_9));
    Odrv4 I__6487 (
            .O(N__36041),
            .I(throttle_order_9));
    InMux I__6486 (
            .O(N__36036),
            .I(N__36033));
    LocalMux I__6485 (
            .O(N__36033),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__6484 (
            .O(N__36030),
            .I(N__36027));
    LocalMux I__6483 (
            .O(N__36027),
            .I(N__36024));
    Odrv4 I__6482 (
            .O(N__36024),
            .I(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ));
    CascadeMux I__6481 (
            .O(N__36021),
            .I(N__36017));
    InMux I__6480 (
            .O(N__36020),
            .I(N__36014));
    InMux I__6479 (
            .O(N__36017),
            .I(N__36011));
    LocalMux I__6478 (
            .O(N__36014),
            .I(N__36008));
    LocalMux I__6477 (
            .O(N__36011),
            .I(N__36005));
    Span4Mux_h I__6476 (
            .O(N__36008),
            .I(N__36002));
    Span4Mux_h I__6475 (
            .O(N__36005),
            .I(N__35999));
    Span4Mux_v I__6474 (
            .O(N__36002),
            .I(N__35996));
    Span4Mux_h I__6473 (
            .O(N__35999),
            .I(N__35993));
    Span4Mux_h I__6472 (
            .O(N__35996),
            .I(N__35990));
    Odrv4 I__6471 (
            .O(N__35993),
            .I(throttle_order_4));
    Odrv4 I__6470 (
            .O(N__35990),
            .I(throttle_order_4));
    InMux I__6469 (
            .O(N__35985),
            .I(N__35982));
    LocalMux I__6468 (
            .O(N__35982),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__6467 (
            .O(N__35979),
            .I(N__35975));
    InMux I__6466 (
            .O(N__35978),
            .I(N__35972));
    LocalMux I__6465 (
            .O(N__35975),
            .I(N__35966));
    LocalMux I__6464 (
            .O(N__35972),
            .I(N__35966));
    CascadeMux I__6463 (
            .O(N__35971),
            .I(N__35963));
    Span4Mux_h I__6462 (
            .O(N__35966),
            .I(N__35960));
    InMux I__6461 (
            .O(N__35963),
            .I(N__35957));
    Span4Mux_h I__6460 (
            .O(N__35960),
            .I(N__35954));
    LocalMux I__6459 (
            .O(N__35957),
            .I(throttle_order_8));
    Odrv4 I__6458 (
            .O(N__35954),
            .I(throttle_order_8));
    InMux I__6457 (
            .O(N__35949),
            .I(N__35946));
    LocalMux I__6456 (
            .O(N__35946),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    InMux I__6455 (
            .O(N__35943),
            .I(N__35940));
    LocalMux I__6454 (
            .O(N__35940),
            .I(N__35936));
    InMux I__6453 (
            .O(N__35939),
            .I(N__35933));
    Span4Mux_h I__6452 (
            .O(N__35936),
            .I(N__35928));
    LocalMux I__6451 (
            .O(N__35933),
            .I(N__35928));
    Span4Mux_h I__6450 (
            .O(N__35928),
            .I(N__35925));
    Span4Mux_v I__6449 (
            .O(N__35925),
            .I(N__35922));
    Sp12to4 I__6448 (
            .O(N__35922),
            .I(N__35919));
    Odrv12 I__6447 (
            .O(N__35919),
            .I(throttle_order_12));
    InMux I__6446 (
            .O(N__35916),
            .I(N__35913));
    LocalMux I__6445 (
            .O(N__35913),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    InMux I__6444 (
            .O(N__35910),
            .I(N__35907));
    LocalMux I__6443 (
            .O(N__35907),
            .I(N__35904));
    Odrv4 I__6442 (
            .O(N__35904),
            .I(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ));
    InMux I__6441 (
            .O(N__35901),
            .I(N__35898));
    LocalMux I__6440 (
            .O(N__35898),
            .I(frame_decoder_CH4data_4));
    CascadeMux I__6439 (
            .O(N__35895),
            .I(N__35892));
    InMux I__6438 (
            .O(N__35892),
            .I(N__35889));
    LocalMux I__6437 (
            .O(N__35889),
            .I(N__35886));
    Span4Mux_h I__6436 (
            .O(N__35886),
            .I(N__35883));
    Odrv4 I__6435 (
            .O(N__35883),
            .I(frame_decoder_OFF4data_4));
    InMux I__6434 (
            .O(N__35880),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__6433 (
            .O(N__35877),
            .I(N__35874));
    LocalMux I__6432 (
            .O(N__35874),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__6431 (
            .O(N__35871),
            .I(N__35868));
    InMux I__6430 (
            .O(N__35868),
            .I(N__35865));
    LocalMux I__6429 (
            .O(N__35865),
            .I(N__35862));
    Odrv12 I__6428 (
            .O(N__35862),
            .I(frame_decoder_OFF4data_5));
    InMux I__6427 (
            .O(N__35859),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__6426 (
            .O(N__35856),
            .I(N__35853));
    LocalMux I__6425 (
            .O(N__35853),
            .I(N__35850));
    Odrv4 I__6424 (
            .O(N__35850),
            .I(frame_decoder_OFF4data_6));
    CascadeMux I__6423 (
            .O(N__35847),
            .I(N__35844));
    InMux I__6422 (
            .O(N__35844),
            .I(N__35841));
    LocalMux I__6421 (
            .O(N__35841),
            .I(frame_decoder_CH4data_6));
    InMux I__6420 (
            .O(N__35838),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__6419 (
            .O(N__35835),
            .I(N__35832));
    LocalMux I__6418 (
            .O(N__35832),
            .I(N__35829));
    Span4Mux_v I__6417 (
            .O(N__35829),
            .I(N__35826));
    Span4Mux_h I__6416 (
            .O(N__35826),
            .I(N__35823));
    Odrv4 I__6415 (
            .O(N__35823),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    InMux I__6414 (
            .O(N__35820),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__6413 (
            .O(N__35817),
            .I(bfn_12_13_0_));
    InMux I__6412 (
            .O(N__35814),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    InMux I__6411 (
            .O(N__35811),
            .I(N__35807));
    InMux I__6410 (
            .O(N__35810),
            .I(N__35804));
    LocalMux I__6409 (
            .O(N__35807),
            .I(N__35801));
    LocalMux I__6408 (
            .O(N__35804),
            .I(N__35798));
    Span4Mux_h I__6407 (
            .O(N__35801),
            .I(N__35795));
    Span12Mux_v I__6406 (
            .O(N__35798),
            .I(N__35792));
    Odrv4 I__6405 (
            .O(N__35795),
            .I(frame_decoder_OFF4data_7));
    Odrv12 I__6404 (
            .O(N__35792),
            .I(frame_decoder_OFF4data_7));
    InMux I__6403 (
            .O(N__35787),
            .I(N__35784));
    LocalMux I__6402 (
            .O(N__35784),
            .I(N__35780));
    InMux I__6401 (
            .O(N__35783),
            .I(N__35777));
    Span4Mux_v I__6400 (
            .O(N__35780),
            .I(N__35774));
    LocalMux I__6399 (
            .O(N__35777),
            .I(N__35769));
    Span4Mux_h I__6398 (
            .O(N__35774),
            .I(N__35769));
    Odrv4 I__6397 (
            .O(N__35769),
            .I(frame_decoder_CH4data_7));
    InMux I__6396 (
            .O(N__35766),
            .I(N__35763));
    LocalMux I__6395 (
            .O(N__35763),
            .I(\scaler_4.N_1849_i_l_ofxZ0 ));
    CEMux I__6394 (
            .O(N__35760),
            .I(N__35757));
    LocalMux I__6393 (
            .O(N__35757),
            .I(N__35754));
    Span4Mux_h I__6392 (
            .O(N__35754),
            .I(N__35751));
    Odrv4 I__6391 (
            .O(N__35751),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__6390 (
            .O(N__35748),
            .I(N__35745));
    LocalMux I__6389 (
            .O(N__35745),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__6388 (
            .O(N__35742),
            .I(N__35739));
    InMux I__6387 (
            .O(N__35739),
            .I(N__35736));
    LocalMux I__6386 (
            .O(N__35736),
            .I(N__35733));
    Odrv4 I__6385 (
            .O(N__35733),
            .I(frame_decoder_OFF4data_1));
    InMux I__6384 (
            .O(N__35730),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__6383 (
            .O(N__35727),
            .I(N__35724));
    LocalMux I__6382 (
            .O(N__35724),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__6381 (
            .O(N__35721),
            .I(N__35718));
    InMux I__6380 (
            .O(N__35718),
            .I(N__35715));
    LocalMux I__6379 (
            .O(N__35715),
            .I(N__35712));
    Odrv4 I__6378 (
            .O(N__35712),
            .I(frame_decoder_OFF4data_2));
    InMux I__6377 (
            .O(N__35709),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__6376 (
            .O(N__35706),
            .I(N__35703));
    LocalMux I__6375 (
            .O(N__35703),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__6374 (
            .O(N__35700),
            .I(N__35697));
    InMux I__6373 (
            .O(N__35697),
            .I(N__35694));
    LocalMux I__6372 (
            .O(N__35694),
            .I(N__35691));
    Odrv4 I__6371 (
            .O(N__35691),
            .I(frame_decoder_OFF4data_3));
    InMux I__6370 (
            .O(N__35688),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__6369 (
            .O(N__35685),
            .I(N__35679));
    InMux I__6368 (
            .O(N__35684),
            .I(N__35679));
    LocalMux I__6367 (
            .O(N__35679),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    InMux I__6366 (
            .O(N__35676),
            .I(N__35671));
    InMux I__6365 (
            .O(N__35675),
            .I(N__35666));
    InMux I__6364 (
            .O(N__35674),
            .I(N__35666));
    LocalMux I__6363 (
            .O(N__35671),
            .I(\pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11 ));
    LocalMux I__6362 (
            .O(N__35666),
            .I(\pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11 ));
    InMux I__6361 (
            .O(N__35661),
            .I(N__35658));
    LocalMux I__6360 (
            .O(N__35658),
            .I(N__35654));
    InMux I__6359 (
            .O(N__35657),
            .I(N__35651));
    Odrv4 I__6358 (
            .O(N__35654),
            .I(\pid_front.error_p_reg_esr_RNI653NZ0Z_10 ));
    LocalMux I__6357 (
            .O(N__35651),
            .I(\pid_front.error_p_reg_esr_RNI653NZ0Z_10 ));
    InMux I__6356 (
            .O(N__35646),
            .I(N__35642));
    InMux I__6355 (
            .O(N__35645),
            .I(N__35639));
    LocalMux I__6354 (
            .O(N__35642),
            .I(\pid_front.N_1463_i ));
    LocalMux I__6353 (
            .O(N__35639),
            .I(\pid_front.N_1463_i ));
    InMux I__6352 (
            .O(N__35634),
            .I(N__35630));
    InMux I__6351 (
            .O(N__35633),
            .I(N__35627));
    LocalMux I__6350 (
            .O(N__35630),
            .I(N__35622));
    LocalMux I__6349 (
            .O(N__35627),
            .I(N__35622));
    Span4Mux_v I__6348 (
            .O(N__35622),
            .I(N__35619));
    Odrv4 I__6347 (
            .O(N__35619),
            .I(\pid_front.error_p_reg_esr_RNIM6G7Z0Z_9 ));
    InMux I__6346 (
            .O(N__35616),
            .I(N__35612));
    InMux I__6345 (
            .O(N__35615),
            .I(N__35609));
    LocalMux I__6344 (
            .O(N__35612),
            .I(N__35604));
    LocalMux I__6343 (
            .O(N__35609),
            .I(N__35601));
    InMux I__6342 (
            .O(N__35608),
            .I(N__35596));
    InMux I__6341 (
            .O(N__35607),
            .I(N__35596));
    Span4Mux_h I__6340 (
            .O(N__35604),
            .I(N__35591));
    Span4Mux_h I__6339 (
            .O(N__35601),
            .I(N__35591));
    LocalMux I__6338 (
            .O(N__35596),
            .I(\uart_drone.N_152 ));
    Odrv4 I__6337 (
            .O(N__35591),
            .I(\uart_drone.N_152 ));
    IoInMux I__6336 (
            .O(N__35586),
            .I(N__35583));
    LocalMux I__6335 (
            .O(N__35583),
            .I(N__35580));
    Odrv12 I__6334 (
            .O(N__35580),
            .I(\pid_side.state_0_0 ));
    InMux I__6333 (
            .O(N__35577),
            .I(N__35573));
    InMux I__6332 (
            .O(N__35576),
            .I(N__35568));
    LocalMux I__6331 (
            .O(N__35573),
            .I(N__35565));
    CascadeMux I__6330 (
            .O(N__35572),
            .I(N__35561));
    CascadeMux I__6329 (
            .O(N__35571),
            .I(N__35556));
    LocalMux I__6328 (
            .O(N__35568),
            .I(N__35553));
    Span4Mux_v I__6327 (
            .O(N__35565),
            .I(N__35550));
    InMux I__6326 (
            .O(N__35564),
            .I(N__35547));
    InMux I__6325 (
            .O(N__35561),
            .I(N__35542));
    InMux I__6324 (
            .O(N__35560),
            .I(N__35542));
    InMux I__6323 (
            .O(N__35559),
            .I(N__35539));
    InMux I__6322 (
            .O(N__35556),
            .I(N__35534));
    Span4Mux_v I__6321 (
            .O(N__35553),
            .I(N__35531));
    Span4Mux_h I__6320 (
            .O(N__35550),
            .I(N__35526));
    LocalMux I__6319 (
            .O(N__35547),
            .I(N__35526));
    LocalMux I__6318 (
            .O(N__35542),
            .I(N__35521));
    LocalMux I__6317 (
            .O(N__35539),
            .I(N__35521));
    InMux I__6316 (
            .O(N__35538),
            .I(N__35518));
    InMux I__6315 (
            .O(N__35537),
            .I(N__35515));
    LocalMux I__6314 (
            .O(N__35534),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__6313 (
            .O(N__35531),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__6312 (
            .O(N__35526),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__6311 (
            .O(N__35521),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    LocalMux I__6310 (
            .O(N__35518),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    LocalMux I__6309 (
            .O(N__35515),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__6308 (
            .O(N__35502),
            .I(N__35499));
    LocalMux I__6307 (
            .O(N__35499),
            .I(N__35494));
    InMux I__6306 (
            .O(N__35498),
            .I(N__35491));
    InMux I__6305 (
            .O(N__35497),
            .I(N__35488));
    Span4Mux_h I__6304 (
            .O(N__35494),
            .I(N__35480));
    LocalMux I__6303 (
            .O(N__35491),
            .I(N__35477));
    LocalMux I__6302 (
            .O(N__35488),
            .I(N__35474));
    InMux I__6301 (
            .O(N__35487),
            .I(N__35469));
    InMux I__6300 (
            .O(N__35486),
            .I(N__35469));
    InMux I__6299 (
            .O(N__35485),
            .I(N__35466));
    InMux I__6298 (
            .O(N__35484),
            .I(N__35459));
    InMux I__6297 (
            .O(N__35483),
            .I(N__35459));
    Span4Mux_v I__6296 (
            .O(N__35480),
            .I(N__35456));
    Span4Mux_v I__6295 (
            .O(N__35477),
            .I(N__35447));
    Span4Mux_h I__6294 (
            .O(N__35474),
            .I(N__35447));
    LocalMux I__6293 (
            .O(N__35469),
            .I(N__35447));
    LocalMux I__6292 (
            .O(N__35466),
            .I(N__35447));
    InMux I__6291 (
            .O(N__35465),
            .I(N__35444));
    InMux I__6290 (
            .O(N__35464),
            .I(N__35441));
    LocalMux I__6289 (
            .O(N__35459),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__6288 (
            .O(N__35456),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__6287 (
            .O(N__35447),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__6286 (
            .O(N__35444),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__6285 (
            .O(N__35441),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    CascadeMux I__6284 (
            .O(N__35430),
            .I(N__35427));
    InMux I__6283 (
            .O(N__35427),
            .I(N__35423));
    CascadeMux I__6282 (
            .O(N__35426),
            .I(N__35416));
    LocalMux I__6281 (
            .O(N__35423),
            .I(N__35413));
    InMux I__6280 (
            .O(N__35422),
            .I(N__35410));
    InMux I__6279 (
            .O(N__35421),
            .I(N__35401));
    InMux I__6278 (
            .O(N__35420),
            .I(N__35401));
    InMux I__6277 (
            .O(N__35419),
            .I(N__35398));
    InMux I__6276 (
            .O(N__35416),
            .I(N__35395));
    Span4Mux_h I__6275 (
            .O(N__35413),
            .I(N__35390));
    LocalMux I__6274 (
            .O(N__35410),
            .I(N__35390));
    InMux I__6273 (
            .O(N__35409),
            .I(N__35384));
    InMux I__6272 (
            .O(N__35408),
            .I(N__35384));
    InMux I__6271 (
            .O(N__35407),
            .I(N__35381));
    InMux I__6270 (
            .O(N__35406),
            .I(N__35378));
    LocalMux I__6269 (
            .O(N__35401),
            .I(N__35375));
    LocalMux I__6268 (
            .O(N__35398),
            .I(N__35370));
    LocalMux I__6267 (
            .O(N__35395),
            .I(N__35370));
    Span4Mux_v I__6266 (
            .O(N__35390),
            .I(N__35367));
    InMux I__6265 (
            .O(N__35389),
            .I(N__35364));
    LocalMux I__6264 (
            .O(N__35384),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__6263 (
            .O(N__35381),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__6262 (
            .O(N__35378),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__6261 (
            .O(N__35375),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__6260 (
            .O(N__35370),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__6259 (
            .O(N__35367),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__6258 (
            .O(N__35364),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    InMux I__6257 (
            .O(N__35349),
            .I(N__35346));
    LocalMux I__6256 (
            .O(N__35346),
            .I(N__35343));
    Odrv4 I__6255 (
            .O(N__35343),
            .I(\uart_drone.data_Auxce_0_3 ));
    CascadeMux I__6254 (
            .O(N__35340),
            .I(\pid_front.m9_e_4_cascade_ ));
    InMux I__6253 (
            .O(N__35337),
            .I(N__35334));
    LocalMux I__6252 (
            .O(N__35334),
            .I(\pid_front.m9_e_5 ));
    CascadeMux I__6251 (
            .O(N__35331),
            .I(N__35327));
    InMux I__6250 (
            .O(N__35330),
            .I(N__35322));
    InMux I__6249 (
            .O(N__35327),
            .I(N__35319));
    InMux I__6248 (
            .O(N__35326),
            .I(N__35313));
    InMux I__6247 (
            .O(N__35325),
            .I(N__35313));
    LocalMux I__6246 (
            .O(N__35322),
            .I(N__35308));
    LocalMux I__6245 (
            .O(N__35319),
            .I(N__35308));
    InMux I__6244 (
            .O(N__35318),
            .I(N__35305));
    LocalMux I__6243 (
            .O(N__35313),
            .I(\pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20 ));
    Odrv4 I__6242 (
            .O(N__35308),
            .I(\pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20 ));
    LocalMux I__6241 (
            .O(N__35305),
            .I(\pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20 ));
    InMux I__6240 (
            .O(N__35298),
            .I(N__35291));
    InMux I__6239 (
            .O(N__35297),
            .I(N__35291));
    InMux I__6238 (
            .O(N__35296),
            .I(N__35288));
    LocalMux I__6237 (
            .O(N__35291),
            .I(N__35285));
    LocalMux I__6236 (
            .O(N__35288),
            .I(\pid_front.pid_prereg_esr_RNIVDO51Z0Z_10 ));
    Odrv12 I__6235 (
            .O(N__35285),
            .I(\pid_front.pid_prereg_esr_RNIVDO51Z0Z_10 ));
    InMux I__6234 (
            .O(N__35280),
            .I(N__35277));
    LocalMux I__6233 (
            .O(N__35277),
            .I(N__35266));
    InMux I__6232 (
            .O(N__35276),
            .I(N__35253));
    InMux I__6231 (
            .O(N__35275),
            .I(N__35253));
    InMux I__6230 (
            .O(N__35274),
            .I(N__35253));
    InMux I__6229 (
            .O(N__35273),
            .I(N__35253));
    InMux I__6228 (
            .O(N__35272),
            .I(N__35253));
    InMux I__6227 (
            .O(N__35271),
            .I(N__35253));
    InMux I__6226 (
            .O(N__35270),
            .I(N__35248));
    InMux I__6225 (
            .O(N__35269),
            .I(N__35248));
    Odrv12 I__6224 (
            .O(N__35266),
            .I(\pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12 ));
    LocalMux I__6223 (
            .O(N__35253),
            .I(\pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12 ));
    LocalMux I__6222 (
            .O(N__35248),
            .I(\pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12 ));
    InMux I__6221 (
            .O(N__35241),
            .I(N__35238));
    LocalMux I__6220 (
            .O(N__35238),
            .I(N__35235));
    Span4Mux_v I__6219 (
            .O(N__35235),
            .I(N__35230));
    InMux I__6218 (
            .O(N__35234),
            .I(N__35225));
    InMux I__6217 (
            .O(N__35233),
            .I(N__35225));
    Odrv4 I__6216 (
            .O(N__35230),
            .I(\pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13 ));
    LocalMux I__6215 (
            .O(N__35225),
            .I(\pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13 ));
    CEMux I__6214 (
            .O(N__35220),
            .I(N__35216));
    CEMux I__6213 (
            .O(N__35219),
            .I(N__35213));
    LocalMux I__6212 (
            .O(N__35216),
            .I(N__35210));
    LocalMux I__6211 (
            .O(N__35213),
            .I(N__35206));
    Span4Mux_v I__6210 (
            .O(N__35210),
            .I(N__35203));
    CEMux I__6209 (
            .O(N__35209),
            .I(N__35200));
    Odrv4 I__6208 (
            .O(N__35206),
            .I(\pid_front.state_0_1 ));
    Odrv4 I__6207 (
            .O(N__35203),
            .I(\pid_front.state_0_1 ));
    LocalMux I__6206 (
            .O(N__35200),
            .I(\pid_front.state_0_1 ));
    SRMux I__6205 (
            .O(N__35193),
            .I(N__35190));
    LocalMux I__6204 (
            .O(N__35190),
            .I(N__35184));
    SRMux I__6203 (
            .O(N__35189),
            .I(N__35181));
    SRMux I__6202 (
            .O(N__35188),
            .I(N__35178));
    SRMux I__6201 (
            .O(N__35187),
            .I(N__35175));
    Span4Mux_v I__6200 (
            .O(N__35184),
            .I(N__35170));
    LocalMux I__6199 (
            .O(N__35181),
            .I(N__35170));
    LocalMux I__6198 (
            .O(N__35178),
            .I(N__35163));
    LocalMux I__6197 (
            .O(N__35175),
            .I(N__35163));
    Span4Mux_h I__6196 (
            .O(N__35170),
            .I(N__35163));
    Odrv4 I__6195 (
            .O(N__35163),
            .I(\pid_front.un1_reset_0_i ));
    CascadeMux I__6194 (
            .O(N__35160),
            .I(\pid_front.state_RNIVIRQZ0Z_0_cascade_ ));
    CascadeMux I__6193 (
            .O(N__35157),
            .I(N__35154));
    InMux I__6192 (
            .O(N__35154),
            .I(N__35148));
    InMux I__6191 (
            .O(N__35153),
            .I(N__35148));
    LocalMux I__6190 (
            .O(N__35148),
            .I(N__35145));
    Span4Mux_v I__6189 (
            .O(N__35145),
            .I(N__35142));
    Span4Mux_v I__6188 (
            .O(N__35142),
            .I(N__35139));
    Sp12to4 I__6187 (
            .O(N__35139),
            .I(N__35136));
    Odrv12 I__6186 (
            .O(N__35136),
            .I(\pid_front.error_p_regZ0Z_10 ));
    CascadeMux I__6185 (
            .O(N__35133),
            .I(\pid_front.error_p_reg_esr_RNI653NZ0Z_10_cascade_ ));
    InMux I__6184 (
            .O(N__35130),
            .I(N__35125));
    InMux I__6183 (
            .O(N__35129),
            .I(N__35120));
    InMux I__6182 (
            .O(N__35128),
            .I(N__35120));
    LocalMux I__6181 (
            .O(N__35125),
            .I(N__35114));
    LocalMux I__6180 (
            .O(N__35120),
            .I(N__35114));
    InMux I__6179 (
            .O(N__35119),
            .I(N__35111));
    Odrv4 I__6178 (
            .O(N__35114),
            .I(\pid_front.error_d_reg_prevZ0Z_7 ));
    LocalMux I__6177 (
            .O(N__35111),
            .I(\pid_front.error_d_reg_prevZ0Z_7 ));
    CascadeMux I__6176 (
            .O(N__35106),
            .I(\pid_front.m26_e_5_cascade_ ));
    CascadeMux I__6175 (
            .O(N__35103),
            .I(\pid_front.m26_e_1_cascade_ ));
    InMux I__6174 (
            .O(N__35100),
            .I(N__35097));
    LocalMux I__6173 (
            .O(N__35097),
            .I(\pid_front.m26_e_5 ));
    CascadeMux I__6172 (
            .O(N__35094),
            .I(N__35091));
    InMux I__6171 (
            .O(N__35091),
            .I(N__35088));
    LocalMux I__6170 (
            .O(N__35088),
            .I(\pid_front.pid_prereg_esr_RNIGSMQ1Z0Z_10 ));
    InMux I__6169 (
            .O(N__35085),
            .I(N__35082));
    LocalMux I__6168 (
            .O(N__35082),
            .I(N__35079));
    Odrv4 I__6167 (
            .O(N__35079),
            .I(\pid_front.m18_s_5 ));
    InMux I__6166 (
            .O(N__35076),
            .I(N__35073));
    LocalMux I__6165 (
            .O(N__35073),
            .I(N__35070));
    Odrv4 I__6164 (
            .O(N__35070),
            .I(\pid_front.m18_s_4 ));
    InMux I__6163 (
            .O(N__35067),
            .I(N__35058));
    InMux I__6162 (
            .O(N__35066),
            .I(N__35058));
    InMux I__6161 (
            .O(N__35065),
            .I(N__35058));
    LocalMux I__6160 (
            .O(N__35058),
            .I(\pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5 ));
    InMux I__6159 (
            .O(N__35055),
            .I(N__35043));
    InMux I__6158 (
            .O(N__35054),
            .I(N__35043));
    InMux I__6157 (
            .O(N__35053),
            .I(N__35043));
    InMux I__6156 (
            .O(N__35052),
            .I(N__35043));
    LocalMux I__6155 (
            .O(N__35043),
            .I(\pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10 ));
    InMux I__6154 (
            .O(N__35040),
            .I(N__35034));
    InMux I__6153 (
            .O(N__35039),
            .I(N__35031));
    InMux I__6152 (
            .O(N__35038),
            .I(N__35026));
    InMux I__6151 (
            .O(N__35037),
            .I(N__35026));
    LocalMux I__6150 (
            .O(N__35034),
            .I(N__35023));
    LocalMux I__6149 (
            .O(N__35031),
            .I(\pid_front.error_p_regZ0Z_7 ));
    LocalMux I__6148 (
            .O(N__35026),
            .I(\pid_front.error_p_regZ0Z_7 ));
    Odrv4 I__6147 (
            .O(N__35023),
            .I(\pid_front.error_p_regZ0Z_7 ));
    CascadeMux I__6146 (
            .O(N__35016),
            .I(\pid_front.un1_pid_prereg_60_0_cascade_ ));
    CascadeMux I__6145 (
            .O(N__35013),
            .I(\pid_front.N_1447_i_cascade_ ));
    InMux I__6144 (
            .O(N__35010),
            .I(N__35004));
    InMux I__6143 (
            .O(N__35009),
            .I(N__35001));
    InMux I__6142 (
            .O(N__35008),
            .I(N__34996));
    InMux I__6141 (
            .O(N__35007),
            .I(N__34996));
    LocalMux I__6140 (
            .O(N__35004),
            .I(N__34989));
    LocalMux I__6139 (
            .O(N__35001),
            .I(N__34989));
    LocalMux I__6138 (
            .O(N__34996),
            .I(N__34989));
    Span12Mux_h I__6137 (
            .O(N__34989),
            .I(N__34986));
    Odrv12 I__6136 (
            .O(N__34986),
            .I(\pid_front.error_p_regZ0Z_6 ));
    InMux I__6135 (
            .O(N__34983),
            .I(N__34980));
    LocalMux I__6134 (
            .O(N__34980),
            .I(N__34974));
    InMux I__6133 (
            .O(N__34979),
            .I(N__34967));
    InMux I__6132 (
            .O(N__34978),
            .I(N__34967));
    InMux I__6131 (
            .O(N__34977),
            .I(N__34967));
    Odrv4 I__6130 (
            .O(N__34974),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    LocalMux I__6129 (
            .O(N__34967),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    CascadeMux I__6128 (
            .O(N__34962),
            .I(\pid_front.un1_pid_prereg_50_0_cascade_ ));
    InMux I__6127 (
            .O(N__34959),
            .I(N__34956));
    LocalMux I__6126 (
            .O(N__34956),
            .I(drone_altitude_3));
    CEMux I__6125 (
            .O(N__34953),
            .I(N__34950));
    LocalMux I__6124 (
            .O(N__34950),
            .I(N__34947));
    Span4Mux_v I__6123 (
            .O(N__34947),
            .I(N__34943));
    CEMux I__6122 (
            .O(N__34946),
            .I(N__34940));
    Sp12to4 I__6121 (
            .O(N__34943),
            .I(N__34937));
    LocalMux I__6120 (
            .O(N__34940),
            .I(N__34934));
    Span12Mux_s9_h I__6119 (
            .O(N__34937),
            .I(N__34931));
    Span4Mux_v I__6118 (
            .O(N__34934),
            .I(N__34928));
    Odrv12 I__6117 (
            .O(N__34931),
            .I(\dron_frame_decoder_1.N_521_0 ));
    Odrv4 I__6116 (
            .O(N__34928),
            .I(\dron_frame_decoder_1.N_521_0 ));
    InMux I__6115 (
            .O(N__34923),
            .I(N__34920));
    LocalMux I__6114 (
            .O(N__34920),
            .I(N__34917));
    Span12Mux_v I__6113 (
            .O(N__34917),
            .I(N__34914));
    Odrv12 I__6112 (
            .O(N__34914),
            .I(\pid_alt.error_d_reg_prevZ0Z_0 ));
    CascadeMux I__6111 (
            .O(N__34911),
            .I(N__34908));
    InMux I__6110 (
            .O(N__34908),
            .I(N__34905));
    LocalMux I__6109 (
            .O(N__34905),
            .I(N__34901));
    InMux I__6108 (
            .O(N__34904),
            .I(N__34898));
    Span4Mux_v I__6107 (
            .O(N__34901),
            .I(N__34895));
    LocalMux I__6106 (
            .O(N__34898),
            .I(N__34892));
    Sp12to4 I__6105 (
            .O(N__34895),
            .I(N__34887));
    Span12Mux_v I__6104 (
            .O(N__34892),
            .I(N__34887));
    Odrv12 I__6103 (
            .O(N__34887),
            .I(\pid_alt.error_d_reg_prev_i_0 ));
    CascadeMux I__6102 (
            .O(N__34884),
            .I(\pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12_cascade_ ));
    CascadeMux I__6101 (
            .O(N__34881),
            .I(\pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10_cascade_ ));
    CascadeMux I__6100 (
            .O(N__34878),
            .I(\pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5_cascade_ ));
    InMux I__6099 (
            .O(N__34875),
            .I(N__34872));
    LocalMux I__6098 (
            .O(N__34872),
            .I(N__34869));
    Odrv4 I__6097 (
            .O(N__34869),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__6096 (
            .O(N__34866),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__6095 (
            .O(N__34863),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__6094 (
            .O(N__34860),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__6093 (
            .O(N__34857),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__6092 (
            .O(N__34854),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__6091 (
            .O(N__34851),
            .I(\ppm_encoder_1.un1_aileron_cry_13 ));
    InMux I__6090 (
            .O(N__34848),
            .I(N__34845));
    LocalMux I__6089 (
            .O(N__34845),
            .I(N__34842));
    Span12Mux_s7_h I__6088 (
            .O(N__34842),
            .I(N__34839));
    Odrv12 I__6087 (
            .O(N__34839),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__6086 (
            .O(N__34836),
            .I(N__34833));
    LocalMux I__6085 (
            .O(N__34833),
            .I(drone_altitude_2));
    InMux I__6084 (
            .O(N__34830),
            .I(N__34827));
    LocalMux I__6083 (
            .O(N__34827),
            .I(N__34824));
    Span4Mux_h I__6082 (
            .O(N__34824),
            .I(N__34821));
    Span4Mux_h I__6081 (
            .O(N__34821),
            .I(N__34818));
    Odrv4 I__6080 (
            .O(N__34818),
            .I(\pid_alt.error_axbZ0Z_3 ));
    InMux I__6079 (
            .O(N__34815),
            .I(N__34812));
    LocalMux I__6078 (
            .O(N__34812),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__6077 (
            .O(N__34809),
            .I(\ppm_encoder_1.un1_aileron_cry_0 ));
    InMux I__6076 (
            .O(N__34806),
            .I(\ppm_encoder_1.un1_aileron_cry_1 ));
    InMux I__6075 (
            .O(N__34803),
            .I(\ppm_encoder_1.un1_aileron_cry_2 ));
    InMux I__6074 (
            .O(N__34800),
            .I(\ppm_encoder_1.un1_aileron_cry_3 ));
    InMux I__6073 (
            .O(N__34797),
            .I(\ppm_encoder_1.un1_aileron_cry_4 ));
    InMux I__6072 (
            .O(N__34794),
            .I(\ppm_encoder_1.un1_aileron_cry_5 ));
    InMux I__6071 (
            .O(N__34791),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__6070 (
            .O(N__34788),
            .I(bfn_11_18_0_));
    InMux I__6069 (
            .O(N__34785),
            .I(bfn_11_15_0_));
    InMux I__6068 (
            .O(N__34782),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__6067 (
            .O(N__34779),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__6066 (
            .O(N__34776),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__6065 (
            .O(N__34773),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__6064 (
            .O(N__34770),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__6063 (
            .O(N__34767),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    CascadeMux I__6062 (
            .O(N__34764),
            .I(N__34761));
    InMux I__6061 (
            .O(N__34761),
            .I(N__34757));
    InMux I__6060 (
            .O(N__34760),
            .I(N__34754));
    LocalMux I__6059 (
            .O(N__34757),
            .I(N__34751));
    LocalMux I__6058 (
            .O(N__34754),
            .I(N__34748));
    Span4Mux_h I__6057 (
            .O(N__34751),
            .I(N__34745));
    Span4Mux_v I__6056 (
            .O(N__34748),
            .I(N__34742));
    Span4Mux_v I__6055 (
            .O(N__34745),
            .I(N__34737));
    Span4Mux_h I__6054 (
            .O(N__34742),
            .I(N__34737));
    Odrv4 I__6053 (
            .O(N__34737),
            .I(throttle_order_13));
    InMux I__6052 (
            .O(N__34734),
            .I(N__34731));
    LocalMux I__6051 (
            .O(N__34731),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    InMux I__6050 (
            .O(N__34728),
            .I(N__34724));
    InMux I__6049 (
            .O(N__34727),
            .I(N__34721));
    LocalMux I__6048 (
            .O(N__34724),
            .I(N__34718));
    LocalMux I__6047 (
            .O(N__34721),
            .I(N__34714));
    Span4Mux_v I__6046 (
            .O(N__34718),
            .I(N__34711));
    InMux I__6045 (
            .O(N__34717),
            .I(N__34708));
    Span4Mux_h I__6044 (
            .O(N__34714),
            .I(N__34703));
    Span4Mux_h I__6043 (
            .O(N__34711),
            .I(N__34703));
    LocalMux I__6042 (
            .O(N__34708),
            .I(throttle_order_10));
    Odrv4 I__6041 (
            .O(N__34703),
            .I(throttle_order_10));
    InMux I__6040 (
            .O(N__34698),
            .I(N__34695));
    LocalMux I__6039 (
            .O(N__34695),
            .I(N__34688));
    InMux I__6038 (
            .O(N__34694),
            .I(N__34685));
    InMux I__6037 (
            .O(N__34693),
            .I(N__34680));
    InMux I__6036 (
            .O(N__34692),
            .I(N__34680));
    InMux I__6035 (
            .O(N__34691),
            .I(N__34674));
    Span4Mux_h I__6034 (
            .O(N__34688),
            .I(N__34667));
    LocalMux I__6033 (
            .O(N__34685),
            .I(N__34667));
    LocalMux I__6032 (
            .O(N__34680),
            .I(N__34667));
    InMux I__6031 (
            .O(N__34679),
            .I(N__34662));
    InMux I__6030 (
            .O(N__34678),
            .I(N__34662));
    InMux I__6029 (
            .O(N__34677),
            .I(N__34659));
    LocalMux I__6028 (
            .O(N__34674),
            .I(N__34656));
    Span4Mux_v I__6027 (
            .O(N__34667),
            .I(N__34649));
    LocalMux I__6026 (
            .O(N__34662),
            .I(N__34649));
    LocalMux I__6025 (
            .O(N__34659),
            .I(N__34649));
    Odrv4 I__6024 (
            .O(N__34656),
            .I(\dron_frame_decoder_1.N_218 ));
    Odrv4 I__6023 (
            .O(N__34649),
            .I(\dron_frame_decoder_1.N_218 ));
    InMux I__6022 (
            .O(N__34644),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    InMux I__6021 (
            .O(N__34641),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__6020 (
            .O(N__34638),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    InMux I__6019 (
            .O(N__34635),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__6018 (
            .O(N__34632),
            .I(N__34628));
    InMux I__6017 (
            .O(N__34631),
            .I(N__34625));
    LocalMux I__6016 (
            .O(N__34628),
            .I(N__34622));
    LocalMux I__6015 (
            .O(N__34625),
            .I(N__34619));
    Span4Mux_h I__6014 (
            .O(N__34622),
            .I(N__34616));
    Span4Mux_h I__6013 (
            .O(N__34619),
            .I(N__34613));
    Span4Mux_v I__6012 (
            .O(N__34616),
            .I(N__34610));
    Span4Mux_v I__6011 (
            .O(N__34613),
            .I(N__34607));
    Span4Mux_h I__6010 (
            .O(N__34610),
            .I(N__34604));
    Span4Mux_h I__6009 (
            .O(N__34607),
            .I(N__34601));
    Odrv4 I__6008 (
            .O(N__34604),
            .I(throttle_order_5));
    Odrv4 I__6007 (
            .O(N__34601),
            .I(throttle_order_5));
    InMux I__6006 (
            .O(N__34596),
            .I(N__34593));
    LocalMux I__6005 (
            .O(N__34593),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__6004 (
            .O(N__34590),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    InMux I__6003 (
            .O(N__34587),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__6002 (
            .O(N__34584),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__6001 (
            .O(N__34581),
            .I(N__34576));
    InMux I__6000 (
            .O(N__34580),
            .I(N__34571));
    InMux I__5999 (
            .O(N__34579),
            .I(N__34571));
    LocalMux I__5998 (
            .O(N__34576),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__5997 (
            .O(N__34571),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    InMux I__5996 (
            .O(N__34566),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__5995 (
            .O(N__34563),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    CascadeMux I__5994 (
            .O(N__34560),
            .I(N__34556));
    InMux I__5993 (
            .O(N__34559),
            .I(N__34552));
    InMux I__5992 (
            .O(N__34556),
            .I(N__34547));
    InMux I__5991 (
            .O(N__34555),
            .I(N__34547));
    LocalMux I__5990 (
            .O(N__34552),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__5989 (
            .O(N__34547),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    InMux I__5988 (
            .O(N__34542),
            .I(N__34538));
    InMux I__5987 (
            .O(N__34541),
            .I(N__34535));
    LocalMux I__5986 (
            .O(N__34538),
            .I(N__34532));
    LocalMux I__5985 (
            .O(N__34535),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    Odrv12 I__5984 (
            .O(N__34532),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    InMux I__5983 (
            .O(N__34527),
            .I(N__34523));
    InMux I__5982 (
            .O(N__34526),
            .I(N__34520));
    LocalMux I__5981 (
            .O(N__34523),
            .I(N__34517));
    LocalMux I__5980 (
            .O(N__34520),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    Odrv4 I__5979 (
            .O(N__34517),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    CascadeMux I__5978 (
            .O(N__34512),
            .I(N__34509));
    InMux I__5977 (
            .O(N__34509),
            .I(N__34505));
    InMux I__5976 (
            .O(N__34508),
            .I(N__34502));
    LocalMux I__5975 (
            .O(N__34505),
            .I(N__34499));
    LocalMux I__5974 (
            .O(N__34502),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    Odrv4 I__5973 (
            .O(N__34499),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__5972 (
            .O(N__34494),
            .I(N__34490));
    InMux I__5971 (
            .O(N__34493),
            .I(N__34487));
    LocalMux I__5970 (
            .O(N__34490),
            .I(N__34484));
    LocalMux I__5969 (
            .O(N__34487),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    Odrv4 I__5968 (
            .O(N__34484),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    InMux I__5967 (
            .O(N__34479),
            .I(N__34475));
    InMux I__5966 (
            .O(N__34478),
            .I(N__34472));
    LocalMux I__5965 (
            .O(N__34475),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    LocalMux I__5964 (
            .O(N__34472),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    CascadeMux I__5963 (
            .O(N__34467),
            .I(\dron_frame_decoder_1.WDT_RNIIVJ1Z0Z_4_cascade_ ));
    InMux I__5962 (
            .O(N__34464),
            .I(N__34458));
    InMux I__5961 (
            .O(N__34463),
            .I(N__34458));
    LocalMux I__5960 (
            .O(N__34458),
            .I(\dron_frame_decoder_1.WDT10lt14_0 ));
    InMux I__5959 (
            .O(N__34455),
            .I(N__34451));
    InMux I__5958 (
            .O(N__34454),
            .I(N__34448));
    LocalMux I__5957 (
            .O(N__34451),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__5956 (
            .O(N__34448),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    CascadeMux I__5955 (
            .O(N__34443),
            .I(N__34439));
    InMux I__5954 (
            .O(N__34442),
            .I(N__34436));
    InMux I__5953 (
            .O(N__34439),
            .I(N__34433));
    LocalMux I__5952 (
            .O(N__34436),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    LocalMux I__5951 (
            .O(N__34433),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    InMux I__5950 (
            .O(N__34428),
            .I(N__34425));
    LocalMux I__5949 (
            .O(N__34425),
            .I(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ));
    InMux I__5948 (
            .O(N__34422),
            .I(N__34417));
    InMux I__5947 (
            .O(N__34421),
            .I(N__34412));
    InMux I__5946 (
            .O(N__34420),
            .I(N__34412));
    LocalMux I__5945 (
            .O(N__34417),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__5944 (
            .O(N__34412),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__5943 (
            .O(N__34407),
            .I(N__34403));
    InMux I__5942 (
            .O(N__34406),
            .I(N__34400));
    LocalMux I__5941 (
            .O(N__34403),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    LocalMux I__5940 (
            .O(N__34400),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    CascadeMux I__5939 (
            .O(N__34395),
            .I(N__34390));
    InMux I__5938 (
            .O(N__34394),
            .I(N__34387));
    InMux I__5937 (
            .O(N__34393),
            .I(N__34382));
    InMux I__5936 (
            .O(N__34390),
            .I(N__34382));
    LocalMux I__5935 (
            .O(N__34387),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__5934 (
            .O(N__34382),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    InMux I__5933 (
            .O(N__34377),
            .I(N__34374));
    LocalMux I__5932 (
            .O(N__34374),
            .I(\dron_frame_decoder_1.WDT10lto13_1 ));
    CascadeMux I__5931 (
            .O(N__34371),
            .I(N__34367));
    CascadeMux I__5930 (
            .O(N__34370),
            .I(N__34363));
    InMux I__5929 (
            .O(N__34367),
            .I(N__34360));
    InMux I__5928 (
            .O(N__34366),
            .I(N__34357));
    InMux I__5927 (
            .O(N__34363),
            .I(N__34354));
    LocalMux I__5926 (
            .O(N__34360),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    LocalMux I__5925 (
            .O(N__34357),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    LocalMux I__5924 (
            .O(N__34354),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    InMux I__5923 (
            .O(N__34347),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__5922 (
            .O(N__34344),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    InMux I__5921 (
            .O(N__34341),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__5920 (
            .O(N__34338),
            .I(bfn_11_11_0_));
    InMux I__5919 (
            .O(N__34335),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    InMux I__5918 (
            .O(N__34332),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    InMux I__5917 (
            .O(N__34329),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    InMux I__5916 (
            .O(N__34326),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    InMux I__5915 (
            .O(N__34323),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__5914 (
            .O(N__34320),
            .I(N__34317));
    LocalMux I__5913 (
            .O(N__34317),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__5912 (
            .O(N__34314),
            .I(N__34310));
    InMux I__5911 (
            .O(N__34313),
            .I(N__34307));
    LocalMux I__5910 (
            .O(N__34310),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__5909 (
            .O(N__34307),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__5908 (
            .O(N__34302),
            .I(N__34298));
    InMux I__5907 (
            .O(N__34301),
            .I(N__34295));
    LocalMux I__5906 (
            .O(N__34298),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__5905 (
            .O(N__34295),
            .I(\reset_module_System.countZ0Z_11 ));
    CascadeMux I__5904 (
            .O(N__34290),
            .I(N__34287));
    InMux I__5903 (
            .O(N__34287),
            .I(N__34283));
    InMux I__5902 (
            .O(N__34286),
            .I(N__34280));
    LocalMux I__5901 (
            .O(N__34283),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__5900 (
            .O(N__34280),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__5899 (
            .O(N__34275),
            .I(N__34269));
    InMux I__5898 (
            .O(N__34274),
            .I(N__34269));
    LocalMux I__5897 (
            .O(N__34269),
            .I(\reset_module_System.countZ0Z_17 ));
    CascadeMux I__5896 (
            .O(N__34266),
            .I(N__34263));
    InMux I__5895 (
            .O(N__34263),
            .I(N__34254));
    InMux I__5894 (
            .O(N__34262),
            .I(N__34254));
    InMux I__5893 (
            .O(N__34261),
            .I(N__34254));
    LocalMux I__5892 (
            .O(N__34254),
            .I(N__34251));
    Span4Mux_h I__5891 (
            .O(N__34251),
            .I(N__34247));
    InMux I__5890 (
            .O(N__34250),
            .I(N__34244));
    Odrv4 I__5889 (
            .O(N__34247),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__5888 (
            .O(N__34244),
            .I(\reset_module_System.reset6_14 ));
    InMux I__5887 (
            .O(N__34239),
            .I(N__34233));
    InMux I__5886 (
            .O(N__34238),
            .I(N__34233));
    LocalMux I__5885 (
            .O(N__34233),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__5884 (
            .O(N__34230),
            .I(N__34226));
    InMux I__5883 (
            .O(N__34229),
            .I(N__34223));
    LocalMux I__5882 (
            .O(N__34226),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__5881 (
            .O(N__34223),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__5880 (
            .O(N__34218),
            .I(N__34214));
    InMux I__5879 (
            .O(N__34217),
            .I(N__34209));
    InMux I__5878 (
            .O(N__34214),
            .I(N__34209));
    LocalMux I__5877 (
            .O(N__34209),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__5876 (
            .O(N__34206),
            .I(N__34202));
    InMux I__5875 (
            .O(N__34205),
            .I(N__34199));
    LocalMux I__5874 (
            .O(N__34202),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__5873 (
            .O(N__34199),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__5872 (
            .O(N__34194),
            .I(N__34191));
    LocalMux I__5871 (
            .O(N__34191),
            .I(\reset_module_System.reset6_11 ));
    CascadeMux I__5870 (
            .O(N__34188),
            .I(N__34184));
    InMux I__5869 (
            .O(N__34187),
            .I(N__34181));
    InMux I__5868 (
            .O(N__34184),
            .I(N__34178));
    LocalMux I__5867 (
            .O(N__34181),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    LocalMux I__5866 (
            .O(N__34178),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__5865 (
            .O(N__34173),
            .I(N__34170));
    LocalMux I__5864 (
            .O(N__34170),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__5863 (
            .O(N__34167),
            .I(N__34164));
    LocalMux I__5862 (
            .O(N__34164),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__5861 (
            .O(N__34161),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    InMux I__5860 (
            .O(N__34158),
            .I(N__34155));
    LocalMux I__5859 (
            .O(N__34155),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__5858 (
            .O(N__34152),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    InMux I__5857 (
            .O(N__34149),
            .I(N__34146));
    LocalMux I__5856 (
            .O(N__34146),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__5855 (
            .O(N__34143),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    InMux I__5854 (
            .O(N__34140),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__5853 (
            .O(N__34137),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__5852 (
            .O(N__34134),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__5851 (
            .O(N__34131),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__5850 (
            .O(N__34128),
            .I(N__34124));
    InMux I__5849 (
            .O(N__34127),
            .I(N__34121));
    LocalMux I__5848 (
            .O(N__34124),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__5847 (
            .O(N__34121),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__5846 (
            .O(N__34116),
            .I(\reset_module_System.count_1_cry_15 ));
    InMux I__5845 (
            .O(N__34113),
            .I(bfn_11_9_0_));
    InMux I__5844 (
            .O(N__34110),
            .I(N__34106));
    InMux I__5843 (
            .O(N__34109),
            .I(N__34103));
    LocalMux I__5842 (
            .O(N__34106),
            .I(\reset_module_System.countZ0Z_18 ));
    LocalMux I__5841 (
            .O(N__34103),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__5840 (
            .O(N__34098),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__5839 (
            .O(N__34095),
            .I(\reset_module_System.count_1_cry_18 ));
    CascadeMux I__5838 (
            .O(N__34092),
            .I(N__34089));
    InMux I__5837 (
            .O(N__34089),
            .I(N__34085));
    InMux I__5836 (
            .O(N__34088),
            .I(N__34082));
    LocalMux I__5835 (
            .O(N__34085),
            .I(N__34079));
    LocalMux I__5834 (
            .O(N__34082),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__5833 (
            .O(N__34079),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__5832 (
            .O(N__34074),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__5831 (
            .O(N__34071),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__5830 (
            .O(N__34068),
            .I(N__34064));
    InMux I__5829 (
            .O(N__34067),
            .I(N__34061));
    LocalMux I__5828 (
            .O(N__34064),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__5827 (
            .O(N__34061),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__5826 (
            .O(N__34056),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__5825 (
            .O(N__34053),
            .I(N__34049));
    InMux I__5824 (
            .O(N__34052),
            .I(N__34046));
    LocalMux I__5823 (
            .O(N__34049),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__5822 (
            .O(N__34046),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__5821 (
            .O(N__34041),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__5820 (
            .O(N__34038),
            .I(N__34034));
    InMux I__5819 (
            .O(N__34037),
            .I(N__34031));
    LocalMux I__5818 (
            .O(N__34034),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__5817 (
            .O(N__34031),
            .I(\reset_module_System.countZ0Z_7 ));
    InMux I__5816 (
            .O(N__34026),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__5815 (
            .O(N__34023),
            .I(N__34019));
    InMux I__5814 (
            .O(N__34022),
            .I(N__34016));
    LocalMux I__5813 (
            .O(N__34019),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__5812 (
            .O(N__34016),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__5811 (
            .O(N__34011),
            .I(\reset_module_System.count_1_cry_7 ));
    CascadeMux I__5810 (
            .O(N__34008),
            .I(N__34004));
    InMux I__5809 (
            .O(N__34007),
            .I(N__34001));
    InMux I__5808 (
            .O(N__34004),
            .I(N__33998));
    LocalMux I__5807 (
            .O(N__34001),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__5806 (
            .O(N__33998),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__5805 (
            .O(N__33993),
            .I(bfn_11_8_0_));
    InMux I__5804 (
            .O(N__33990),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__5803 (
            .O(N__33987),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__5802 (
            .O(N__33984),
            .I(N__33980));
    InMux I__5801 (
            .O(N__33983),
            .I(N__33977));
    LocalMux I__5800 (
            .O(N__33980),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__5799 (
            .O(N__33977),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__5798 (
            .O(N__33972),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__5797 (
            .O(N__33969),
            .I(N__33965));
    InMux I__5796 (
            .O(N__33968),
            .I(N__33962));
    LocalMux I__5795 (
            .O(N__33965),
            .I(N__33959));
    LocalMux I__5794 (
            .O(N__33962),
            .I(N__33954));
    Span4Mux_v I__5793 (
            .O(N__33959),
            .I(N__33954));
    Span4Mux_h I__5792 (
            .O(N__33954),
            .I(N__33951));
    Span4Mux_v I__5791 (
            .O(N__33951),
            .I(N__33948));
    Odrv4 I__5790 (
            .O(N__33948),
            .I(\pid_front.error_p_regZ0Z_11 ));
    InMux I__5789 (
            .O(N__33945),
            .I(N__33939));
    InMux I__5788 (
            .O(N__33944),
            .I(N__33939));
    LocalMux I__5787 (
            .O(N__33939),
            .I(\uart_drone.un1_state_7_0 ));
    InMux I__5786 (
            .O(N__33936),
            .I(N__33933));
    LocalMux I__5785 (
            .O(N__33933),
            .I(\uart_drone.CO0 ));
    InMux I__5784 (
            .O(N__33930),
            .I(N__33923));
    InMux I__5783 (
            .O(N__33929),
            .I(N__33923));
    InMux I__5782 (
            .O(N__33928),
            .I(N__33920));
    LocalMux I__5781 (
            .O(N__33923),
            .I(N__33913));
    LocalMux I__5780 (
            .O(N__33920),
            .I(N__33913));
    CascadeMux I__5779 (
            .O(N__33919),
            .I(N__33907));
    InMux I__5778 (
            .O(N__33918),
            .I(N__33904));
    Span4Mux_h I__5777 (
            .O(N__33913),
            .I(N__33901));
    InMux I__5776 (
            .O(N__33912),
            .I(N__33898));
    InMux I__5775 (
            .O(N__33911),
            .I(N__33891));
    InMux I__5774 (
            .O(N__33910),
            .I(N__33891));
    InMux I__5773 (
            .O(N__33907),
            .I(N__33891));
    LocalMux I__5772 (
            .O(N__33904),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__5771 (
            .O(N__33901),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__5770 (
            .O(N__33898),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__5769 (
            .O(N__33891),
            .I(\uart_drone.stateZ0Z_3 ));
    CascadeMux I__5768 (
            .O(N__33882),
            .I(N__33878));
    CascadeMux I__5767 (
            .O(N__33881),
            .I(N__33875));
    InMux I__5766 (
            .O(N__33878),
            .I(N__33869));
    InMux I__5765 (
            .O(N__33875),
            .I(N__33869));
    InMux I__5764 (
            .O(N__33874),
            .I(N__33866));
    LocalMux I__5763 (
            .O(N__33869),
            .I(\uart_drone.un1_state_4_0 ));
    LocalMux I__5762 (
            .O(N__33866),
            .I(\uart_drone.un1_state_4_0 ));
    CascadeMux I__5761 (
            .O(N__33861),
            .I(N__33856));
    InMux I__5760 (
            .O(N__33860),
            .I(N__33853));
    InMux I__5759 (
            .O(N__33859),
            .I(N__33848));
    InMux I__5758 (
            .O(N__33856),
            .I(N__33845));
    LocalMux I__5757 (
            .O(N__33853),
            .I(N__33842));
    InMux I__5756 (
            .O(N__33852),
            .I(N__33837));
    InMux I__5755 (
            .O(N__33851),
            .I(N__33837));
    LocalMux I__5754 (
            .O(N__33848),
            .I(N__33831));
    LocalMux I__5753 (
            .O(N__33845),
            .I(N__33831));
    Span4Mux_v I__5752 (
            .O(N__33842),
            .I(N__33826));
    LocalMux I__5751 (
            .O(N__33837),
            .I(N__33826));
    CascadeMux I__5750 (
            .O(N__33836),
            .I(N__33822));
    Span4Mux_h I__5749 (
            .O(N__33831),
            .I(N__33818));
    Span4Mux_h I__5748 (
            .O(N__33826),
            .I(N__33815));
    InMux I__5747 (
            .O(N__33825),
            .I(N__33812));
    InMux I__5746 (
            .O(N__33822),
            .I(N__33807));
    InMux I__5745 (
            .O(N__33821),
            .I(N__33807));
    Odrv4 I__5744 (
            .O(N__33818),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__5743 (
            .O(N__33815),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__5742 (
            .O(N__33812),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__5741 (
            .O(N__33807),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__5740 (
            .O(N__33798),
            .I(N__33794));
    CascadeMux I__5739 (
            .O(N__33797),
            .I(N__33791));
    LocalMux I__5738 (
            .O(N__33794),
            .I(N__33782));
    InMux I__5737 (
            .O(N__33791),
            .I(N__33777));
    InMux I__5736 (
            .O(N__33790),
            .I(N__33777));
    CascadeMux I__5735 (
            .O(N__33789),
            .I(N__33773));
    InMux I__5734 (
            .O(N__33788),
            .I(N__33770));
    InMux I__5733 (
            .O(N__33787),
            .I(N__33763));
    InMux I__5732 (
            .O(N__33786),
            .I(N__33763));
    InMux I__5731 (
            .O(N__33785),
            .I(N__33763));
    Span4Mux_h I__5730 (
            .O(N__33782),
            .I(N__33760));
    LocalMux I__5729 (
            .O(N__33777),
            .I(N__33757));
    InMux I__5728 (
            .O(N__33776),
            .I(N__33752));
    InMux I__5727 (
            .O(N__33773),
            .I(N__33752));
    LocalMux I__5726 (
            .O(N__33770),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__5725 (
            .O(N__33763),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__5724 (
            .O(N__33760),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__5723 (
            .O(N__33757),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__5722 (
            .O(N__33752),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    InMux I__5721 (
            .O(N__33741),
            .I(N__33738));
    LocalMux I__5720 (
            .O(N__33738),
            .I(N__33735));
    Span4Mux_h I__5719 (
            .O(N__33735),
            .I(N__33731));
    InMux I__5718 (
            .O(N__33734),
            .I(N__33728));
    Odrv4 I__5717 (
            .O(N__33731),
            .I(\uart_drone.N_144_1 ));
    LocalMux I__5716 (
            .O(N__33728),
            .I(\uart_drone.N_144_1 ));
    InMux I__5715 (
            .O(N__33723),
            .I(N__33718));
    InMux I__5714 (
            .O(N__33722),
            .I(N__33715));
    InMux I__5713 (
            .O(N__33721),
            .I(N__33712));
    LocalMux I__5712 (
            .O(N__33718),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__5711 (
            .O(N__33715),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__5710 (
            .O(N__33712),
            .I(\reset_module_System.countZ0Z_1 ));
    CascadeMux I__5709 (
            .O(N__33705),
            .I(N__33699));
    InMux I__5708 (
            .O(N__33704),
            .I(N__33694));
    InMux I__5707 (
            .O(N__33703),
            .I(N__33694));
    InMux I__5706 (
            .O(N__33702),
            .I(N__33691));
    InMux I__5705 (
            .O(N__33699),
            .I(N__33688));
    LocalMux I__5704 (
            .O(N__33694),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__5703 (
            .O(N__33691),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__5702 (
            .O(N__33688),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__5701 (
            .O(N__33681),
            .I(N__33677));
    InMux I__5700 (
            .O(N__33680),
            .I(N__33674));
    LocalMux I__5699 (
            .O(N__33677),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__5698 (
            .O(N__33674),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__5697 (
            .O(N__33669),
            .I(N__33666));
    LocalMux I__5696 (
            .O(N__33666),
            .I(\reset_module_System.count_1_2 ));
    InMux I__5695 (
            .O(N__33663),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__5694 (
            .O(N__33660),
            .I(N__33656));
    InMux I__5693 (
            .O(N__33659),
            .I(N__33653));
    LocalMux I__5692 (
            .O(N__33656),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__5691 (
            .O(N__33653),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__5690 (
            .O(N__33648),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__5689 (
            .O(N__33645),
            .I(N__33641));
    InMux I__5688 (
            .O(N__33644),
            .I(N__33638));
    LocalMux I__5687 (
            .O(N__33641),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__5686 (
            .O(N__33638),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__5685 (
            .O(N__33633),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__5684 (
            .O(N__33630),
            .I(N__33627));
    LocalMux I__5683 (
            .O(N__33627),
            .I(N__33624));
    Odrv4 I__5682 (
            .O(N__33624),
            .I(\pid_front.pid_prereg_esr_RNI6FQ75Z0Z_23 ));
    InMux I__5681 (
            .O(N__33621),
            .I(N__33617));
    InMux I__5680 (
            .O(N__33620),
            .I(N__33614));
    LocalMux I__5679 (
            .O(N__33617),
            .I(\pid_front.un1_pid_prereg_42 ));
    LocalMux I__5678 (
            .O(N__33614),
            .I(\pid_front.un1_pid_prereg_42 ));
    InMux I__5677 (
            .O(N__33609),
            .I(N__33606));
    LocalMux I__5676 (
            .O(N__33606),
            .I(N__33601));
    InMux I__5675 (
            .O(N__33605),
            .I(N__33596));
    InMux I__5674 (
            .O(N__33604),
            .I(N__33596));
    Span4Mux_v I__5673 (
            .O(N__33601),
            .I(N__33593));
    LocalMux I__5672 (
            .O(N__33596),
            .I(N__33590));
    Odrv4 I__5671 (
            .O(N__33593),
            .I(\pid_front.un1_pid_prereg_47 ));
    Odrv4 I__5670 (
            .O(N__33590),
            .I(\pid_front.un1_pid_prereg_47 ));
    CascadeMux I__5669 (
            .O(N__33585),
            .I(\pid_front.un1_pid_prereg_42_cascade_ ));
    InMux I__5668 (
            .O(N__33582),
            .I(N__33578));
    InMux I__5667 (
            .O(N__33581),
            .I(N__33575));
    LocalMux I__5666 (
            .O(N__33578),
            .I(N__33570));
    LocalMux I__5665 (
            .O(N__33575),
            .I(N__33570));
    Span4Mux_v I__5664 (
            .O(N__33570),
            .I(N__33567));
    Span4Mux_h I__5663 (
            .O(N__33567),
            .I(N__33564));
    Span4Mux_h I__5662 (
            .O(N__33564),
            .I(N__33561));
    Odrv4 I__5661 (
            .O(N__33561),
            .I(\pid_front.error_p_regZ0Z_16 ));
    InMux I__5660 (
            .O(N__33558),
            .I(N__33555));
    LocalMux I__5659 (
            .O(N__33555),
            .I(N__33551));
    InMux I__5658 (
            .O(N__33554),
            .I(N__33548));
    Span4Mux_v I__5657 (
            .O(N__33551),
            .I(N__33543));
    LocalMux I__5656 (
            .O(N__33548),
            .I(N__33543));
    Span4Mux_v I__5655 (
            .O(N__33543),
            .I(N__33540));
    Odrv4 I__5654 (
            .O(N__33540),
            .I(\pid_front.error_d_reg_prevZ0Z_16 ));
    InMux I__5653 (
            .O(N__33537),
            .I(N__33530));
    InMux I__5652 (
            .O(N__33536),
            .I(N__33530));
    InMux I__5651 (
            .O(N__33535),
            .I(N__33527));
    LocalMux I__5650 (
            .O(N__33530),
            .I(N__33524));
    LocalMux I__5649 (
            .O(N__33527),
            .I(N__33519));
    Span4Mux_h I__5648 (
            .O(N__33524),
            .I(N__33519));
    Odrv4 I__5647 (
            .O(N__33519),
            .I(\pid_front.un1_pid_prereg_35 ));
    CascadeMux I__5646 (
            .O(N__33516),
            .I(\pid_front.un1_pid_prereg_36_cascade_ ));
    InMux I__5645 (
            .O(N__33513),
            .I(N__33510));
    LocalMux I__5644 (
            .O(N__33510),
            .I(N__33506));
    InMux I__5643 (
            .O(N__33509),
            .I(N__33503));
    Odrv4 I__5642 (
            .O(N__33506),
            .I(\pid_front.un1_pid_prereg_30 ));
    LocalMux I__5641 (
            .O(N__33503),
            .I(\pid_front.un1_pid_prereg_30 ));
    InMux I__5640 (
            .O(N__33498),
            .I(N__33492));
    InMux I__5639 (
            .O(N__33497),
            .I(N__33492));
    LocalMux I__5638 (
            .O(N__33492),
            .I(N__33489));
    Span4Mux_v I__5637 (
            .O(N__33489),
            .I(N__33486));
    Sp12to4 I__5636 (
            .O(N__33486),
            .I(N__33483));
    Span12Mux_h I__5635 (
            .O(N__33483),
            .I(N__33480));
    Odrv12 I__5634 (
            .O(N__33480),
            .I(\pid_front.error_p_regZ0Z_17 ));
    CascadeMux I__5633 (
            .O(N__33477),
            .I(N__33474));
    InMux I__5632 (
            .O(N__33474),
            .I(N__33468));
    InMux I__5631 (
            .O(N__33473),
            .I(N__33468));
    LocalMux I__5630 (
            .O(N__33468),
            .I(\pid_front.error_d_reg_prevZ0Z_17 ));
    InMux I__5629 (
            .O(N__33465),
            .I(N__33459));
    InMux I__5628 (
            .O(N__33464),
            .I(N__33459));
    LocalMux I__5627 (
            .O(N__33459),
            .I(\pid_front.un1_pid_prereg_41 ));
    CascadeMux I__5626 (
            .O(N__33456),
            .I(\pid_front.un1_pid_prereg_41_cascade_ ));
    InMux I__5625 (
            .O(N__33453),
            .I(N__33449));
    InMux I__5624 (
            .O(N__33452),
            .I(N__33446));
    LocalMux I__5623 (
            .O(N__33449),
            .I(\pid_front.un1_pid_prereg_36 ));
    LocalMux I__5622 (
            .O(N__33446),
            .I(\pid_front.un1_pid_prereg_36 ));
    InMux I__5621 (
            .O(N__33441),
            .I(N__33438));
    LocalMux I__5620 (
            .O(N__33438),
            .I(\pid_front.un1_reset_0_i_sn ));
    CascadeMux I__5619 (
            .O(N__33435),
            .I(N__33432));
    InMux I__5618 (
            .O(N__33432),
            .I(N__33429));
    LocalMux I__5617 (
            .O(N__33429),
            .I(N__33425));
    CascadeMux I__5616 (
            .O(N__33428),
            .I(N__33421));
    Span12Mux_v I__5615 (
            .O(N__33425),
            .I(N__33417));
    InMux I__5614 (
            .O(N__33424),
            .I(N__33412));
    InMux I__5613 (
            .O(N__33421),
            .I(N__33412));
    InMux I__5612 (
            .O(N__33420),
            .I(N__33409));
    Odrv12 I__5611 (
            .O(N__33417),
            .I(\pid_alt.error_i_acumm7lto5 ));
    LocalMux I__5610 (
            .O(N__33412),
            .I(\pid_alt.error_i_acumm7lto5 ));
    LocalMux I__5609 (
            .O(N__33409),
            .I(\pid_alt.error_i_acumm7lto5 ));
    InMux I__5608 (
            .O(N__33402),
            .I(N__33399));
    LocalMux I__5607 (
            .O(N__33399),
            .I(N__33396));
    Span4Mux_h I__5606 (
            .O(N__33396),
            .I(N__33393));
    Span4Mux_h I__5605 (
            .O(N__33393),
            .I(N__33390));
    Span4Mux_v I__5604 (
            .O(N__33390),
            .I(N__33382));
    InMux I__5603 (
            .O(N__33389),
            .I(N__33371));
    InMux I__5602 (
            .O(N__33388),
            .I(N__33371));
    InMux I__5601 (
            .O(N__33387),
            .I(N__33371));
    InMux I__5600 (
            .O(N__33386),
            .I(N__33371));
    InMux I__5599 (
            .O(N__33385),
            .I(N__33371));
    Odrv4 I__5598 (
            .O(N__33382),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__5597 (
            .O(N__33371),
            .I(\pid_alt.N_62_mux ));
    InMux I__5596 (
            .O(N__33366),
            .I(N__33363));
    LocalMux I__5595 (
            .O(N__33363),
            .I(N__33360));
    Span4Mux_h I__5594 (
            .O(N__33360),
            .I(N__33357));
    Span4Mux_v I__5593 (
            .O(N__33357),
            .I(N__33353));
    InMux I__5592 (
            .O(N__33356),
            .I(N__33350));
    Span4Mux_h I__5591 (
            .O(N__33353),
            .I(N__33347));
    LocalMux I__5590 (
            .O(N__33350),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    Odrv4 I__5589 (
            .O(N__33347),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    SRMux I__5588 (
            .O(N__33342),
            .I(N__33339));
    LocalMux I__5587 (
            .O(N__33339),
            .I(N__33335));
    SRMux I__5586 (
            .O(N__33338),
            .I(N__33332));
    Span4Mux_v I__5585 (
            .O(N__33335),
            .I(N__33327));
    LocalMux I__5584 (
            .O(N__33332),
            .I(N__33324));
    SRMux I__5583 (
            .O(N__33331),
            .I(N__33321));
    SRMux I__5582 (
            .O(N__33330),
            .I(N__33318));
    Span4Mux_h I__5581 (
            .O(N__33327),
            .I(N__33315));
    Span4Mux_h I__5580 (
            .O(N__33324),
            .I(N__33310));
    LocalMux I__5579 (
            .O(N__33321),
            .I(N__33310));
    LocalMux I__5578 (
            .O(N__33318),
            .I(N__33307));
    Odrv4 I__5577 (
            .O(N__33315),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__5576 (
            .O(N__33310),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__5575 (
            .O(N__33307),
            .I(\pid_alt.un1_reset_1_0_i ));
    CascadeMux I__5574 (
            .O(N__33300),
            .I(N__33297));
    InMux I__5573 (
            .O(N__33297),
            .I(N__33294));
    LocalMux I__5572 (
            .O(N__33294),
            .I(N__33290));
    InMux I__5571 (
            .O(N__33293),
            .I(N__33287));
    Span4Mux_h I__5570 (
            .O(N__33290),
            .I(N__33284));
    LocalMux I__5569 (
            .O(N__33287),
            .I(N__33281));
    Odrv4 I__5568 (
            .O(N__33284),
            .I(\pid_front.un1_pid_prereg_57 ));
    Odrv4 I__5567 (
            .O(N__33281),
            .I(\pid_front.un1_pid_prereg_57 ));
    InMux I__5566 (
            .O(N__33276),
            .I(N__33273));
    LocalMux I__5565 (
            .O(N__33273),
            .I(N__33269));
    InMux I__5564 (
            .O(N__33272),
            .I(N__33266));
    Span4Mux_v I__5563 (
            .O(N__33269),
            .I(N__33263));
    LocalMux I__5562 (
            .O(N__33266),
            .I(N__33260));
    Span4Mux_v I__5561 (
            .O(N__33263),
            .I(N__33257));
    Sp12to4 I__5560 (
            .O(N__33260),
            .I(N__33254));
    Sp12to4 I__5559 (
            .O(N__33257),
            .I(N__33249));
    Span12Mux_v I__5558 (
            .O(N__33254),
            .I(N__33249));
    Odrv12 I__5557 (
            .O(N__33249),
            .I(\pid_front.error_p_regZ0Z_18 ));
    CascadeMux I__5556 (
            .O(N__33246),
            .I(N__33242));
    InMux I__5555 (
            .O(N__33245),
            .I(N__33238));
    InMux I__5554 (
            .O(N__33242),
            .I(N__33233));
    InMux I__5553 (
            .O(N__33241),
            .I(N__33233));
    LocalMux I__5552 (
            .O(N__33238),
            .I(N__33230));
    LocalMux I__5551 (
            .O(N__33233),
            .I(N__33227));
    Span4Mux_h I__5550 (
            .O(N__33230),
            .I(N__33224));
    Odrv4 I__5549 (
            .O(N__33227),
            .I(\pid_front.un1_pid_prereg_18 ));
    Odrv4 I__5548 (
            .O(N__33224),
            .I(\pid_front.un1_pid_prereg_18 ));
    InMux I__5547 (
            .O(N__33219),
            .I(N__33213));
    InMux I__5546 (
            .O(N__33218),
            .I(N__33213));
    LocalMux I__5545 (
            .O(N__33213),
            .I(N__33210));
    Span4Mux_v I__5544 (
            .O(N__33210),
            .I(N__33207));
    Span4Mux_v I__5543 (
            .O(N__33207),
            .I(N__33204));
    Sp12to4 I__5542 (
            .O(N__33204),
            .I(N__33201));
    Odrv12 I__5541 (
            .O(N__33201),
            .I(\pid_front.error_p_regZ0Z_13 ));
    InMux I__5540 (
            .O(N__33198),
            .I(N__33192));
    InMux I__5539 (
            .O(N__33197),
            .I(N__33192));
    LocalMux I__5538 (
            .O(N__33192),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    InMux I__5537 (
            .O(N__33189),
            .I(N__33183));
    InMux I__5536 (
            .O(N__33188),
            .I(N__33183));
    LocalMux I__5535 (
            .O(N__33183),
            .I(N__33179));
    InMux I__5534 (
            .O(N__33182),
            .I(N__33176));
    Odrv4 I__5533 (
            .O(N__33179),
            .I(\pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ));
    LocalMux I__5532 (
            .O(N__33176),
            .I(\pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ));
    CascadeMux I__5531 (
            .O(N__33171),
            .I(\pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13_cascade_ ));
    CascadeMux I__5530 (
            .O(N__33168),
            .I(\pid_front.pid_prereg_esr_RNICUKFAZ0Z_6_cascade_ ));
    CascadeMux I__5529 (
            .O(N__33165),
            .I(\pid_front.un1_reset_0_i_cascade_ ));
    InMux I__5528 (
            .O(N__33162),
            .I(N__33159));
    LocalMux I__5527 (
            .O(N__33159),
            .I(\pid_front.un1_reset_0_i_rn_0 ));
    CascadeMux I__5526 (
            .O(N__33156),
            .I(\pid_front.m32_1_cascade_ ));
    InMux I__5525 (
            .O(N__33153),
            .I(N__33150));
    LocalMux I__5524 (
            .O(N__33150),
            .I(N__33147));
    Odrv12 I__5523 (
            .O(N__33147),
            .I(\pid_front.O_0_5 ));
    InMux I__5522 (
            .O(N__33144),
            .I(N__33138));
    InMux I__5521 (
            .O(N__33143),
            .I(N__33138));
    LocalMux I__5520 (
            .O(N__33138),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ));
    CascadeMux I__5519 (
            .O(N__33135),
            .I(N__33132));
    InMux I__5518 (
            .O(N__33132),
            .I(N__33120));
    InMux I__5517 (
            .O(N__33131),
            .I(N__33120));
    InMux I__5516 (
            .O(N__33130),
            .I(N__33120));
    InMux I__5515 (
            .O(N__33129),
            .I(N__33120));
    LocalMux I__5514 (
            .O(N__33120),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    CascadeMux I__5513 (
            .O(N__33117),
            .I(N__33113));
    CascadeMux I__5512 (
            .O(N__33116),
            .I(N__33110));
    InMux I__5511 (
            .O(N__33113),
            .I(N__33102));
    InMux I__5510 (
            .O(N__33110),
            .I(N__33102));
    InMux I__5509 (
            .O(N__33109),
            .I(N__33099));
    InMux I__5508 (
            .O(N__33108),
            .I(N__33094));
    InMux I__5507 (
            .O(N__33107),
            .I(N__33094));
    LocalMux I__5506 (
            .O(N__33102),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__5505 (
            .O(N__33099),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__5504 (
            .O(N__33094),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    InMux I__5503 (
            .O(N__33087),
            .I(N__33084));
    LocalMux I__5502 (
            .O(N__33084),
            .I(\dron_frame_decoder_1.drone_H_disp_side_10 ));
    CEMux I__5501 (
            .O(N__33081),
            .I(N__33078));
    LocalMux I__5500 (
            .O(N__33078),
            .I(N__33074));
    CEMux I__5499 (
            .O(N__33077),
            .I(N__33071));
    Span4Mux_v I__5498 (
            .O(N__33074),
            .I(N__33068));
    LocalMux I__5497 (
            .O(N__33071),
            .I(N__33065));
    Odrv4 I__5496 (
            .O(N__33068),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    Odrv4 I__5495 (
            .O(N__33065),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    InMux I__5494 (
            .O(N__33060),
            .I(N__33057));
    LocalMux I__5493 (
            .O(N__33057),
            .I(N__33054));
    Odrv4 I__5492 (
            .O(N__33054),
            .I(\dron_frame_decoder_1.N_219_4 ));
    CascadeMux I__5491 (
            .O(N__33051),
            .I(\dron_frame_decoder_1.N_219_4_cascade_ ));
    InMux I__5490 (
            .O(N__33048),
            .I(N__33045));
    LocalMux I__5489 (
            .O(N__33045),
            .I(N__33042));
    Odrv4 I__5488 (
            .O(N__33042),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_1_3 ));
    InMux I__5487 (
            .O(N__33039),
            .I(N__33036));
    LocalMux I__5486 (
            .O(N__33036),
            .I(N__33033));
    Span4Mux_v I__5485 (
            .O(N__33033),
            .I(N__33030));
    Odrv4 I__5484 (
            .O(N__33030),
            .I(scaler_4_data_5));
    CascadeMux I__5483 (
            .O(N__33027),
            .I(N__33023));
    InMux I__5482 (
            .O(N__33026),
            .I(N__33020));
    InMux I__5481 (
            .O(N__33023),
            .I(N__33017));
    LocalMux I__5480 (
            .O(N__33020),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__5479 (
            .O(N__33017),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    CascadeMux I__5478 (
            .O(N__33012),
            .I(N__33008));
    InMux I__5477 (
            .O(N__33011),
            .I(N__33005));
    InMux I__5476 (
            .O(N__33008),
            .I(N__33002));
    LocalMux I__5475 (
            .O(N__33005),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__5474 (
            .O(N__33002),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    CEMux I__5473 (
            .O(N__32997),
            .I(N__32993));
    CEMux I__5472 (
            .O(N__32996),
            .I(N__32990));
    LocalMux I__5471 (
            .O(N__32993),
            .I(\uart_drone.data_rdyc_1_0 ));
    LocalMux I__5470 (
            .O(N__32990),
            .I(\uart_drone.data_rdyc_1_0 ));
    SRMux I__5469 (
            .O(N__32985),
            .I(N__32982));
    LocalMux I__5468 (
            .O(N__32982),
            .I(N__32978));
    SRMux I__5467 (
            .O(N__32981),
            .I(N__32975));
    Span4Mux_h I__5466 (
            .O(N__32978),
            .I(N__32972));
    LocalMux I__5465 (
            .O(N__32975),
            .I(N__32969));
    Odrv4 I__5464 (
            .O(N__32972),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    Odrv4 I__5463 (
            .O(N__32969),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    InMux I__5462 (
            .O(N__32964),
            .I(N__32961));
    LocalMux I__5461 (
            .O(N__32961),
            .I(N__32958));
    Odrv12 I__5460 (
            .O(N__32958),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__5459 (
            .O(N__32955),
            .I(N__32952));
    LocalMux I__5458 (
            .O(N__32952),
            .I(\dron_frame_decoder_1.N_263_5 ));
    CascadeMux I__5457 (
            .O(N__32949),
            .I(\dron_frame_decoder_1.N_263_5_cascade_ ));
    InMux I__5456 (
            .O(N__32946),
            .I(N__32942));
    InMux I__5455 (
            .O(N__32945),
            .I(N__32938));
    LocalMux I__5454 (
            .O(N__32942),
            .I(N__32935));
    InMux I__5453 (
            .O(N__32941),
            .I(N__32932));
    LocalMux I__5452 (
            .O(N__32938),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    Odrv4 I__5451 (
            .O(N__32935),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    LocalMux I__5450 (
            .O(N__32932),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    InMux I__5449 (
            .O(N__32925),
            .I(N__32922));
    LocalMux I__5448 (
            .O(N__32922),
            .I(N__32919));
    Span4Mux_h I__5447 (
            .O(N__32919),
            .I(N__32916));
    Odrv4 I__5446 (
            .O(N__32916),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__5445 (
            .O(N__32913),
            .I(N__32910));
    LocalMux I__5444 (
            .O(N__32910),
            .I(N__32907));
    Odrv4 I__5443 (
            .O(N__32907),
            .I(\uart_drone.data_Auxce_0_6 ));
    IoInMux I__5442 (
            .O(N__32904),
            .I(N__32901));
    LocalMux I__5441 (
            .O(N__32901),
            .I(N__32898));
    IoSpan4Mux I__5440 (
            .O(N__32898),
            .I(N__32885));
    InMux I__5439 (
            .O(N__32897),
            .I(N__32882));
    InMux I__5438 (
            .O(N__32896),
            .I(N__32865));
    InMux I__5437 (
            .O(N__32895),
            .I(N__32865));
    InMux I__5436 (
            .O(N__32894),
            .I(N__32865));
    InMux I__5435 (
            .O(N__32893),
            .I(N__32865));
    InMux I__5434 (
            .O(N__32892),
            .I(N__32865));
    InMux I__5433 (
            .O(N__32891),
            .I(N__32865));
    InMux I__5432 (
            .O(N__32890),
            .I(N__32865));
    InMux I__5431 (
            .O(N__32889),
            .I(N__32865));
    CascadeMux I__5430 (
            .O(N__32888),
            .I(N__32861));
    IoSpan4Mux I__5429 (
            .O(N__32885),
            .I(N__32856));
    LocalMux I__5428 (
            .O(N__32882),
            .I(N__32851));
    LocalMux I__5427 (
            .O(N__32865),
            .I(N__32851));
    InMux I__5426 (
            .O(N__32864),
            .I(N__32848));
    InMux I__5425 (
            .O(N__32861),
            .I(N__32843));
    InMux I__5424 (
            .O(N__32860),
            .I(N__32843));
    InMux I__5423 (
            .O(N__32859),
            .I(N__32840));
    Span4Mux_s2_v I__5422 (
            .O(N__32856),
            .I(N__32835));
    Span4Mux_v I__5421 (
            .O(N__32851),
            .I(N__32835));
    LocalMux I__5420 (
            .O(N__32848),
            .I(N__32832));
    LocalMux I__5419 (
            .O(N__32843),
            .I(debug_CH0_16A_c));
    LocalMux I__5418 (
            .O(N__32840),
            .I(debug_CH0_16A_c));
    Odrv4 I__5417 (
            .O(N__32835),
            .I(debug_CH0_16A_c));
    Odrv12 I__5416 (
            .O(N__32832),
            .I(debug_CH0_16A_c));
    InMux I__5415 (
            .O(N__32823),
            .I(N__32807));
    InMux I__5414 (
            .O(N__32822),
            .I(N__32807));
    InMux I__5413 (
            .O(N__32821),
            .I(N__32807));
    InMux I__5412 (
            .O(N__32820),
            .I(N__32807));
    InMux I__5411 (
            .O(N__32819),
            .I(N__32798));
    InMux I__5410 (
            .O(N__32818),
            .I(N__32798));
    InMux I__5409 (
            .O(N__32817),
            .I(N__32798));
    InMux I__5408 (
            .O(N__32816),
            .I(N__32798));
    LocalMux I__5407 (
            .O(N__32807),
            .I(N__32793));
    LocalMux I__5406 (
            .O(N__32798),
            .I(N__32793));
    Odrv4 I__5405 (
            .O(N__32793),
            .I(\uart_drone.un1_state_2_0 ));
    SRMux I__5404 (
            .O(N__32790),
            .I(N__32787));
    LocalMux I__5403 (
            .O(N__32787),
            .I(N__32784));
    Span4Mux_h I__5402 (
            .O(N__32784),
            .I(N__32781));
    Odrv4 I__5401 (
            .O(N__32781),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    CascadeMux I__5400 (
            .O(N__32778),
            .I(N__32774));
    InMux I__5399 (
            .O(N__32777),
            .I(N__32771));
    InMux I__5398 (
            .O(N__32774),
            .I(N__32768));
    LocalMux I__5397 (
            .O(N__32771),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__5396 (
            .O(N__32768),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    CascadeMux I__5395 (
            .O(N__32763),
            .I(N__32759));
    InMux I__5394 (
            .O(N__32762),
            .I(N__32756));
    InMux I__5393 (
            .O(N__32759),
            .I(N__32753));
    LocalMux I__5392 (
            .O(N__32756),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__5391 (
            .O(N__32753),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    CascadeMux I__5390 (
            .O(N__32748),
            .I(N__32744));
    InMux I__5389 (
            .O(N__32747),
            .I(N__32741));
    InMux I__5388 (
            .O(N__32744),
            .I(N__32738));
    LocalMux I__5387 (
            .O(N__32741),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__5386 (
            .O(N__32738),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    CascadeMux I__5385 (
            .O(N__32733),
            .I(N__32729));
    InMux I__5384 (
            .O(N__32732),
            .I(N__32726));
    InMux I__5383 (
            .O(N__32729),
            .I(N__32723));
    LocalMux I__5382 (
            .O(N__32726),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__5381 (
            .O(N__32723),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    CascadeMux I__5380 (
            .O(N__32718),
            .I(N__32715));
    InMux I__5379 (
            .O(N__32715),
            .I(N__32711));
    InMux I__5378 (
            .O(N__32714),
            .I(N__32708));
    LocalMux I__5377 (
            .O(N__32711),
            .I(N__32705));
    LocalMux I__5376 (
            .O(N__32708),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    Odrv4 I__5375 (
            .O(N__32705),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    CascadeMux I__5374 (
            .O(N__32700),
            .I(\reset_module_System.reset6_3_cascade_ ));
    InMux I__5373 (
            .O(N__32697),
            .I(N__32694));
    LocalMux I__5372 (
            .O(N__32694),
            .I(\reset_module_System.reset6_13 ));
    CascadeMux I__5371 (
            .O(N__32691),
            .I(\reset_module_System.reset6_17_cascade_ ));
    InMux I__5370 (
            .O(N__32688),
            .I(N__32679));
    InMux I__5369 (
            .O(N__32687),
            .I(N__32679));
    InMux I__5368 (
            .O(N__32686),
            .I(N__32679));
    LocalMux I__5367 (
            .O(N__32679),
            .I(\reset_module_System.reset6_19 ));
    InMux I__5366 (
            .O(N__32676),
            .I(N__32669));
    InMux I__5365 (
            .O(N__32675),
            .I(N__32669));
    InMux I__5364 (
            .O(N__32674),
            .I(N__32666));
    LocalMux I__5363 (
            .O(N__32669),
            .I(\reset_module_System.reset6_15 ));
    LocalMux I__5362 (
            .O(N__32666),
            .I(\reset_module_System.reset6_15 ));
    CascadeMux I__5361 (
            .O(N__32661),
            .I(\reset_module_System.reset6_19_cascade_ ));
    InMux I__5360 (
            .O(N__32658),
            .I(N__32655));
    LocalMux I__5359 (
            .O(N__32655),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    InMux I__5358 (
            .O(N__32652),
            .I(N__32649));
    LocalMux I__5357 (
            .O(N__32649),
            .I(N__32646));
    Odrv4 I__5356 (
            .O(N__32646),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    InMux I__5355 (
            .O(N__32643),
            .I(N__32639));
    CascadeMux I__5354 (
            .O(N__32642),
            .I(N__32636));
    LocalMux I__5353 (
            .O(N__32639),
            .I(N__32633));
    InMux I__5352 (
            .O(N__32636),
            .I(N__32630));
    Odrv4 I__5351 (
            .O(N__32633),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__5350 (
            .O(N__32630),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    InMux I__5349 (
            .O(N__32625),
            .I(N__32621));
    InMux I__5348 (
            .O(N__32624),
            .I(N__32618));
    LocalMux I__5347 (
            .O(N__32621),
            .I(\uart_drone.N_126_li ));
    LocalMux I__5346 (
            .O(N__32618),
            .I(\uart_drone.N_126_li ));
    CascadeMux I__5345 (
            .O(N__32613),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    InMux I__5344 (
            .O(N__32610),
            .I(N__32603));
    InMux I__5343 (
            .O(N__32609),
            .I(N__32599));
    InMux I__5342 (
            .O(N__32608),
            .I(N__32592));
    InMux I__5341 (
            .O(N__32607),
            .I(N__32592));
    InMux I__5340 (
            .O(N__32606),
            .I(N__32592));
    LocalMux I__5339 (
            .O(N__32603),
            .I(N__32589));
    InMux I__5338 (
            .O(N__32602),
            .I(N__32586));
    LocalMux I__5337 (
            .O(N__32599),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__5336 (
            .O(N__32592),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__5335 (
            .O(N__32589),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__5334 (
            .O(N__32586),
            .I(\uart_drone.stateZ0Z_4 ));
    InMux I__5333 (
            .O(N__32577),
            .I(N__32571));
    InMux I__5332 (
            .O(N__32576),
            .I(N__32571));
    LocalMux I__5331 (
            .O(N__32571),
            .I(\uart_drone.stateZ0Z_0 ));
    CascadeMux I__5330 (
            .O(N__32568),
            .I(N__32563));
    InMux I__5329 (
            .O(N__32567),
            .I(N__32560));
    InMux I__5328 (
            .O(N__32566),
            .I(N__32555));
    InMux I__5327 (
            .O(N__32563),
            .I(N__32555));
    LocalMux I__5326 (
            .O(N__32560),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__5325 (
            .O(N__32555),
            .I(\uart_drone.stateZ0Z_1 ));
    CascadeMux I__5324 (
            .O(N__32550),
            .I(\reset_module_System.reset6_15_cascade_ ));
    CascadeMux I__5323 (
            .O(N__32547),
            .I(\reset_module_System.count_1_1_cascade_ ));
    InMux I__5322 (
            .O(N__32544),
            .I(N__32541));
    LocalMux I__5321 (
            .O(N__32541),
            .I(N__32538));
    Odrv4 I__5320 (
            .O(N__32538),
            .I(\pid_front.error_p_reg_esr_RNI8NB61Z0Z_11 ));
    CascadeMux I__5319 (
            .O(N__32535),
            .I(\uart_drone.N_145_cascade_ ));
    CascadeMux I__5318 (
            .O(N__32532),
            .I(\uart_drone.un1_state_4_0_cascade_ ));
    CascadeMux I__5317 (
            .O(N__32529),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    InMux I__5316 (
            .O(N__32526),
            .I(N__32520));
    InMux I__5315 (
            .O(N__32525),
            .I(N__32520));
    LocalMux I__5314 (
            .O(N__32520),
            .I(N__32515));
    InMux I__5313 (
            .O(N__32519),
            .I(N__32510));
    InMux I__5312 (
            .O(N__32518),
            .I(N__32510));
    Odrv4 I__5311 (
            .O(N__32515),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__5310 (
            .O(N__32510),
            .I(\uart_drone.stateZ0Z_2 ));
    CascadeMux I__5309 (
            .O(N__32505),
            .I(N__32501));
    InMux I__5308 (
            .O(N__32504),
            .I(N__32495));
    InMux I__5307 (
            .O(N__32501),
            .I(N__32495));
    InMux I__5306 (
            .O(N__32500),
            .I(N__32492));
    LocalMux I__5305 (
            .O(N__32495),
            .I(N__32487));
    LocalMux I__5304 (
            .O(N__32492),
            .I(N__32484));
    InMux I__5303 (
            .O(N__32491),
            .I(N__32481));
    CascadeMux I__5302 (
            .O(N__32490),
            .I(N__32478));
    Span4Mux_v I__5301 (
            .O(N__32487),
            .I(N__32475));
    Span4Mux_h I__5300 (
            .O(N__32484),
            .I(N__32472));
    LocalMux I__5299 (
            .O(N__32481),
            .I(N__32469));
    InMux I__5298 (
            .O(N__32478),
            .I(N__32466));
    Odrv4 I__5297 (
            .O(N__32475),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    Odrv4 I__5296 (
            .O(N__32472),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    Odrv4 I__5295 (
            .O(N__32469),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__5294 (
            .O(N__32466),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    CascadeMux I__5293 (
            .O(N__32457),
            .I(\pid_front.un1_pid_prereg_48_cascade_ ));
    CascadeMux I__5292 (
            .O(N__32454),
            .I(N__32451));
    InMux I__5291 (
            .O(N__32451),
            .I(N__32445));
    InMux I__5290 (
            .O(N__32450),
            .I(N__32445));
    LocalMux I__5289 (
            .O(N__32445),
            .I(\pid_front.error_d_reg_prevZ0Z_19 ));
    InMux I__5288 (
            .O(N__32442),
            .I(N__32436));
    InMux I__5287 (
            .O(N__32441),
            .I(N__32436));
    LocalMux I__5286 (
            .O(N__32436),
            .I(N__32433));
    Span4Mux_v I__5285 (
            .O(N__32433),
            .I(N__32430));
    Span4Mux_v I__5284 (
            .O(N__32430),
            .I(N__32427));
    Sp12to4 I__5283 (
            .O(N__32427),
            .I(N__32424));
    Odrv12 I__5282 (
            .O(N__32424),
            .I(\pid_front.error_p_regZ0Z_19 ));
    InMux I__5281 (
            .O(N__32421),
            .I(N__32418));
    LocalMux I__5280 (
            .O(N__32418),
            .I(N__32414));
    InMux I__5279 (
            .O(N__32417),
            .I(N__32411));
    Odrv4 I__5278 (
            .O(N__32414),
            .I(\pid_front.un1_pid_prereg_56 ));
    LocalMux I__5277 (
            .O(N__32411),
            .I(\pid_front.un1_pid_prereg_56 ));
    CascadeMux I__5276 (
            .O(N__32406),
            .I(\pid_front.un1_pid_prereg_56_cascade_ ));
    InMux I__5275 (
            .O(N__32403),
            .I(N__32400));
    LocalMux I__5274 (
            .O(N__32400),
            .I(N__32396));
    InMux I__5273 (
            .O(N__32399),
            .I(N__32393));
    Odrv4 I__5272 (
            .O(N__32396),
            .I(\pid_front.un1_pid_prereg_48 ));
    LocalMux I__5271 (
            .O(N__32393),
            .I(\pid_front.un1_pid_prereg_48 ));
    InMux I__5270 (
            .O(N__32388),
            .I(N__32385));
    LocalMux I__5269 (
            .O(N__32385),
            .I(N__32382));
    Odrv4 I__5268 (
            .O(N__32382),
            .I(\pid_front.N_1471_i ));
    InMux I__5267 (
            .O(N__32379),
            .I(N__32372));
    InMux I__5266 (
            .O(N__32378),
            .I(N__32372));
    InMux I__5265 (
            .O(N__32377),
            .I(N__32369));
    LocalMux I__5264 (
            .O(N__32372),
            .I(N__32364));
    LocalMux I__5263 (
            .O(N__32369),
            .I(N__32364));
    Odrv4 I__5262 (
            .O(N__32364),
            .I(\pid_front.error_p_reg_esr_RNIA93NZ0Z_12 ));
    InMux I__5261 (
            .O(N__32361),
            .I(N__32352));
    InMux I__5260 (
            .O(N__32360),
            .I(N__32352));
    InMux I__5259 (
            .O(N__32359),
            .I(N__32352));
    LocalMux I__5258 (
            .O(N__32352),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    InMux I__5257 (
            .O(N__32349),
            .I(N__32344));
    InMux I__5256 (
            .O(N__32348),
            .I(N__32339));
    InMux I__5255 (
            .O(N__32347),
            .I(N__32339));
    LocalMux I__5254 (
            .O(N__32344),
            .I(N__32334));
    LocalMux I__5253 (
            .O(N__32339),
            .I(N__32334));
    Span12Mux_v I__5252 (
            .O(N__32334),
            .I(N__32331));
    Odrv12 I__5251 (
            .O(N__32331),
            .I(\pid_front.error_p_regZ0Z_12 ));
    CascadeMux I__5250 (
            .O(N__32328),
            .I(\pid_front.un1_pid_prereg_107_0_cascade_ ));
    InMux I__5249 (
            .O(N__32325),
            .I(N__32322));
    LocalMux I__5248 (
            .O(N__32322),
            .I(drone_altitude_1));
    InMux I__5247 (
            .O(N__32319),
            .I(N__32316));
    LocalMux I__5246 (
            .O(N__32316),
            .I(N__32313));
    Odrv12 I__5245 (
            .O(N__32313),
            .I(\pid_alt.error_axbZ0Z_1 ));
    CascadeMux I__5244 (
            .O(N__32310),
            .I(N__32306));
    InMux I__5243 (
            .O(N__32309),
            .I(N__32301));
    InMux I__5242 (
            .O(N__32306),
            .I(N__32296));
    InMux I__5241 (
            .O(N__32305),
            .I(N__32296));
    InMux I__5240 (
            .O(N__32304),
            .I(N__32293));
    LocalMux I__5239 (
            .O(N__32301),
            .I(N__32288));
    LocalMux I__5238 (
            .O(N__32296),
            .I(N__32288));
    LocalMux I__5237 (
            .O(N__32293),
            .I(N__32285));
    Span4Mux_v I__5236 (
            .O(N__32288),
            .I(N__32282));
    Span4Mux_v I__5235 (
            .O(N__32285),
            .I(N__32277));
    Span4Mux_h I__5234 (
            .O(N__32282),
            .I(N__32277));
    Span4Mux_h I__5233 (
            .O(N__32277),
            .I(N__32274));
    Odrv4 I__5232 (
            .O(N__32274),
            .I(\pid_front.error_p_regZ0Z_8 ));
    InMux I__5231 (
            .O(N__32271),
            .I(N__32268));
    LocalMux I__5230 (
            .O(N__32268),
            .I(N__32263));
    InMux I__5229 (
            .O(N__32267),
            .I(N__32257));
    InMux I__5228 (
            .O(N__32266),
            .I(N__32257));
    Span4Mux_v I__5227 (
            .O(N__32263),
            .I(N__32254));
    InMux I__5226 (
            .O(N__32262),
            .I(N__32251));
    LocalMux I__5225 (
            .O(N__32257),
            .I(N__32248));
    Span4Mux_h I__5224 (
            .O(N__32254),
            .I(N__32243));
    LocalMux I__5223 (
            .O(N__32251),
            .I(N__32243));
    Span4Mux_v I__5222 (
            .O(N__32248),
            .I(N__32240));
    Odrv4 I__5221 (
            .O(N__32243),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    Odrv4 I__5220 (
            .O(N__32240),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    CascadeMux I__5219 (
            .O(N__32235),
            .I(N__32232));
    InMux I__5218 (
            .O(N__32232),
            .I(N__32229));
    LocalMux I__5217 (
            .O(N__32229),
            .I(\pid_front.un1_pid_prereg_80_0 ));
    InMux I__5216 (
            .O(N__32226),
            .I(N__32223));
    LocalMux I__5215 (
            .O(N__32223),
            .I(\pid_front.N_1455_i ));
    CascadeMux I__5214 (
            .O(N__32220),
            .I(\pid_front.error_p_reg_esr_RNI8NB61Z0Z_11_cascade_ ));
    CascadeMux I__5213 (
            .O(N__32217),
            .I(\pid_front.un1_pid_prereg_57_cascade_ ));
    InMux I__5212 (
            .O(N__32214),
            .I(N__32209));
    InMux I__5211 (
            .O(N__32213),
            .I(N__32203));
    InMux I__5210 (
            .O(N__32212),
            .I(N__32200));
    LocalMux I__5209 (
            .O(N__32209),
            .I(N__32197));
    InMux I__5208 (
            .O(N__32208),
            .I(N__32192));
    InMux I__5207 (
            .O(N__32207),
            .I(N__32192));
    InMux I__5206 (
            .O(N__32206),
            .I(N__32189));
    LocalMux I__5205 (
            .O(N__32203),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__5204 (
            .O(N__32200),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv4 I__5203 (
            .O(N__32197),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__5202 (
            .O(N__32192),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__5201 (
            .O(N__32189),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    CascadeMux I__5200 (
            .O(N__32178),
            .I(N__32174));
    CascadeMux I__5199 (
            .O(N__32177),
            .I(N__32171));
    InMux I__5198 (
            .O(N__32174),
            .I(N__32167));
    InMux I__5197 (
            .O(N__32171),
            .I(N__32164));
    InMux I__5196 (
            .O(N__32170),
            .I(N__32161));
    LocalMux I__5195 (
            .O(N__32167),
            .I(N__32156));
    LocalMux I__5194 (
            .O(N__32164),
            .I(N__32156));
    LocalMux I__5193 (
            .O(N__32161),
            .I(N__32151));
    Span4Mux_v I__5192 (
            .O(N__32156),
            .I(N__32151));
    Odrv4 I__5191 (
            .O(N__32151),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    InMux I__5190 (
            .O(N__32148),
            .I(N__32145));
    LocalMux I__5189 (
            .O(N__32145),
            .I(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ));
    InMux I__5188 (
            .O(N__32142),
            .I(N__32139));
    LocalMux I__5187 (
            .O(N__32139),
            .I(N__32136));
    Odrv12 I__5186 (
            .O(N__32136),
            .I(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ));
    CascadeMux I__5185 (
            .O(N__32133),
            .I(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ));
    InMux I__5184 (
            .O(N__32130),
            .I(N__32127));
    LocalMux I__5183 (
            .O(N__32127),
            .I(\dron_frame_decoder_1.drone_H_disp_side_9 ));
    CascadeMux I__5182 (
            .O(N__32124),
            .I(\dron_frame_decoder_1.N_198_cascade_ ));
    InMux I__5181 (
            .O(N__32121),
            .I(N__32118));
    LocalMux I__5180 (
            .O(N__32118),
            .I(\dron_frame_decoder_1.N_200 ));
    InMux I__5179 (
            .O(N__32115),
            .I(N__32112));
    LocalMux I__5178 (
            .O(N__32112),
            .I(N__32108));
    InMux I__5177 (
            .O(N__32111),
            .I(N__32105));
    Span4Mux_s3_h I__5176 (
            .O(N__32108),
            .I(N__32102));
    LocalMux I__5175 (
            .O(N__32105),
            .I(N__32099));
    Span4Mux_h I__5174 (
            .O(N__32102),
            .I(N__32096));
    Span4Mux_s1_h I__5173 (
            .O(N__32099),
            .I(N__32093));
    Span4Mux_h I__5172 (
            .O(N__32096),
            .I(N__32090));
    Span4Mux_h I__5171 (
            .O(N__32093),
            .I(N__32087));
    Span4Mux_h I__5170 (
            .O(N__32090),
            .I(N__32084));
    Span4Mux_h I__5169 (
            .O(N__32087),
            .I(N__32081));
    Odrv4 I__5168 (
            .O(N__32084),
            .I(xy_kp_0));
    Odrv4 I__5167 (
            .O(N__32081),
            .I(xy_kp_0));
    InMux I__5166 (
            .O(N__32076),
            .I(N__32072));
    InMux I__5165 (
            .O(N__32075),
            .I(N__32069));
    LocalMux I__5164 (
            .O(N__32072),
            .I(N__32066));
    LocalMux I__5163 (
            .O(N__32069),
            .I(N__32063));
    Span4Mux_s2_h I__5162 (
            .O(N__32066),
            .I(N__32060));
    Span12Mux_s4_h I__5161 (
            .O(N__32063),
            .I(N__32057));
    Span4Mux_h I__5160 (
            .O(N__32060),
            .I(N__32054));
    Span12Mux_h I__5159 (
            .O(N__32057),
            .I(N__32051));
    Span4Mux_h I__5158 (
            .O(N__32054),
            .I(N__32048));
    Odrv12 I__5157 (
            .O(N__32051),
            .I(xy_kp_1));
    Odrv4 I__5156 (
            .O(N__32048),
            .I(xy_kp_1));
    InMux I__5155 (
            .O(N__32043),
            .I(N__32040));
    LocalMux I__5154 (
            .O(N__32040),
            .I(N__32037));
    Span4Mux_s3_h I__5153 (
            .O(N__32037),
            .I(N__32034));
    Span4Mux_h I__5152 (
            .O(N__32034),
            .I(N__32030));
    InMux I__5151 (
            .O(N__32033),
            .I(N__32027));
    Span4Mux_h I__5150 (
            .O(N__32030),
            .I(N__32024));
    LocalMux I__5149 (
            .O(N__32027),
            .I(N__32021));
    Span4Mux_h I__5148 (
            .O(N__32024),
            .I(N__32018));
    Span12Mux_s9_h I__5147 (
            .O(N__32021),
            .I(N__32015));
    Odrv4 I__5146 (
            .O(N__32018),
            .I(xy_kp_2));
    Odrv12 I__5145 (
            .O(N__32015),
            .I(xy_kp_2));
    InMux I__5144 (
            .O(N__32010),
            .I(N__32007));
    LocalMux I__5143 (
            .O(N__32007),
            .I(N__32003));
    InMux I__5142 (
            .O(N__32006),
            .I(N__32000));
    Span4Mux_s3_h I__5141 (
            .O(N__32003),
            .I(N__31997));
    LocalMux I__5140 (
            .O(N__32000),
            .I(N__31994));
    Span4Mux_h I__5139 (
            .O(N__31997),
            .I(N__31991));
    Span4Mux_v I__5138 (
            .O(N__31994),
            .I(N__31988));
    Span4Mux_h I__5137 (
            .O(N__31991),
            .I(N__31985));
    Span4Mux_h I__5136 (
            .O(N__31988),
            .I(N__31982));
    Span4Mux_h I__5135 (
            .O(N__31985),
            .I(N__31979));
    Span4Mux_h I__5134 (
            .O(N__31982),
            .I(N__31976));
    Odrv4 I__5133 (
            .O(N__31979),
            .I(xy_kp_3));
    Odrv4 I__5132 (
            .O(N__31976),
            .I(xy_kp_3));
    InMux I__5131 (
            .O(N__31971),
            .I(N__31968));
    LocalMux I__5130 (
            .O(N__31968),
            .I(N__31964));
    InMux I__5129 (
            .O(N__31967),
            .I(N__31961));
    Span4Mux_s3_h I__5128 (
            .O(N__31964),
            .I(N__31958));
    LocalMux I__5127 (
            .O(N__31961),
            .I(N__31955));
    Span4Mux_h I__5126 (
            .O(N__31958),
            .I(N__31952));
    Span4Mux_s1_h I__5125 (
            .O(N__31955),
            .I(N__31949));
    Span4Mux_h I__5124 (
            .O(N__31952),
            .I(N__31946));
    Span4Mux_h I__5123 (
            .O(N__31949),
            .I(N__31943));
    Span4Mux_h I__5122 (
            .O(N__31946),
            .I(N__31940));
    Span4Mux_h I__5121 (
            .O(N__31943),
            .I(N__31937));
    Odrv4 I__5120 (
            .O(N__31940),
            .I(xy_kp_7));
    Odrv4 I__5119 (
            .O(N__31937),
            .I(xy_kp_7));
    CEMux I__5118 (
            .O(N__31932),
            .I(N__31929));
    LocalMux I__5117 (
            .O(N__31929),
            .I(N__31926));
    Span4Mux_v I__5116 (
            .O(N__31926),
            .I(N__31922));
    CEMux I__5115 (
            .O(N__31925),
            .I(N__31919));
    Odrv4 I__5114 (
            .O(N__31922),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    LocalMux I__5113 (
            .O(N__31919),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    CascadeMux I__5112 (
            .O(N__31914),
            .I(N__31910));
    InMux I__5111 (
            .O(N__31913),
            .I(N__31901));
    InMux I__5110 (
            .O(N__31910),
            .I(N__31901));
    InMux I__5109 (
            .O(N__31909),
            .I(N__31901));
    InMux I__5108 (
            .O(N__31908),
            .I(N__31898));
    LocalMux I__5107 (
            .O(N__31901),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__5106 (
            .O(N__31898),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    InMux I__5105 (
            .O(N__31893),
            .I(N__31890));
    LocalMux I__5104 (
            .O(N__31890),
            .I(\dron_frame_decoder_1.state_ns_i_a2_0_0_0 ));
    InMux I__5103 (
            .O(N__31887),
            .I(N__31880));
    InMux I__5102 (
            .O(N__31886),
            .I(N__31880));
    InMux I__5101 (
            .O(N__31885),
            .I(N__31877));
    LocalMux I__5100 (
            .O(N__31880),
            .I(N__31874));
    LocalMux I__5099 (
            .O(N__31877),
            .I(\uart_drone.data_rdyc_1 ));
    Odrv4 I__5098 (
            .O(N__31874),
            .I(\uart_drone.data_rdyc_1 ));
    CascadeMux I__5097 (
            .O(N__31869),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ));
    CascadeMux I__5096 (
            .O(N__31866),
            .I(N__31861));
    InMux I__5095 (
            .O(N__31865),
            .I(N__31858));
    InMux I__5094 (
            .O(N__31864),
            .I(N__31853));
    InMux I__5093 (
            .O(N__31861),
            .I(N__31853));
    LocalMux I__5092 (
            .O(N__31858),
            .I(N__31850));
    LocalMux I__5091 (
            .O(N__31853),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    Odrv4 I__5090 (
            .O(N__31850),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    InMux I__5089 (
            .O(N__31845),
            .I(N__31842));
    LocalMux I__5088 (
            .O(N__31842),
            .I(N__31837));
    InMux I__5087 (
            .O(N__31841),
            .I(N__31832));
    InMux I__5086 (
            .O(N__31840),
            .I(N__31832));
    Span4Mux_h I__5085 (
            .O(N__31837),
            .I(N__31826));
    LocalMux I__5084 (
            .O(N__31832),
            .I(N__31826));
    InMux I__5083 (
            .O(N__31831),
            .I(N__31823));
    Odrv4 I__5082 (
            .O(N__31826),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    LocalMux I__5081 (
            .O(N__31823),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    InMux I__5080 (
            .O(N__31818),
            .I(N__31815));
    LocalMux I__5079 (
            .O(N__31815),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    InMux I__5078 (
            .O(N__31812),
            .I(N__31809));
    LocalMux I__5077 (
            .O(N__31809),
            .I(N__31805));
    InMux I__5076 (
            .O(N__31808),
            .I(N__31801));
    Span4Mux_v I__5075 (
            .O(N__31805),
            .I(N__31798));
    InMux I__5074 (
            .O(N__31804),
            .I(N__31795));
    LocalMux I__5073 (
            .O(N__31801),
            .I(N__31790));
    Span4Mux_h I__5072 (
            .O(N__31798),
            .I(N__31790));
    LocalMux I__5071 (
            .O(N__31795),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    Odrv4 I__5070 (
            .O(N__31790),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    CascadeMux I__5069 (
            .O(N__31785),
            .I(N__31768));
    InMux I__5068 (
            .O(N__31784),
            .I(N__31759));
    InMux I__5067 (
            .O(N__31783),
            .I(N__31754));
    InMux I__5066 (
            .O(N__31782),
            .I(N__31754));
    InMux I__5065 (
            .O(N__31781),
            .I(N__31747));
    InMux I__5064 (
            .O(N__31780),
            .I(N__31747));
    InMux I__5063 (
            .O(N__31779),
            .I(N__31747));
    InMux I__5062 (
            .O(N__31778),
            .I(N__31742));
    InMux I__5061 (
            .O(N__31777),
            .I(N__31742));
    InMux I__5060 (
            .O(N__31776),
            .I(N__31735));
    InMux I__5059 (
            .O(N__31775),
            .I(N__31732));
    CascadeMux I__5058 (
            .O(N__31774),
            .I(N__31729));
    InMux I__5057 (
            .O(N__31773),
            .I(N__31722));
    InMux I__5056 (
            .O(N__31772),
            .I(N__31719));
    InMux I__5055 (
            .O(N__31771),
            .I(N__31716));
    InMux I__5054 (
            .O(N__31768),
            .I(N__31713));
    InMux I__5053 (
            .O(N__31767),
            .I(N__31704));
    InMux I__5052 (
            .O(N__31766),
            .I(N__31704));
    InMux I__5051 (
            .O(N__31765),
            .I(N__31704));
    InMux I__5050 (
            .O(N__31764),
            .I(N__31704));
    InMux I__5049 (
            .O(N__31763),
            .I(N__31701));
    InMux I__5048 (
            .O(N__31762),
            .I(N__31698));
    LocalMux I__5047 (
            .O(N__31759),
            .I(N__31695));
    LocalMux I__5046 (
            .O(N__31754),
            .I(N__31690));
    LocalMux I__5045 (
            .O(N__31747),
            .I(N__31690));
    LocalMux I__5044 (
            .O(N__31742),
            .I(N__31687));
    InMux I__5043 (
            .O(N__31741),
            .I(N__31680));
    InMux I__5042 (
            .O(N__31740),
            .I(N__31680));
    InMux I__5041 (
            .O(N__31739),
            .I(N__31680));
    CascadeMux I__5040 (
            .O(N__31738),
            .I(N__31675));
    LocalMux I__5039 (
            .O(N__31735),
            .I(N__31671));
    LocalMux I__5038 (
            .O(N__31732),
            .I(N__31668));
    InMux I__5037 (
            .O(N__31729),
            .I(N__31663));
    InMux I__5036 (
            .O(N__31728),
            .I(N__31663));
    InMux I__5035 (
            .O(N__31727),
            .I(N__31656));
    InMux I__5034 (
            .O(N__31726),
            .I(N__31656));
    InMux I__5033 (
            .O(N__31725),
            .I(N__31656));
    LocalMux I__5032 (
            .O(N__31722),
            .I(N__31650));
    LocalMux I__5031 (
            .O(N__31719),
            .I(N__31650));
    LocalMux I__5030 (
            .O(N__31716),
            .I(N__31647));
    LocalMux I__5029 (
            .O(N__31713),
            .I(N__31634));
    LocalMux I__5028 (
            .O(N__31704),
            .I(N__31634));
    LocalMux I__5027 (
            .O(N__31701),
            .I(N__31634));
    LocalMux I__5026 (
            .O(N__31698),
            .I(N__31634));
    Span4Mux_h I__5025 (
            .O(N__31695),
            .I(N__31634));
    Span4Mux_v I__5024 (
            .O(N__31690),
            .I(N__31634));
    Span4Mux_h I__5023 (
            .O(N__31687),
            .I(N__31629));
    LocalMux I__5022 (
            .O(N__31680),
            .I(N__31629));
    InMux I__5021 (
            .O(N__31679),
            .I(N__31626));
    InMux I__5020 (
            .O(N__31678),
            .I(N__31621));
    InMux I__5019 (
            .O(N__31675),
            .I(N__31621));
    InMux I__5018 (
            .O(N__31674),
            .I(N__31618));
    Span4Mux_v I__5017 (
            .O(N__31671),
            .I(N__31613));
    Span4Mux_v I__5016 (
            .O(N__31668),
            .I(N__31613));
    LocalMux I__5015 (
            .O(N__31663),
            .I(N__31608));
    LocalMux I__5014 (
            .O(N__31656),
            .I(N__31608));
    InMux I__5013 (
            .O(N__31655),
            .I(N__31605));
    Span4Mux_v I__5012 (
            .O(N__31650),
            .I(N__31596));
    Span4Mux_v I__5011 (
            .O(N__31647),
            .I(N__31596));
    Span4Mux_v I__5010 (
            .O(N__31634),
            .I(N__31596));
    Span4Mux_v I__5009 (
            .O(N__31629),
            .I(N__31596));
    LocalMux I__5008 (
            .O(N__31626),
            .I(uart_pc_data_rdy));
    LocalMux I__5007 (
            .O(N__31621),
            .I(uart_pc_data_rdy));
    LocalMux I__5006 (
            .O(N__31618),
            .I(uart_pc_data_rdy));
    Odrv4 I__5005 (
            .O(N__31613),
            .I(uart_pc_data_rdy));
    Odrv12 I__5004 (
            .O(N__31608),
            .I(uart_pc_data_rdy));
    LocalMux I__5003 (
            .O(N__31605),
            .I(uart_pc_data_rdy));
    Odrv4 I__5002 (
            .O(N__31596),
            .I(uart_pc_data_rdy));
    CascadeMux I__5001 (
            .O(N__31581),
            .I(\dron_frame_decoder_1.state_ns_0_a3_0_1Z0Z_1_cascade_ ));
    InMux I__5000 (
            .O(N__31578),
            .I(N__31575));
    LocalMux I__4999 (
            .O(N__31575),
            .I(\dron_frame_decoder_1.N_220 ));
    CascadeMux I__4998 (
            .O(N__31572),
            .I(\dron_frame_decoder_1.N_220_cascade_ ));
    CascadeMux I__4997 (
            .O(N__31569),
            .I(N__31566));
    InMux I__4996 (
            .O(N__31566),
            .I(N__31560));
    InMux I__4995 (
            .O(N__31565),
            .I(N__31560));
    LocalMux I__4994 (
            .O(N__31560),
            .I(\dron_frame_decoder_1.N_224 ));
    InMux I__4993 (
            .O(N__31557),
            .I(N__31553));
    InMux I__4992 (
            .O(N__31556),
            .I(N__31550));
    LocalMux I__4991 (
            .O(N__31553),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    LocalMux I__4990 (
            .O(N__31550),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    CascadeMux I__4989 (
            .O(N__31545),
            .I(N__31540));
    InMux I__4988 (
            .O(N__31544),
            .I(N__31534));
    InMux I__4987 (
            .O(N__31543),
            .I(N__31534));
    InMux I__4986 (
            .O(N__31540),
            .I(N__31529));
    InMux I__4985 (
            .O(N__31539),
            .I(N__31529));
    LocalMux I__4984 (
            .O(N__31534),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__4983 (
            .O(N__31529),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    CascadeMux I__4982 (
            .O(N__31524),
            .I(N__31521));
    InMux I__4981 (
            .O(N__31521),
            .I(N__31518));
    LocalMux I__4980 (
            .O(N__31518),
            .I(N__31515));
    Odrv4 I__4979 (
            .O(N__31515),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    InMux I__4978 (
            .O(N__31512),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__4977 (
            .O(N__31509),
            .I(N__31506));
    LocalMux I__4976 (
            .O(N__31506),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__4975 (
            .O(N__31503),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__4974 (
            .O(N__31500),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__4973 (
            .O(N__31497),
            .I(N__31494));
    LocalMux I__4972 (
            .O(N__31494),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    InMux I__4971 (
            .O(N__31491),
            .I(N__31488));
    LocalMux I__4970 (
            .O(N__31488),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__4969 (
            .O(N__31485),
            .I(N__31478));
    InMux I__4968 (
            .O(N__31484),
            .I(N__31475));
    InMux I__4967 (
            .O(N__31483),
            .I(N__31472));
    InMux I__4966 (
            .O(N__31482),
            .I(N__31467));
    InMux I__4965 (
            .O(N__31481),
            .I(N__31467));
    LocalMux I__4964 (
            .O(N__31478),
            .I(\uart_drone.N_143 ));
    LocalMux I__4963 (
            .O(N__31475),
            .I(\uart_drone.N_143 ));
    LocalMux I__4962 (
            .O(N__31472),
            .I(\uart_drone.N_143 ));
    LocalMux I__4961 (
            .O(N__31467),
            .I(\uart_drone.N_143 ));
    CascadeMux I__4960 (
            .O(N__31458),
            .I(N__31454));
    InMux I__4959 (
            .O(N__31457),
            .I(N__31450));
    InMux I__4958 (
            .O(N__31454),
            .I(N__31445));
    InMux I__4957 (
            .O(N__31453),
            .I(N__31445));
    LocalMux I__4956 (
            .O(N__31450),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__4955 (
            .O(N__31445),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    InMux I__4954 (
            .O(N__31440),
            .I(N__31437));
    LocalMux I__4953 (
            .O(N__31437),
            .I(N__31432));
    InMux I__4952 (
            .O(N__31436),
            .I(N__31429));
    InMux I__4951 (
            .O(N__31435),
            .I(N__31426));
    Odrv4 I__4950 (
            .O(N__31432),
            .I(\Commands_frame_decoder.preinitZ0 ));
    LocalMux I__4949 (
            .O(N__31429),
            .I(\Commands_frame_decoder.preinitZ0 ));
    LocalMux I__4948 (
            .O(N__31426),
            .I(\Commands_frame_decoder.preinitZ0 ));
    InMux I__4947 (
            .O(N__31419),
            .I(N__31415));
    InMux I__4946 (
            .O(N__31418),
            .I(N__31412));
    LocalMux I__4945 (
            .O(N__31415),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__4944 (
            .O(N__31412),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__4943 (
            .O(N__31407),
            .I(N__31402));
    InMux I__4942 (
            .O(N__31406),
            .I(N__31397));
    InMux I__4941 (
            .O(N__31405),
            .I(N__31397));
    LocalMux I__4940 (
            .O(N__31402),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__4939 (
            .O(N__31397),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    CascadeMux I__4938 (
            .O(N__31392),
            .I(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4_cascade_ ));
    InMux I__4937 (
            .O(N__31389),
            .I(N__31386));
    LocalMux I__4936 (
            .O(N__31386),
            .I(\Commands_frame_decoder.WDT8lto15_N_5L7_1 ));
    InMux I__4935 (
            .O(N__31383),
            .I(N__31380));
    LocalMux I__4934 (
            .O(N__31380),
            .I(\Commands_frame_decoder.WDT_RNIAERH3Z0Z_12 ));
    InMux I__4933 (
            .O(N__31377),
            .I(N__31372));
    InMux I__4932 (
            .O(N__31376),
            .I(N__31369));
    InMux I__4931 (
            .O(N__31375),
            .I(N__31366));
    LocalMux I__4930 (
            .O(N__31372),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__4929 (
            .O(N__31369),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__4928 (
            .O(N__31366),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    InMux I__4927 (
            .O(N__31359),
            .I(N__31353));
    InMux I__4926 (
            .O(N__31358),
            .I(N__31350));
    InMux I__4925 (
            .O(N__31357),
            .I(N__31345));
    InMux I__4924 (
            .O(N__31356),
            .I(N__31345));
    LocalMux I__4923 (
            .O(N__31353),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__4922 (
            .O(N__31350),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__4921 (
            .O(N__31345),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    CascadeMux I__4920 (
            .O(N__31338),
            .I(\Commands_frame_decoder.WDT_RNIAERH3Z0Z_12_cascade_ ));
    InMux I__4919 (
            .O(N__31335),
            .I(N__31330));
    InMux I__4918 (
            .O(N__31334),
            .I(N__31327));
    InMux I__4917 (
            .O(N__31333),
            .I(N__31324));
    LocalMux I__4916 (
            .O(N__31330),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__4915 (
            .O(N__31327),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__4914 (
            .O(N__31324),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    InMux I__4913 (
            .O(N__31317),
            .I(N__31310));
    InMux I__4912 (
            .O(N__31316),
            .I(N__31300));
    InMux I__4911 (
            .O(N__31315),
            .I(N__31297));
    InMux I__4910 (
            .O(N__31314),
            .I(N__31292));
    InMux I__4909 (
            .O(N__31313),
            .I(N__31292));
    LocalMux I__4908 (
            .O(N__31310),
            .I(N__31287));
    InMux I__4907 (
            .O(N__31309),
            .I(N__31280));
    InMux I__4906 (
            .O(N__31308),
            .I(N__31280));
    InMux I__4905 (
            .O(N__31307),
            .I(N__31280));
    InMux I__4904 (
            .O(N__31306),
            .I(N__31275));
    InMux I__4903 (
            .O(N__31305),
            .I(N__31275));
    InMux I__4902 (
            .O(N__31304),
            .I(N__31270));
    InMux I__4901 (
            .O(N__31303),
            .I(N__31270));
    LocalMux I__4900 (
            .O(N__31300),
            .I(N__31264));
    LocalMux I__4899 (
            .O(N__31297),
            .I(N__31264));
    LocalMux I__4898 (
            .O(N__31292),
            .I(N__31261));
    InMux I__4897 (
            .O(N__31291),
            .I(N__31256));
    InMux I__4896 (
            .O(N__31290),
            .I(N__31256));
    Span4Mux_v I__4895 (
            .O(N__31287),
            .I(N__31253));
    LocalMux I__4894 (
            .O(N__31280),
            .I(N__31248));
    LocalMux I__4893 (
            .O(N__31275),
            .I(N__31248));
    LocalMux I__4892 (
            .O(N__31270),
            .I(N__31245));
    InMux I__4891 (
            .O(N__31269),
            .I(N__31242));
    Span4Mux_v I__4890 (
            .O(N__31264),
            .I(N__31239));
    Span4Mux_v I__4889 (
            .O(N__31261),
            .I(N__31234));
    LocalMux I__4888 (
            .O(N__31256),
            .I(N__31234));
    Span4Mux_h I__4887 (
            .O(N__31253),
            .I(N__31225));
    Span4Mux_v I__4886 (
            .O(N__31248),
            .I(N__31225));
    Span4Mux_h I__4885 (
            .O(N__31245),
            .I(N__31225));
    LocalMux I__4884 (
            .O(N__31242),
            .I(N__31225));
    Span4Mux_h I__4883 (
            .O(N__31239),
            .I(N__31222));
    Span4Mux_v I__4882 (
            .O(N__31234),
            .I(N__31219));
    Span4Mux_v I__4881 (
            .O(N__31225),
            .I(N__31216));
    Odrv4 I__4880 (
            .O(N__31222),
            .I(\Commands_frame_decoder.WDT8_0 ));
    Odrv4 I__4879 (
            .O(N__31219),
            .I(\Commands_frame_decoder.WDT8_0 ));
    Odrv4 I__4878 (
            .O(N__31216),
            .I(\Commands_frame_decoder.WDT8_0 ));
    CascadeMux I__4877 (
            .O(N__31209),
            .I(\uart_drone.N_126_li_cascade_ ));
    CascadeMux I__4876 (
            .O(N__31206),
            .I(\uart_drone.N_143_cascade_ ));
    IoInMux I__4875 (
            .O(N__31203),
            .I(N__31200));
    LocalMux I__4874 (
            .O(N__31200),
            .I(N__31197));
    Span4Mux_s3_v I__4873 (
            .O(N__31197),
            .I(N__31194));
    Odrv4 I__4872 (
            .O(N__31194),
            .I(\pid_front.state_0_0 ));
    InMux I__4871 (
            .O(N__31191),
            .I(N__31188));
    LocalMux I__4870 (
            .O(N__31188),
            .I(uart_input_pc_c));
    InMux I__4869 (
            .O(N__31185),
            .I(N__31182));
    LocalMux I__4868 (
            .O(N__31182),
            .I(N__31179));
    Odrv4 I__4867 (
            .O(N__31179),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    InMux I__4866 (
            .O(N__31176),
            .I(N__31173));
    LocalMux I__4865 (
            .O(N__31173),
            .I(N__31170));
    Odrv4 I__4864 (
            .O(N__31170),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    CascadeMux I__4863 (
            .O(N__31167),
            .I(\Commands_frame_decoder.state_0_sqmuxa_1_cascade_ ));
    CascadeMux I__4862 (
            .O(N__31164),
            .I(N__31160));
    InMux I__4861 (
            .O(N__31163),
            .I(N__31157));
    InMux I__4860 (
            .O(N__31160),
            .I(N__31154));
    LocalMux I__4859 (
            .O(N__31157),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__4858 (
            .O(N__31154),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    InMux I__4857 (
            .O(N__31149),
            .I(N__31146));
    LocalMux I__4856 (
            .O(N__31146),
            .I(N__31143));
    Odrv4 I__4855 (
            .O(N__31143),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    InMux I__4854 (
            .O(N__31140),
            .I(N__31137));
    LocalMux I__4853 (
            .O(N__31137),
            .I(N__31134));
    Odrv4 I__4852 (
            .O(N__31134),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    InMux I__4851 (
            .O(N__31131),
            .I(N__31127));
    InMux I__4850 (
            .O(N__31130),
            .I(N__31124));
    LocalMux I__4849 (
            .O(N__31127),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__4848 (
            .O(N__31124),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    CascadeMux I__4847 (
            .O(N__31119),
            .I(N__31115));
    InMux I__4846 (
            .O(N__31118),
            .I(N__31112));
    InMux I__4845 (
            .O(N__31115),
            .I(N__31109));
    LocalMux I__4844 (
            .O(N__31112),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__4843 (
            .O(N__31109),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__4842 (
            .O(N__31104),
            .I(N__31100));
    InMux I__4841 (
            .O(N__31103),
            .I(N__31097));
    LocalMux I__4840 (
            .O(N__31100),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__4839 (
            .O(N__31097),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__4838 (
            .O(N__31092),
            .I(N__31088));
    InMux I__4837 (
            .O(N__31091),
            .I(N__31085));
    LocalMux I__4836 (
            .O(N__31088),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__4835 (
            .O(N__31085),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__4834 (
            .O(N__31080),
            .I(N__31076));
    InMux I__4833 (
            .O(N__31079),
            .I(N__31073));
    LocalMux I__4832 (
            .O(N__31076),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__4831 (
            .O(N__31073),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    CascadeMux I__4830 (
            .O(N__31068),
            .I(N__31064));
    InMux I__4829 (
            .O(N__31067),
            .I(N__31061));
    InMux I__4828 (
            .O(N__31064),
            .I(N__31058));
    LocalMux I__4827 (
            .O(N__31061),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__4826 (
            .O(N__31058),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    InMux I__4825 (
            .O(N__31053),
            .I(N__31049));
    InMux I__4824 (
            .O(N__31052),
            .I(N__31046));
    LocalMux I__4823 (
            .O(N__31049),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__4822 (
            .O(N__31046),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    CascadeMux I__4821 (
            .O(N__31041),
            .I(\pid_front.un1_pid_prereg_23_cascade_ ));
    CascadeMux I__4820 (
            .O(N__31038),
            .I(\pid_front.un1_pid_prereg_30_cascade_ ));
    InMux I__4819 (
            .O(N__31035),
            .I(N__31029));
    InMux I__4818 (
            .O(N__31034),
            .I(N__31029));
    LocalMux I__4817 (
            .O(N__31029),
            .I(N__31026));
    Span4Mux_v I__4816 (
            .O(N__31026),
            .I(N__31023));
    Span4Mux_v I__4815 (
            .O(N__31023),
            .I(N__31020));
    Span4Mux_h I__4814 (
            .O(N__31020),
            .I(N__31017));
    Odrv4 I__4813 (
            .O(N__31017),
            .I(\pid_front.error_p_regZ0Z_15 ));
    CascadeMux I__4812 (
            .O(N__31014),
            .I(N__31011));
    InMux I__4811 (
            .O(N__31011),
            .I(N__31005));
    InMux I__4810 (
            .O(N__31010),
            .I(N__31005));
    LocalMux I__4809 (
            .O(N__31005),
            .I(\pid_front.error_d_reg_prevZ0Z_15 ));
    InMux I__4808 (
            .O(N__31002),
            .I(N__30998));
    InMux I__4807 (
            .O(N__31001),
            .I(N__30995));
    LocalMux I__4806 (
            .O(N__30998),
            .I(\pid_front.un1_pid_prereg_29 ));
    LocalMux I__4805 (
            .O(N__30995),
            .I(\pid_front.un1_pid_prereg_29 ));
    CascadeMux I__4804 (
            .O(N__30990),
            .I(\pid_front.un1_pid_prereg_29_cascade_ ));
    InMux I__4803 (
            .O(N__30987),
            .I(N__30983));
    InMux I__4802 (
            .O(N__30986),
            .I(N__30980));
    LocalMux I__4801 (
            .O(N__30983),
            .I(N__30975));
    LocalMux I__4800 (
            .O(N__30980),
            .I(N__30975));
    Span4Mux_v I__4799 (
            .O(N__30975),
            .I(N__30972));
    Span4Mux_h I__4798 (
            .O(N__30972),
            .I(N__30969));
    Span4Mux_v I__4797 (
            .O(N__30969),
            .I(N__30966));
    Odrv4 I__4796 (
            .O(N__30966),
            .I(\pid_front.error_p_regZ0Z_14 ));
    InMux I__4795 (
            .O(N__30963),
            .I(N__30956));
    InMux I__4794 (
            .O(N__30962),
            .I(N__30956));
    InMux I__4793 (
            .O(N__30961),
            .I(N__30953));
    LocalMux I__4792 (
            .O(N__30956),
            .I(\pid_front.un1_pid_prereg_24 ));
    LocalMux I__4791 (
            .O(N__30953),
            .I(\pid_front.un1_pid_prereg_24 ));
    InMux I__4790 (
            .O(N__30948),
            .I(N__30945));
    LocalMux I__4789 (
            .O(N__30945),
            .I(N__30942));
    Span4Mux_v I__4788 (
            .O(N__30942),
            .I(N__30939));
    Span4Mux_h I__4787 (
            .O(N__30939),
            .I(N__30936));
    Span4Mux_h I__4786 (
            .O(N__30936),
            .I(N__30933));
    Odrv4 I__4785 (
            .O(N__30933),
            .I(\pid_front.O_0_11 ));
    CascadeMux I__4784 (
            .O(N__30930),
            .I(\pid_front.N_1451_i_cascade_ ));
    CascadeMux I__4783 (
            .O(N__30927),
            .I(\pid_front.error_d_reg_esr_RNINKUFZ0Z_7_cascade_ ));
    InMux I__4782 (
            .O(N__30924),
            .I(N__30921));
    LocalMux I__4781 (
            .O(N__30921),
            .I(\pid_front.un1_pid_prereg_70_0 ));
    InMux I__4780 (
            .O(N__30918),
            .I(N__30914));
    InMux I__4779 (
            .O(N__30917),
            .I(N__30911));
    LocalMux I__4778 (
            .O(N__30914),
            .I(N__30908));
    LocalMux I__4777 (
            .O(N__30911),
            .I(\pid_front.un1_pid_prereg_23 ));
    Odrv4 I__4776 (
            .O(N__30908),
            .I(\pid_front.un1_pid_prereg_23 ));
    InMux I__4775 (
            .O(N__30903),
            .I(N__30900));
    LocalMux I__4774 (
            .O(N__30900),
            .I(\dron_frame_decoder_1.drone_altitude_5 ));
    InMux I__4773 (
            .O(N__30897),
            .I(N__30894));
    LocalMux I__4772 (
            .O(N__30894),
            .I(\dron_frame_decoder_1.drone_altitude_6 ));
    InMux I__4771 (
            .O(N__30891),
            .I(N__30888));
    LocalMux I__4770 (
            .O(N__30888),
            .I(\dron_frame_decoder_1.drone_altitude_7 ));
    InMux I__4769 (
            .O(N__30885),
            .I(N__30882));
    LocalMux I__4768 (
            .O(N__30882),
            .I(\dron_frame_decoder_1.drone_altitude_8 ));
    InMux I__4767 (
            .O(N__30879),
            .I(N__30876));
    LocalMux I__4766 (
            .O(N__30876),
            .I(drone_altitude_14));
    InMux I__4765 (
            .O(N__30873),
            .I(N__30870));
    LocalMux I__4764 (
            .O(N__30870),
            .I(drone_altitude_13));
    InMux I__4763 (
            .O(N__30867),
            .I(N__30864));
    LocalMux I__4762 (
            .O(N__30864),
            .I(drone_altitude_12));
    CEMux I__4761 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__4760 (
            .O(N__30858),
            .I(N__30855));
    Span4Mux_h I__4759 (
            .O(N__30855),
            .I(N__30851));
    CEMux I__4758 (
            .O(N__30854),
            .I(N__30847));
    Span4Mux_h I__4757 (
            .O(N__30851),
            .I(N__30844));
    CEMux I__4756 (
            .O(N__30850),
            .I(N__30841));
    LocalMux I__4755 (
            .O(N__30847),
            .I(N__30838));
    Sp12to4 I__4754 (
            .O(N__30844),
            .I(N__30833));
    LocalMux I__4753 (
            .O(N__30841),
            .I(N__30833));
    Sp12to4 I__4752 (
            .O(N__30838),
            .I(N__30830));
    Odrv12 I__4751 (
            .O(N__30833),
            .I(\dron_frame_decoder_1.N_513_0 ));
    Odrv12 I__4750 (
            .O(N__30830),
            .I(\dron_frame_decoder_1.N_513_0 ));
    InMux I__4749 (
            .O(N__30825),
            .I(N__30820));
    InMux I__4748 (
            .O(N__30824),
            .I(N__30815));
    InMux I__4747 (
            .O(N__30823),
            .I(N__30815));
    LocalMux I__4746 (
            .O(N__30820),
            .I(N__30812));
    LocalMux I__4745 (
            .O(N__30815),
            .I(N__30809));
    Span4Mux_h I__4744 (
            .O(N__30812),
            .I(N__30806));
    Span4Mux_v I__4743 (
            .O(N__30809),
            .I(N__30803));
    Span4Mux_v I__4742 (
            .O(N__30806),
            .I(N__30800));
    Span4Mux_h I__4741 (
            .O(N__30803),
            .I(N__30797));
    Span4Mux_h I__4740 (
            .O(N__30800),
            .I(N__30794));
    Odrv4 I__4739 (
            .O(N__30797),
            .I(\pid_front.error_p_regZ0Z_9 ));
    Odrv4 I__4738 (
            .O(N__30794),
            .I(\pid_front.error_p_regZ0Z_9 ));
    InMux I__4737 (
            .O(N__30789),
            .I(N__30782));
    InMux I__4736 (
            .O(N__30788),
            .I(N__30782));
    InMux I__4735 (
            .O(N__30787),
            .I(N__30779));
    LocalMux I__4734 (
            .O(N__30782),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    LocalMux I__4733 (
            .O(N__30779),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    InMux I__4732 (
            .O(N__30774),
            .I(N__30771));
    LocalMux I__4731 (
            .O(N__30771),
            .I(N__30768));
    Span4Mux_v I__4730 (
            .O(N__30768),
            .I(N__30765));
    Odrv4 I__4729 (
            .O(N__30765),
            .I(\pid_front.N_1459_i ));
    InMux I__4728 (
            .O(N__30762),
            .I(N__30759));
    LocalMux I__4727 (
            .O(N__30759),
            .I(N__30755));
    InMux I__4726 (
            .O(N__30758),
            .I(N__30752));
    Span4Mux_v I__4725 (
            .O(N__30755),
            .I(N__30749));
    LocalMux I__4724 (
            .O(N__30752),
            .I(N__30746));
    Sp12to4 I__4723 (
            .O(N__30749),
            .I(N__30743));
    Span4Mux_h I__4722 (
            .O(N__30746),
            .I(N__30740));
    Span12Mux_s11_h I__4721 (
            .O(N__30743),
            .I(N__30737));
    Span4Mux_h I__4720 (
            .O(N__30740),
            .I(N__30734));
    Odrv12 I__4719 (
            .O(N__30737),
            .I(xy_kp_6));
    Odrv4 I__4718 (
            .O(N__30734),
            .I(xy_kp_6));
    InMux I__4717 (
            .O(N__30729),
            .I(N__30726));
    LocalMux I__4716 (
            .O(N__30726),
            .I(N__30723));
    Span4Mux_v I__4715 (
            .O(N__30723),
            .I(N__30719));
    InMux I__4714 (
            .O(N__30722),
            .I(N__30716));
    Span4Mux_h I__4713 (
            .O(N__30719),
            .I(N__30713));
    LocalMux I__4712 (
            .O(N__30716),
            .I(N__30710));
    Span4Mux_h I__4711 (
            .O(N__30713),
            .I(N__30707));
    Span4Mux_h I__4710 (
            .O(N__30710),
            .I(N__30704));
    Sp12to4 I__4709 (
            .O(N__30707),
            .I(N__30701));
    Span4Mux_h I__4708 (
            .O(N__30704),
            .I(N__30698));
    Odrv12 I__4707 (
            .O(N__30701),
            .I(xy_kp_5));
    Odrv4 I__4706 (
            .O(N__30698),
            .I(xy_kp_5));
    InMux I__4705 (
            .O(N__30693),
            .I(N__30690));
    LocalMux I__4704 (
            .O(N__30690),
            .I(N__30687));
    Span4Mux_v I__4703 (
            .O(N__30687),
            .I(N__30682));
    InMux I__4702 (
            .O(N__30686),
            .I(N__30679));
    InMux I__4701 (
            .O(N__30685),
            .I(N__30676));
    Span4Mux_v I__4700 (
            .O(N__30682),
            .I(N__30671));
    LocalMux I__4699 (
            .O(N__30679),
            .I(N__30671));
    LocalMux I__4698 (
            .O(N__30676),
            .I(N__30668));
    Span4Mux_h I__4697 (
            .O(N__30671),
            .I(N__30665));
    Span4Mux_v I__4696 (
            .O(N__30668),
            .I(N__30662));
    Span4Mux_h I__4695 (
            .O(N__30665),
            .I(N__30659));
    Sp12to4 I__4694 (
            .O(N__30662),
            .I(N__30656));
    Sp12to4 I__4693 (
            .O(N__30659),
            .I(N__30650));
    Span12Mux_s8_h I__4692 (
            .O(N__30656),
            .I(N__30650));
    InMux I__4691 (
            .O(N__30655),
            .I(N__30647));
    Odrv12 I__4690 (
            .O(N__30650),
            .I(drone_altitude_0));
    LocalMux I__4689 (
            .O(N__30647),
            .I(drone_altitude_0));
    InMux I__4688 (
            .O(N__30642),
            .I(N__30639));
    LocalMux I__4687 (
            .O(N__30639),
            .I(\dron_frame_decoder_1.drone_altitude_4 ));
    CascadeMux I__4686 (
            .O(N__30636),
            .I(N__30633));
    InMux I__4685 (
            .O(N__30633),
            .I(N__30630));
    LocalMux I__4684 (
            .O(N__30630),
            .I(\uart_pc.data_Auxce_0_5 ));
    InMux I__4683 (
            .O(N__30627),
            .I(N__30624));
    LocalMux I__4682 (
            .O(N__30624),
            .I(\uart_pc.data_Auxce_0_6 ));
    InMux I__4681 (
            .O(N__30621),
            .I(N__30615));
    InMux I__4680 (
            .O(N__30620),
            .I(N__30612));
    InMux I__4679 (
            .O(N__30619),
            .I(N__30609));
    InMux I__4678 (
            .O(N__30618),
            .I(N__30606));
    LocalMux I__4677 (
            .O(N__30615),
            .I(N__30603));
    LocalMux I__4676 (
            .O(N__30612),
            .I(N__30598));
    LocalMux I__4675 (
            .O(N__30609),
            .I(N__30598));
    LocalMux I__4674 (
            .O(N__30606),
            .I(\uart_pc.N_152 ));
    Odrv4 I__4673 (
            .O(N__30603),
            .I(\uart_pc.N_152 ));
    Odrv4 I__4672 (
            .O(N__30598),
            .I(\uart_pc.N_152 ));
    InMux I__4671 (
            .O(N__30591),
            .I(N__30588));
    LocalMux I__4670 (
            .O(N__30588),
            .I(N__30585));
    Odrv4 I__4669 (
            .O(N__30585),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    InMux I__4668 (
            .O(N__30582),
            .I(N__30579));
    LocalMux I__4667 (
            .O(N__30579),
            .I(N__30576));
    Odrv4 I__4666 (
            .O(N__30576),
            .I(\uart_pc.data_Auxce_0_1 ));
    InMux I__4665 (
            .O(N__30573),
            .I(N__30570));
    LocalMux I__4664 (
            .O(N__30570),
            .I(N__30567));
    Odrv4 I__4663 (
            .O(N__30567),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    InMux I__4662 (
            .O(N__30564),
            .I(N__30553));
    InMux I__4661 (
            .O(N__30563),
            .I(N__30546));
    InMux I__4660 (
            .O(N__30562),
            .I(N__30546));
    InMux I__4659 (
            .O(N__30561),
            .I(N__30546));
    InMux I__4658 (
            .O(N__30560),
            .I(N__30535));
    InMux I__4657 (
            .O(N__30559),
            .I(N__30535));
    InMux I__4656 (
            .O(N__30558),
            .I(N__30535));
    InMux I__4655 (
            .O(N__30557),
            .I(N__30535));
    InMux I__4654 (
            .O(N__30556),
            .I(N__30535));
    LocalMux I__4653 (
            .O(N__30553),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__4652 (
            .O(N__30546),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__4651 (
            .O(N__30535),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    InMux I__4650 (
            .O(N__30528),
            .I(N__30505));
    InMux I__4649 (
            .O(N__30527),
            .I(N__30505));
    InMux I__4648 (
            .O(N__30526),
            .I(N__30505));
    InMux I__4647 (
            .O(N__30525),
            .I(N__30505));
    InMux I__4646 (
            .O(N__30524),
            .I(N__30505));
    InMux I__4645 (
            .O(N__30523),
            .I(N__30505));
    InMux I__4644 (
            .O(N__30522),
            .I(N__30494));
    InMux I__4643 (
            .O(N__30521),
            .I(N__30494));
    InMux I__4642 (
            .O(N__30520),
            .I(N__30494));
    InMux I__4641 (
            .O(N__30519),
            .I(N__30494));
    InMux I__4640 (
            .O(N__30518),
            .I(N__30494));
    LocalMux I__4639 (
            .O(N__30505),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__4638 (
            .O(N__30494),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    CascadeMux I__4637 (
            .O(N__30489),
            .I(N__30482));
    CascadeMux I__4636 (
            .O(N__30488),
            .I(N__30478));
    CascadeMux I__4635 (
            .O(N__30487),
            .I(N__30473));
    CascadeMux I__4634 (
            .O(N__30486),
            .I(N__30469));
    InMux I__4633 (
            .O(N__30485),
            .I(N__30457));
    InMux I__4632 (
            .O(N__30482),
            .I(N__30457));
    InMux I__4631 (
            .O(N__30481),
            .I(N__30457));
    InMux I__4630 (
            .O(N__30478),
            .I(N__30457));
    InMux I__4629 (
            .O(N__30477),
            .I(N__30457));
    InMux I__4628 (
            .O(N__30476),
            .I(N__30446));
    InMux I__4627 (
            .O(N__30473),
            .I(N__30446));
    InMux I__4626 (
            .O(N__30472),
            .I(N__30446));
    InMux I__4625 (
            .O(N__30469),
            .I(N__30446));
    InMux I__4624 (
            .O(N__30468),
            .I(N__30446));
    LocalMux I__4623 (
            .O(N__30457),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__4622 (
            .O(N__30446),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    CascadeMux I__4621 (
            .O(N__30441),
            .I(N__30438));
    InMux I__4620 (
            .O(N__30438),
            .I(N__30435));
    LocalMux I__4619 (
            .O(N__30435),
            .I(N__30432));
    Odrv4 I__4618 (
            .O(N__30432),
            .I(\uart_pc.data_Auxce_0_3 ));
    CascadeMux I__4617 (
            .O(N__30429),
            .I(N__30426));
    InMux I__4616 (
            .O(N__30426),
            .I(N__30423));
    LocalMux I__4615 (
            .O(N__30423),
            .I(N__30419));
    InMux I__4614 (
            .O(N__30422),
            .I(N__30416));
    Odrv4 I__4613 (
            .O(N__30419),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    LocalMux I__4612 (
            .O(N__30416),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    InMux I__4611 (
            .O(N__30411),
            .I(N__30408));
    LocalMux I__4610 (
            .O(N__30408),
            .I(N__30404));
    InMux I__4609 (
            .O(N__30407),
            .I(N__30401));
    Odrv4 I__4608 (
            .O(N__30404),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__4607 (
            .O(N__30401),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    CascadeMux I__4606 (
            .O(N__30396),
            .I(N__30393));
    InMux I__4605 (
            .O(N__30393),
            .I(N__30389));
    InMux I__4604 (
            .O(N__30392),
            .I(N__30386));
    LocalMux I__4603 (
            .O(N__30389),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__4602 (
            .O(N__30386),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    InMux I__4601 (
            .O(N__30381),
            .I(N__30357));
    InMux I__4600 (
            .O(N__30380),
            .I(N__30357));
    InMux I__4599 (
            .O(N__30379),
            .I(N__30357));
    InMux I__4598 (
            .O(N__30378),
            .I(N__30357));
    InMux I__4597 (
            .O(N__30377),
            .I(N__30357));
    InMux I__4596 (
            .O(N__30376),
            .I(N__30357));
    InMux I__4595 (
            .O(N__30375),
            .I(N__30357));
    InMux I__4594 (
            .O(N__30374),
            .I(N__30357));
    LocalMux I__4593 (
            .O(N__30357),
            .I(\uart_pc.un1_state_2_0 ));
    IoInMux I__4592 (
            .O(N__30354),
            .I(N__30351));
    LocalMux I__4591 (
            .O(N__30351),
            .I(N__30348));
    Span4Mux_s3_v I__4590 (
            .O(N__30348),
            .I(N__30345));
    Span4Mux_v I__4589 (
            .O(N__30345),
            .I(N__30341));
    InMux I__4588 (
            .O(N__30344),
            .I(N__30330));
    Span4Mux_h I__4587 (
            .O(N__30341),
            .I(N__30323));
    InMux I__4586 (
            .O(N__30340),
            .I(N__30314));
    InMux I__4585 (
            .O(N__30339),
            .I(N__30314));
    InMux I__4584 (
            .O(N__30338),
            .I(N__30314));
    InMux I__4583 (
            .O(N__30337),
            .I(N__30314));
    InMux I__4582 (
            .O(N__30336),
            .I(N__30305));
    InMux I__4581 (
            .O(N__30335),
            .I(N__30305));
    InMux I__4580 (
            .O(N__30334),
            .I(N__30305));
    InMux I__4579 (
            .O(N__30333),
            .I(N__30305));
    LocalMux I__4578 (
            .O(N__30330),
            .I(N__30302));
    InMux I__4577 (
            .O(N__30329),
            .I(N__30295));
    InMux I__4576 (
            .O(N__30328),
            .I(N__30295));
    InMux I__4575 (
            .O(N__30327),
            .I(N__30295));
    InMux I__4574 (
            .O(N__30326),
            .I(N__30292));
    Odrv4 I__4573 (
            .O(N__30323),
            .I(debug_CH2_18A_c));
    LocalMux I__4572 (
            .O(N__30314),
            .I(debug_CH2_18A_c));
    LocalMux I__4571 (
            .O(N__30305),
            .I(debug_CH2_18A_c));
    Odrv4 I__4570 (
            .O(N__30302),
            .I(debug_CH2_18A_c));
    LocalMux I__4569 (
            .O(N__30295),
            .I(debug_CH2_18A_c));
    LocalMux I__4568 (
            .O(N__30292),
            .I(debug_CH2_18A_c));
    CascadeMux I__4567 (
            .O(N__30279),
            .I(N__30275));
    InMux I__4566 (
            .O(N__30278),
            .I(N__30272));
    InMux I__4565 (
            .O(N__30275),
            .I(N__30269));
    LocalMux I__4564 (
            .O(N__30272),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    LocalMux I__4563 (
            .O(N__30269),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    SRMux I__4562 (
            .O(N__30264),
            .I(N__30261));
    LocalMux I__4561 (
            .O(N__30261),
            .I(N__30258));
    Span4Mux_h I__4560 (
            .O(N__30258),
            .I(N__30255));
    Span4Mux_h I__4559 (
            .O(N__30255),
            .I(N__30252));
    Odrv4 I__4558 (
            .O(N__30252),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__4557 (
            .O(N__30249),
            .I(N__30245));
    InMux I__4556 (
            .O(N__30248),
            .I(N__30242));
    LocalMux I__4555 (
            .O(N__30245),
            .I(N__30239));
    LocalMux I__4554 (
            .O(N__30242),
            .I(N__30230));
    Span4Mux_v I__4553 (
            .O(N__30239),
            .I(N__30227));
    InMux I__4552 (
            .O(N__30238),
            .I(N__30224));
    InMux I__4551 (
            .O(N__30237),
            .I(N__30219));
    InMux I__4550 (
            .O(N__30236),
            .I(N__30219));
    InMux I__4549 (
            .O(N__30235),
            .I(N__30212));
    InMux I__4548 (
            .O(N__30234),
            .I(N__30212));
    InMux I__4547 (
            .O(N__30233),
            .I(N__30212));
    Odrv4 I__4546 (
            .O(N__30230),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__4545 (
            .O(N__30227),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__4544 (
            .O(N__30224),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__4543 (
            .O(N__30219),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__4542 (
            .O(N__30212),
            .I(\uart_pc.stateZ0Z_3 ));
    CascadeMux I__4541 (
            .O(N__30201),
            .I(\uart_pc.CO0_cascade_ ));
    CascadeMux I__4540 (
            .O(N__30198),
            .I(N__30194));
    InMux I__4539 (
            .O(N__30197),
            .I(N__30186));
    InMux I__4538 (
            .O(N__30194),
            .I(N__30186));
    InMux I__4537 (
            .O(N__30193),
            .I(N__30186));
    LocalMux I__4536 (
            .O(N__30186),
            .I(N__30183));
    Odrv4 I__4535 (
            .O(N__30183),
            .I(\uart_pc.un1_state_4_0 ));
    InMux I__4534 (
            .O(N__30180),
            .I(N__30174));
    InMux I__4533 (
            .O(N__30179),
            .I(N__30174));
    LocalMux I__4532 (
            .O(N__30174),
            .I(N__30171));
    Odrv4 I__4531 (
            .O(N__30171),
            .I(\uart_pc.un1_state_7_0 ));
    InMux I__4530 (
            .O(N__30168),
            .I(N__30165));
    LocalMux I__4529 (
            .O(N__30165),
            .I(N__30162));
    Odrv12 I__4528 (
            .O(N__30162),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    InMux I__4527 (
            .O(N__30159),
            .I(N__30156));
    LocalMux I__4526 (
            .O(N__30156),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__4525 (
            .O(N__30153),
            .I(\uart_pc.N_145_cascade_ ));
    InMux I__4524 (
            .O(N__30150),
            .I(N__30145));
    InMux I__4523 (
            .O(N__30149),
            .I(N__30141));
    CascadeMux I__4522 (
            .O(N__30148),
            .I(N__30138));
    LocalMux I__4521 (
            .O(N__30145),
            .I(N__30135));
    InMux I__4520 (
            .O(N__30144),
            .I(N__30132));
    LocalMux I__4519 (
            .O(N__30141),
            .I(N__30129));
    InMux I__4518 (
            .O(N__30138),
            .I(N__30126));
    Odrv12 I__4517 (
            .O(N__30135),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__4516 (
            .O(N__30132),
            .I(\uart_pc.stateZ0Z_2 ));
    Odrv4 I__4515 (
            .O(N__30129),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__4514 (
            .O(N__30126),
            .I(\uart_pc.stateZ0Z_2 ));
    InMux I__4513 (
            .O(N__30117),
            .I(N__30114));
    LocalMux I__4512 (
            .O(N__30114),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    CascadeMux I__4511 (
            .O(N__30111),
            .I(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ));
    CascadeMux I__4510 (
            .O(N__30108),
            .I(N__30104));
    CascadeMux I__4509 (
            .O(N__30107),
            .I(N__30101));
    InMux I__4508 (
            .O(N__30104),
            .I(N__30098));
    InMux I__4507 (
            .O(N__30101),
            .I(N__30095));
    LocalMux I__4506 (
            .O(N__30098),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__4505 (
            .O(N__30095),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    CascadeMux I__4504 (
            .O(N__30090),
            .I(N__30086));
    InMux I__4503 (
            .O(N__30089),
            .I(N__30083));
    InMux I__4502 (
            .O(N__30086),
            .I(N__30080));
    LocalMux I__4501 (
            .O(N__30083),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    LocalMux I__4500 (
            .O(N__30080),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    CascadeMux I__4499 (
            .O(N__30075),
            .I(N__30071));
    InMux I__4498 (
            .O(N__30074),
            .I(N__30068));
    InMux I__4497 (
            .O(N__30071),
            .I(N__30065));
    LocalMux I__4496 (
            .O(N__30068),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__4495 (
            .O(N__30065),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    CascadeMux I__4494 (
            .O(N__30060),
            .I(N__30057));
    InMux I__4493 (
            .O(N__30057),
            .I(N__30053));
    InMux I__4492 (
            .O(N__30056),
            .I(N__30050));
    LocalMux I__4491 (
            .O(N__30053),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__4490 (
            .O(N__30050),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    CascadeMux I__4489 (
            .O(N__30045),
            .I(N__30040));
    InMux I__4488 (
            .O(N__30044),
            .I(N__30033));
    InMux I__4487 (
            .O(N__30043),
            .I(N__30033));
    InMux I__4486 (
            .O(N__30040),
            .I(N__30033));
    LocalMux I__4485 (
            .O(N__30033),
            .I(\uart_pc.stateZ0Z_1 ));
    InMux I__4484 (
            .O(N__30030),
            .I(N__30026));
    InMux I__4483 (
            .O(N__30029),
            .I(N__30023));
    LocalMux I__4482 (
            .O(N__30026),
            .I(\uart_pc.N_126_li ));
    LocalMux I__4481 (
            .O(N__30023),
            .I(\uart_pc.N_126_li ));
    CascadeMux I__4480 (
            .O(N__30018),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__4479 (
            .O(N__30015),
            .I(N__30012));
    InMux I__4478 (
            .O(N__30012),
            .I(N__30006));
    InMux I__4477 (
            .O(N__30011),
            .I(N__30006));
    LocalMux I__4476 (
            .O(N__30006),
            .I(\uart_pc.stateZ0Z_0 ));
    CascadeMux I__4475 (
            .O(N__30003),
            .I(N__30000));
    InMux I__4474 (
            .O(N__30000),
            .I(N__29993));
    InMux I__4473 (
            .O(N__29999),
            .I(N__29993));
    CascadeMux I__4472 (
            .O(N__29998),
            .I(N__29988));
    LocalMux I__4471 (
            .O(N__29993),
            .I(N__29985));
    InMux I__4470 (
            .O(N__29992),
            .I(N__29978));
    InMux I__4469 (
            .O(N__29991),
            .I(N__29978));
    InMux I__4468 (
            .O(N__29988),
            .I(N__29978));
    Odrv4 I__4467 (
            .O(N__29985),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__4466 (
            .O(N__29978),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    InMux I__4465 (
            .O(N__29973),
            .I(N__29969));
    InMux I__4464 (
            .O(N__29972),
            .I(N__29962));
    LocalMux I__4463 (
            .O(N__29969),
            .I(N__29959));
    InMux I__4462 (
            .O(N__29968),
            .I(N__29956));
    InMux I__4461 (
            .O(N__29967),
            .I(N__29949));
    InMux I__4460 (
            .O(N__29966),
            .I(N__29949));
    InMux I__4459 (
            .O(N__29965),
            .I(N__29949));
    LocalMux I__4458 (
            .O(N__29962),
            .I(\uart_pc.stateZ0Z_4 ));
    Odrv4 I__4457 (
            .O(N__29959),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__4456 (
            .O(N__29956),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__4455 (
            .O(N__29949),
            .I(\uart_pc.stateZ0Z_4 ));
    CascadeMux I__4454 (
            .O(N__29940),
            .I(\uart_pc.un1_state_4_0_cascade_ ));
    CascadeMux I__4453 (
            .O(N__29937),
            .I(N__29927));
    InMux I__4452 (
            .O(N__29936),
            .I(N__29920));
    InMux I__4451 (
            .O(N__29935),
            .I(N__29920));
    InMux I__4450 (
            .O(N__29934),
            .I(N__29920));
    CascadeMux I__4449 (
            .O(N__29933),
            .I(N__29916));
    CascadeMux I__4448 (
            .O(N__29932),
            .I(N__29913));
    InMux I__4447 (
            .O(N__29931),
            .I(N__29906));
    InMux I__4446 (
            .O(N__29930),
            .I(N__29906));
    InMux I__4445 (
            .O(N__29927),
            .I(N__29906));
    LocalMux I__4444 (
            .O(N__29920),
            .I(N__29903));
    InMux I__4443 (
            .O(N__29919),
            .I(N__29900));
    InMux I__4442 (
            .O(N__29916),
            .I(N__29895));
    InMux I__4441 (
            .O(N__29913),
            .I(N__29895));
    LocalMux I__4440 (
            .O(N__29906),
            .I(N__29892));
    Odrv4 I__4439 (
            .O(N__29903),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__4438 (
            .O(N__29900),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__4437 (
            .O(N__29895),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__4436 (
            .O(N__29892),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    InMux I__4435 (
            .O(N__29883),
            .I(N__29871));
    InMux I__4434 (
            .O(N__29882),
            .I(N__29871));
    InMux I__4433 (
            .O(N__29881),
            .I(N__29868));
    InMux I__4432 (
            .O(N__29880),
            .I(N__29863));
    InMux I__4431 (
            .O(N__29879),
            .I(N__29863));
    InMux I__4430 (
            .O(N__29878),
            .I(N__29856));
    InMux I__4429 (
            .O(N__29877),
            .I(N__29856));
    InMux I__4428 (
            .O(N__29876),
            .I(N__29856));
    LocalMux I__4427 (
            .O(N__29871),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4426 (
            .O(N__29868),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4425 (
            .O(N__29863),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4424 (
            .O(N__29856),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    InMux I__4423 (
            .O(N__29847),
            .I(bfn_8_6_0_));
    InMux I__4422 (
            .O(N__29844),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    InMux I__4421 (
            .O(N__29841),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__4420 (
            .O(N__29838),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    InMux I__4419 (
            .O(N__29835),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    InMux I__4418 (
            .O(N__29832),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__4417 (
            .O(N__29829),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__4416 (
            .O(N__29826),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    SRMux I__4415 (
            .O(N__29823),
            .I(N__29820));
    LocalMux I__4414 (
            .O(N__29820),
            .I(N__29816));
    SRMux I__4413 (
            .O(N__29819),
            .I(N__29813));
    Span4Mux_v I__4412 (
            .O(N__29816),
            .I(N__29808));
    LocalMux I__4411 (
            .O(N__29813),
            .I(N__29808));
    Span4Mux_h I__4410 (
            .O(N__29808),
            .I(N__29805));
    Odrv4 I__4409 (
            .O(N__29805),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    CascadeMux I__4408 (
            .O(N__29802),
            .I(\uart_pc.state_srsts_i_0_2_cascade_ ));
    InMux I__4407 (
            .O(N__29799),
            .I(N__29796));
    LocalMux I__4406 (
            .O(N__29796),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__4405 (
            .O(N__29793),
            .I(N__29790));
    LocalMux I__4404 (
            .O(N__29790),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__4403 (
            .O(N__29787),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__4402 (
            .O(N__29784),
            .I(N__29781));
    LocalMux I__4401 (
            .O(N__29781),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__4400 (
            .O(N__29778),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__4399 (
            .O(N__29775),
            .I(N__29772));
    LocalMux I__4398 (
            .O(N__29772),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__4397 (
            .O(N__29769),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__4396 (
            .O(N__29766),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    InMux I__4395 (
            .O(N__29763),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__4394 (
            .O(N__29760),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    InMux I__4393 (
            .O(N__29757),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    InMux I__4392 (
            .O(N__29754),
            .I(N__29751));
    LocalMux I__4391 (
            .O(N__29751),
            .I(N__29748));
    Odrv12 I__4390 (
            .O(N__29748),
            .I(drone_altitude_i_7));
    CascadeMux I__4389 (
            .O(N__29745),
            .I(N__29742));
    InMux I__4388 (
            .O(N__29742),
            .I(N__29739));
    LocalMux I__4387 (
            .O(N__29739),
            .I(N__29735));
    InMux I__4386 (
            .O(N__29738),
            .I(N__29732));
    Span4Mux_h I__4385 (
            .O(N__29735),
            .I(N__29729));
    LocalMux I__4384 (
            .O(N__29732),
            .I(\pid_alt.drone_altitude_i_0 ));
    Odrv4 I__4383 (
            .O(N__29729),
            .I(\pid_alt.drone_altitude_i_0 ));
    InMux I__4382 (
            .O(N__29724),
            .I(N__29721));
    LocalMux I__4381 (
            .O(N__29721),
            .I(N__29718));
    Odrv12 I__4380 (
            .O(N__29718),
            .I(\pid_alt.error_axbZ0Z_13 ));
    InMux I__4379 (
            .O(N__29715),
            .I(N__29712));
    LocalMux I__4378 (
            .O(N__29712),
            .I(N__29709));
    Odrv12 I__4377 (
            .O(N__29709),
            .I(\pid_alt.error_axbZ0Z_14 ));
    InMux I__4376 (
            .O(N__29706),
            .I(N__29703));
    LocalMux I__4375 (
            .O(N__29703),
            .I(N__29700));
    Odrv12 I__4374 (
            .O(N__29700),
            .I(\pid_alt.error_axbZ0Z_12 ));
    InMux I__4373 (
            .O(N__29697),
            .I(N__29694));
    LocalMux I__4372 (
            .O(N__29694),
            .I(uart_input_drone_c));
    InMux I__4371 (
            .O(N__29691),
            .I(N__29688));
    LocalMux I__4370 (
            .O(N__29688),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    InMux I__4369 (
            .O(N__29685),
            .I(N__29682));
    LocalMux I__4368 (
            .O(N__29682),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    InMux I__4367 (
            .O(N__29679),
            .I(N__29676));
    LocalMux I__4366 (
            .O(N__29676),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    InMux I__4365 (
            .O(N__29673),
            .I(N__29670));
    LocalMux I__4364 (
            .O(N__29670),
            .I(N__29667));
    Span4Mux_v I__4363 (
            .O(N__29667),
            .I(N__29664));
    Span4Mux_h I__4362 (
            .O(N__29664),
            .I(N__29661));
    Odrv4 I__4361 (
            .O(N__29661),
            .I(drone_altitude_15));
    InMux I__4360 (
            .O(N__29658),
            .I(N__29655));
    LocalMux I__4359 (
            .O(N__29655),
            .I(N__29652));
    Span4Mux_v I__4358 (
            .O(N__29652),
            .I(N__29649));
    Span4Mux_h I__4357 (
            .O(N__29649),
            .I(N__29646));
    Odrv4 I__4356 (
            .O(N__29646),
            .I(drone_altitude_i_4));
    InMux I__4355 (
            .O(N__29643),
            .I(N__29640));
    LocalMux I__4354 (
            .O(N__29640),
            .I(N__29637));
    Span4Mux_v I__4353 (
            .O(N__29637),
            .I(N__29634));
    Span4Mux_h I__4352 (
            .O(N__29634),
            .I(N__29631));
    Odrv4 I__4351 (
            .O(N__29631),
            .I(drone_altitude_i_5));
    InMux I__4350 (
            .O(N__29628),
            .I(N__29625));
    LocalMux I__4349 (
            .O(N__29625),
            .I(N__29622));
    Span4Mux_s3_h I__4348 (
            .O(N__29622),
            .I(N__29619));
    Span4Mux_h I__4347 (
            .O(N__29619),
            .I(N__29616));
    Odrv4 I__4346 (
            .O(N__29616),
            .I(drone_altitude_i_6));
    InMux I__4345 (
            .O(N__29613),
            .I(N__29610));
    LocalMux I__4344 (
            .O(N__29610),
            .I(\dron_frame_decoder_1.drone_altitude_9 ));
    InMux I__4343 (
            .O(N__29607),
            .I(N__29604));
    LocalMux I__4342 (
            .O(N__29604),
            .I(N__29601));
    Span4Mux_s3_h I__4341 (
            .O(N__29601),
            .I(N__29598));
    Span4Mux_h I__4340 (
            .O(N__29598),
            .I(N__29595));
    Odrv4 I__4339 (
            .O(N__29595),
            .I(drone_altitude_i_9));
    InMux I__4338 (
            .O(N__29592),
            .I(N__29589));
    LocalMux I__4337 (
            .O(N__29589),
            .I(N__29586));
    Span4Mux_s3_h I__4336 (
            .O(N__29586),
            .I(N__29583));
    Span4Mux_h I__4335 (
            .O(N__29583),
            .I(N__29580));
    Odrv4 I__4334 (
            .O(N__29580),
            .I(drone_altitude_i_8));
    CascadeMux I__4333 (
            .O(N__29577),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ));
    InMux I__4332 (
            .O(N__29574),
            .I(N__29570));
    InMux I__4331 (
            .O(N__29573),
            .I(N__29567));
    LocalMux I__4330 (
            .O(N__29570),
            .I(N__29564));
    LocalMux I__4329 (
            .O(N__29567),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    Odrv4 I__4328 (
            .O(N__29564),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    InMux I__4327 (
            .O(N__29559),
            .I(N__29556));
    LocalMux I__4326 (
            .O(N__29556),
            .I(N__29553));
    Odrv4 I__4325 (
            .O(N__29553),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    InMux I__4324 (
            .O(N__29550),
            .I(N__29544));
    CascadeMux I__4323 (
            .O(N__29549),
            .I(N__29541));
    CascadeMux I__4322 (
            .O(N__29548),
            .I(N__29538));
    CascadeMux I__4321 (
            .O(N__29547),
            .I(N__29535));
    LocalMux I__4320 (
            .O(N__29544),
            .I(N__29532));
    InMux I__4319 (
            .O(N__29541),
            .I(N__29529));
    InMux I__4318 (
            .O(N__29538),
            .I(N__29524));
    InMux I__4317 (
            .O(N__29535),
            .I(N__29524));
    Span4Mux_h I__4316 (
            .O(N__29532),
            .I(N__29521));
    LocalMux I__4315 (
            .O(N__29529),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    LocalMux I__4314 (
            .O(N__29524),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv4 I__4313 (
            .O(N__29521),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    InMux I__4312 (
            .O(N__29514),
            .I(N__29510));
    InMux I__4311 (
            .O(N__29513),
            .I(N__29507));
    LocalMux I__4310 (
            .O(N__29510),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    LocalMux I__4309 (
            .O(N__29507),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    InMux I__4308 (
            .O(N__29502),
            .I(N__29499));
    LocalMux I__4307 (
            .O(N__29499),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__4306 (
            .O(N__29496),
            .I(N__29493));
    LocalMux I__4305 (
            .O(N__29493),
            .I(N__29490));
    Odrv12 I__4304 (
            .O(N__29490),
            .I(\pid_front.O_0_6 ));
    InMux I__4303 (
            .O(N__29487),
            .I(N__29484));
    LocalMux I__4302 (
            .O(N__29484),
            .I(N__29481));
    Span4Mux_h I__4301 (
            .O(N__29481),
            .I(N__29478));
    Odrv4 I__4300 (
            .O(N__29478),
            .I(\pid_front.O_0_4 ));
    InMux I__4299 (
            .O(N__29475),
            .I(N__29472));
    LocalMux I__4298 (
            .O(N__29472),
            .I(N__29469));
    Span4Mux_v I__4297 (
            .O(N__29469),
            .I(N__29466));
    Span4Mux_h I__4296 (
            .O(N__29466),
            .I(N__29463));
    Odrv4 I__4295 (
            .O(N__29463),
            .I(\pid_front.O_0_9 ));
    InMux I__4294 (
            .O(N__29460),
            .I(N__29457));
    LocalMux I__4293 (
            .O(N__29457),
            .I(N__29454));
    Span4Mux_h I__4292 (
            .O(N__29454),
            .I(N__29451));
    Span4Mux_h I__4291 (
            .O(N__29451),
            .I(N__29448));
    Odrv4 I__4290 (
            .O(N__29448),
            .I(\pid_front.O_0_15 ));
    InMux I__4289 (
            .O(N__29445),
            .I(N__29442));
    LocalMux I__4288 (
            .O(N__29442),
            .I(N__29439));
    Odrv12 I__4287 (
            .O(N__29439),
            .I(\dron_frame_decoder_1.drone_altitude_11 ));
    CascadeMux I__4286 (
            .O(N__29436),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ));
    InMux I__4285 (
            .O(N__29433),
            .I(N__29430));
    LocalMux I__4284 (
            .O(N__29430),
            .I(N__29427));
    Span4Mux_v I__4283 (
            .O(N__29427),
            .I(N__29424));
    Span4Mux_h I__4282 (
            .O(N__29424),
            .I(N__29420));
    InMux I__4281 (
            .O(N__29423),
            .I(N__29417));
    Span4Mux_h I__4280 (
            .O(N__29420),
            .I(N__29414));
    LocalMux I__4279 (
            .O(N__29417),
            .I(N__29411));
    Span4Mux_h I__4278 (
            .O(N__29414),
            .I(N__29407));
    Span4Mux_v I__4277 (
            .O(N__29411),
            .I(N__29404));
    InMux I__4276 (
            .O(N__29410),
            .I(N__29401));
    Span4Mux_h I__4275 (
            .O(N__29407),
            .I(N__29396));
    Span4Mux_h I__4274 (
            .O(N__29404),
            .I(N__29396));
    LocalMux I__4273 (
            .O(N__29401),
            .I(xy_kp_4));
    Odrv4 I__4272 (
            .O(N__29396),
            .I(xy_kp_4));
    InMux I__4271 (
            .O(N__29391),
            .I(N__29388));
    LocalMux I__4270 (
            .O(N__29388),
            .I(N__29384));
    CascadeMux I__4269 (
            .O(N__29387),
            .I(N__29380));
    Span4Mux_v I__4268 (
            .O(N__29384),
            .I(N__29376));
    InMux I__4267 (
            .O(N__29383),
            .I(N__29369));
    InMux I__4266 (
            .O(N__29380),
            .I(N__29369));
    InMux I__4265 (
            .O(N__29379),
            .I(N__29369));
    Odrv4 I__4264 (
            .O(N__29376),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__4263 (
            .O(N__29369),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    InMux I__4262 (
            .O(N__29364),
            .I(N__29358));
    InMux I__4261 (
            .O(N__29363),
            .I(N__29358));
    LocalMux I__4260 (
            .O(N__29358),
            .I(N__29355));
    Odrv4 I__4259 (
            .O(N__29355),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    InMux I__4258 (
            .O(N__29352),
            .I(N__29348));
    InMux I__4257 (
            .O(N__29351),
            .I(N__29344));
    LocalMux I__4256 (
            .O(N__29348),
            .I(N__29341));
    CascadeMux I__4255 (
            .O(N__29347),
            .I(N__29338));
    LocalMux I__4254 (
            .O(N__29344),
            .I(N__29335));
    Span4Mux_h I__4253 (
            .O(N__29341),
            .I(N__29332));
    InMux I__4252 (
            .O(N__29338),
            .I(N__29329));
    Span12Mux_s11_v I__4251 (
            .O(N__29335),
            .I(N__29326));
    Span4Mux_v I__4250 (
            .O(N__29332),
            .I(N__29323));
    LocalMux I__4249 (
            .O(N__29329),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv12 I__4248 (
            .O(N__29326),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv4 I__4247 (
            .O(N__29323),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    InMux I__4246 (
            .O(N__29316),
            .I(N__29313));
    LocalMux I__4245 (
            .O(N__29313),
            .I(N__29310));
    Span4Mux_v I__4244 (
            .O(N__29310),
            .I(N__29307));
    Sp12to4 I__4243 (
            .O(N__29307),
            .I(N__29303));
    InMux I__4242 (
            .O(N__29306),
            .I(N__29300));
    Span12Mux_s7_h I__4241 (
            .O(N__29303),
            .I(N__29297));
    LocalMux I__4240 (
            .O(N__29300),
            .I(alt_kp_4));
    Odrv12 I__4239 (
            .O(N__29297),
            .I(alt_kp_4));
    InMux I__4238 (
            .O(N__29292),
            .I(N__29289));
    LocalMux I__4237 (
            .O(N__29289),
            .I(N__29283));
    InMux I__4236 (
            .O(N__29288),
            .I(N__29276));
    InMux I__4235 (
            .O(N__29287),
            .I(N__29276));
    InMux I__4234 (
            .O(N__29286),
            .I(N__29276));
    Odrv4 I__4233 (
            .O(N__29283),
            .I(\uart_pc.data_rdyc_1 ));
    LocalMux I__4232 (
            .O(N__29276),
            .I(\uart_pc.data_rdyc_1 ));
    CascadeMux I__4231 (
            .O(N__29271),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ));
    InMux I__4230 (
            .O(N__29268),
            .I(N__29262));
    InMux I__4229 (
            .O(N__29267),
            .I(N__29262));
    LocalMux I__4228 (
            .O(N__29262),
            .I(N__29259));
    Odrv4 I__4227 (
            .O(N__29259),
            .I(\Commands_frame_decoder.N_378 ));
    InMux I__4226 (
            .O(N__29256),
            .I(N__29243));
    InMux I__4225 (
            .O(N__29255),
            .I(N__29243));
    InMux I__4224 (
            .O(N__29254),
            .I(N__29243));
    InMux I__4223 (
            .O(N__29253),
            .I(N__29234));
    InMux I__4222 (
            .O(N__29252),
            .I(N__29234));
    InMux I__4221 (
            .O(N__29251),
            .I(N__29234));
    InMux I__4220 (
            .O(N__29250),
            .I(N__29234));
    LocalMux I__4219 (
            .O(N__29243),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__4218 (
            .O(N__29234),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    CascadeMux I__4217 (
            .O(N__29229),
            .I(N__29224));
    CascadeMux I__4216 (
            .O(N__29228),
            .I(N__29219));
    InMux I__4215 (
            .O(N__29227),
            .I(N__29211));
    InMux I__4214 (
            .O(N__29224),
            .I(N__29211));
    InMux I__4213 (
            .O(N__29223),
            .I(N__29211));
    InMux I__4212 (
            .O(N__29222),
            .I(N__29204));
    InMux I__4211 (
            .O(N__29219),
            .I(N__29204));
    InMux I__4210 (
            .O(N__29218),
            .I(N__29204));
    LocalMux I__4209 (
            .O(N__29211),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__4208 (
            .O(N__29204),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    CascadeMux I__4207 (
            .O(N__29199),
            .I(N__29195));
    CascadeMux I__4206 (
            .O(N__29198),
            .I(N__29192));
    InMux I__4205 (
            .O(N__29195),
            .I(N__29189));
    InMux I__4204 (
            .O(N__29192),
            .I(N__29186));
    LocalMux I__4203 (
            .O(N__29189),
            .I(N__29183));
    LocalMux I__4202 (
            .O(N__29186),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    Odrv4 I__4201 (
            .O(N__29183),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    InMux I__4200 (
            .O(N__29178),
            .I(N__29175));
    LocalMux I__4199 (
            .O(N__29175),
            .I(N__29172));
    Span4Mux_h I__4198 (
            .O(N__29172),
            .I(N__29169));
    Odrv4 I__4197 (
            .O(N__29169),
            .I(\Commands_frame_decoder.state_ns_0_i_1_1 ));
    InMux I__4196 (
            .O(N__29166),
            .I(N__29163));
    LocalMux I__4195 (
            .O(N__29163),
            .I(N__29160));
    Span4Mux_v I__4194 (
            .O(N__29160),
            .I(N__29156));
    InMux I__4193 (
            .O(N__29159),
            .I(N__29153));
    Span4Mux_v I__4192 (
            .O(N__29156),
            .I(N__29150));
    LocalMux I__4191 (
            .O(N__29153),
            .I(N__29147));
    Span4Mux_h I__4190 (
            .O(N__29150),
            .I(N__29144));
    Span4Mux_h I__4189 (
            .O(N__29147),
            .I(N__29141));
    Odrv4 I__4188 (
            .O(N__29144),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ));
    Odrv4 I__4187 (
            .O(N__29141),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ));
    InMux I__4186 (
            .O(N__29136),
            .I(N__29131));
    InMux I__4185 (
            .O(N__29135),
            .I(N__29126));
    InMux I__4184 (
            .O(N__29134),
            .I(N__29126));
    LocalMux I__4183 (
            .O(N__29131),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__4182 (
            .O(N__29126),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    CascadeMux I__4181 (
            .O(N__29121),
            .I(\uart_pc.N_126_li_cascade_ ));
    CascadeMux I__4180 (
            .O(N__29118),
            .I(N__29114));
    CascadeMux I__4179 (
            .O(N__29117),
            .I(N__29111));
    InMux I__4178 (
            .O(N__29114),
            .I(N__29101));
    InMux I__4177 (
            .O(N__29111),
            .I(N__29101));
    InMux I__4176 (
            .O(N__29110),
            .I(N__29101));
    InMux I__4175 (
            .O(N__29109),
            .I(N__29096));
    InMux I__4174 (
            .O(N__29108),
            .I(N__29096));
    LocalMux I__4173 (
            .O(N__29101),
            .I(\uart_pc.N_143 ));
    LocalMux I__4172 (
            .O(N__29096),
            .I(\uart_pc.N_143 ));
    CascadeMux I__4171 (
            .O(N__29091),
            .I(\uart_pc.N_143_cascade_ ));
    CascadeMux I__4170 (
            .O(N__29088),
            .I(N__29082));
    InMux I__4169 (
            .O(N__29087),
            .I(N__29079));
    InMux I__4168 (
            .O(N__29086),
            .I(N__29072));
    InMux I__4167 (
            .O(N__29085),
            .I(N__29072));
    InMux I__4166 (
            .O(N__29082),
            .I(N__29072));
    LocalMux I__4165 (
            .O(N__29079),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__4164 (
            .O(N__29072),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    CascadeMux I__4163 (
            .O(N__29067),
            .I(N__29064));
    InMux I__4162 (
            .O(N__29064),
            .I(N__29061));
    LocalMux I__4161 (
            .O(N__29061),
            .I(N__29058));
    Span4Mux_h I__4160 (
            .O(N__29058),
            .I(N__29055));
    Odrv4 I__4159 (
            .O(N__29055),
            .I(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ));
    CascadeMux I__4158 (
            .O(N__29052),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ));
    InMux I__4157 (
            .O(N__29049),
            .I(N__29046));
    LocalMux I__4156 (
            .O(N__29046),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4 ));
    InMux I__4155 (
            .O(N__29043),
            .I(N__29040));
    LocalMux I__4154 (
            .O(N__29040),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1 ));
    InMux I__4153 (
            .O(N__29037),
            .I(N__29031));
    InMux I__4152 (
            .O(N__29036),
            .I(N__29031));
    LocalMux I__4151 (
            .O(N__29031),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    InMux I__4150 (
            .O(N__29028),
            .I(N__29025));
    LocalMux I__4149 (
            .O(N__29025),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    CascadeMux I__4148 (
            .O(N__29022),
            .I(\uart_pc.N_144_1_cascade_ ));
    CascadeMux I__4147 (
            .O(N__29019),
            .I(N__29016));
    InMux I__4146 (
            .O(N__29016),
            .I(N__29013));
    LocalMux I__4145 (
            .O(N__29013),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    InMux I__4144 (
            .O(N__29010),
            .I(N__29007));
    LocalMux I__4143 (
            .O(N__29007),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    InMux I__4142 (
            .O(N__29004),
            .I(N__28998));
    InMux I__4141 (
            .O(N__29003),
            .I(N__28998));
    LocalMux I__4140 (
            .O(N__28998),
            .I(N__28995));
    Odrv4 I__4139 (
            .O(N__28995),
            .I(\pid_alt.N_44 ));
    InMux I__4138 (
            .O(N__28992),
            .I(N__28988));
    InMux I__4137 (
            .O(N__28991),
            .I(N__28985));
    LocalMux I__4136 (
            .O(N__28988),
            .I(N__28982));
    LocalMux I__4135 (
            .O(N__28985),
            .I(N__28979));
    Span4Mux_v I__4134 (
            .O(N__28982),
            .I(N__28976));
    Span4Mux_h I__4133 (
            .O(N__28979),
            .I(N__28973));
    Odrv4 I__4132 (
            .O(N__28976),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    Odrv4 I__4131 (
            .O(N__28973),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    InMux I__4130 (
            .O(N__28968),
            .I(N__28962));
    InMux I__4129 (
            .O(N__28967),
            .I(N__28962));
    LocalMux I__4128 (
            .O(N__28962),
            .I(N__28956));
    InMux I__4127 (
            .O(N__28961),
            .I(N__28953));
    InMux I__4126 (
            .O(N__28960),
            .I(N__28950));
    InMux I__4125 (
            .O(N__28959),
            .I(N__28947));
    Span4Mux_v I__4124 (
            .O(N__28956),
            .I(N__28942));
    LocalMux I__4123 (
            .O(N__28953),
            .I(N__28942));
    LocalMux I__4122 (
            .O(N__28950),
            .I(N__28938));
    LocalMux I__4121 (
            .O(N__28947),
            .I(N__28935));
    Span4Mux_v I__4120 (
            .O(N__28942),
            .I(N__28932));
    InMux I__4119 (
            .O(N__28941),
            .I(N__28929));
    Span4Mux_h I__4118 (
            .O(N__28938),
            .I(N__28926));
    Span4Mux_h I__4117 (
            .O(N__28935),
            .I(N__28923));
    Span4Mux_h I__4116 (
            .O(N__28932),
            .I(N__28918));
    LocalMux I__4115 (
            .O(N__28929),
            .I(N__28918));
    Odrv4 I__4114 (
            .O(N__28926),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__4113 (
            .O(N__28923),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__4112 (
            .O(N__28918),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    CascadeMux I__4111 (
            .O(N__28911),
            .I(N__28907));
    CascadeMux I__4110 (
            .O(N__28910),
            .I(N__28896));
    InMux I__4109 (
            .O(N__28907),
            .I(N__28891));
    InMux I__4108 (
            .O(N__28906),
            .I(N__28891));
    InMux I__4107 (
            .O(N__28905),
            .I(N__28888));
    InMux I__4106 (
            .O(N__28904),
            .I(N__28881));
    InMux I__4105 (
            .O(N__28903),
            .I(N__28881));
    InMux I__4104 (
            .O(N__28902),
            .I(N__28881));
    InMux I__4103 (
            .O(N__28901),
            .I(N__28876));
    InMux I__4102 (
            .O(N__28900),
            .I(N__28876));
    InMux I__4101 (
            .O(N__28899),
            .I(N__28873));
    InMux I__4100 (
            .O(N__28896),
            .I(N__28870));
    LocalMux I__4099 (
            .O(N__28891),
            .I(N__28867));
    LocalMux I__4098 (
            .O(N__28888),
            .I(N__28862));
    LocalMux I__4097 (
            .O(N__28881),
            .I(N__28862));
    LocalMux I__4096 (
            .O(N__28876),
            .I(N__28855));
    LocalMux I__4095 (
            .O(N__28873),
            .I(N__28855));
    LocalMux I__4094 (
            .O(N__28870),
            .I(N__28855));
    Span4Mux_h I__4093 (
            .O(N__28867),
            .I(N__28848));
    Span4Mux_v I__4092 (
            .O(N__28862),
            .I(N__28848));
    Span4Mux_v I__4091 (
            .O(N__28855),
            .I(N__28848));
    Sp12to4 I__4090 (
            .O(N__28848),
            .I(N__28845));
    Span12Mux_s3_h I__4089 (
            .O(N__28845),
            .I(N__28842));
    Odrv12 I__4088 (
            .O(N__28842),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    CascadeMux I__4087 (
            .O(N__28839),
            .I(N__28829));
    CascadeMux I__4086 (
            .O(N__28838),
            .I(N__28826));
    InMux I__4085 (
            .O(N__28837),
            .I(N__28815));
    InMux I__4084 (
            .O(N__28836),
            .I(N__28815));
    InMux I__4083 (
            .O(N__28835),
            .I(N__28815));
    InMux I__4082 (
            .O(N__28834),
            .I(N__28815));
    InMux I__4081 (
            .O(N__28833),
            .I(N__28812));
    InMux I__4080 (
            .O(N__28832),
            .I(N__28809));
    InMux I__4079 (
            .O(N__28829),
            .I(N__28799));
    InMux I__4078 (
            .O(N__28826),
            .I(N__28799));
    InMux I__4077 (
            .O(N__28825),
            .I(N__28799));
    InMux I__4076 (
            .O(N__28824),
            .I(N__28799));
    LocalMux I__4075 (
            .O(N__28815),
            .I(N__28794));
    LocalMux I__4074 (
            .O(N__28812),
            .I(N__28794));
    LocalMux I__4073 (
            .O(N__28809),
            .I(N__28791));
    InMux I__4072 (
            .O(N__28808),
            .I(N__28788));
    LocalMux I__4071 (
            .O(N__28799),
            .I(\pid_alt.N_305 ));
    Odrv4 I__4070 (
            .O(N__28794),
            .I(\pid_alt.N_305 ));
    Odrv12 I__4069 (
            .O(N__28791),
            .I(\pid_alt.N_305 ));
    LocalMux I__4068 (
            .O(N__28788),
            .I(\pid_alt.N_305 ));
    CascadeMux I__4067 (
            .O(N__28779),
            .I(N__28775));
    InMux I__4066 (
            .O(N__28778),
            .I(N__28771));
    InMux I__4065 (
            .O(N__28775),
            .I(N__28768));
    InMux I__4064 (
            .O(N__28774),
            .I(N__28765));
    LocalMux I__4063 (
            .O(N__28771),
            .I(N__28761));
    LocalMux I__4062 (
            .O(N__28768),
            .I(N__28758));
    LocalMux I__4061 (
            .O(N__28765),
            .I(N__28755));
    InMux I__4060 (
            .O(N__28764),
            .I(N__28752));
    Span4Mux_v I__4059 (
            .O(N__28761),
            .I(N__28749));
    Span4Mux_h I__4058 (
            .O(N__28758),
            .I(N__28746));
    Span4Mux_h I__4057 (
            .O(N__28755),
            .I(N__28743));
    LocalMux I__4056 (
            .O(N__28752),
            .I(N__28740));
    Odrv4 I__4055 (
            .O(N__28749),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv4 I__4054 (
            .O(N__28746),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv4 I__4053 (
            .O(N__28743),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv12 I__4052 (
            .O(N__28740),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    CEMux I__4051 (
            .O(N__28731),
            .I(N__28727));
    CEMux I__4050 (
            .O(N__28730),
            .I(N__28724));
    LocalMux I__4049 (
            .O(N__28727),
            .I(N__28719));
    LocalMux I__4048 (
            .O(N__28724),
            .I(N__28719));
    Odrv4 I__4047 (
            .O(N__28719),
            .I(\pid_alt.N_72_i_1 ));
    SRMux I__4046 (
            .O(N__28716),
            .I(N__28712));
    SRMux I__4045 (
            .O(N__28715),
            .I(N__28709));
    LocalMux I__4044 (
            .O(N__28712),
            .I(N__28703));
    LocalMux I__4043 (
            .O(N__28709),
            .I(N__28703));
    SRMux I__4042 (
            .O(N__28708),
            .I(N__28700));
    Sp12to4 I__4041 (
            .O(N__28703),
            .I(N__28694));
    LocalMux I__4040 (
            .O(N__28700),
            .I(N__28694));
    InMux I__4039 (
            .O(N__28699),
            .I(N__28691));
    Odrv12 I__4038 (
            .O(N__28694),
            .I(\pid_alt.un1_reset_0_i ));
    LocalMux I__4037 (
            .O(N__28691),
            .I(\pid_alt.un1_reset_0_i ));
    InMux I__4036 (
            .O(N__28686),
            .I(N__28682));
    InMux I__4035 (
            .O(N__28685),
            .I(N__28679));
    LocalMux I__4034 (
            .O(N__28682),
            .I(N__28674));
    LocalMux I__4033 (
            .O(N__28679),
            .I(N__28674));
    Span4Mux_v I__4032 (
            .O(N__28674),
            .I(N__28671));
    Span4Mux_v I__4031 (
            .O(N__28671),
            .I(N__28668));
    Odrv4 I__4030 (
            .O(N__28668),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    InMux I__4029 (
            .O(N__28665),
            .I(N__28662));
    LocalMux I__4028 (
            .O(N__28662),
            .I(N__28658));
    InMux I__4027 (
            .O(N__28661),
            .I(N__28655));
    Span4Mux_v I__4026 (
            .O(N__28658),
            .I(N__28650));
    LocalMux I__4025 (
            .O(N__28655),
            .I(N__28650));
    Span4Mux_h I__4024 (
            .O(N__28650),
            .I(N__28647));
    Odrv4 I__4023 (
            .O(N__28647),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    InMux I__4022 (
            .O(N__28644),
            .I(N__28641));
    LocalMux I__4021 (
            .O(N__28641),
            .I(N__28637));
    InMux I__4020 (
            .O(N__28640),
            .I(N__28634));
    Span4Mux_v I__4019 (
            .O(N__28637),
            .I(N__28628));
    LocalMux I__4018 (
            .O(N__28634),
            .I(N__28628));
    InMux I__4017 (
            .O(N__28633),
            .I(N__28625));
    Span4Mux_h I__4016 (
            .O(N__28628),
            .I(N__28622));
    LocalMux I__4015 (
            .O(N__28625),
            .I(N__28619));
    Span4Mux_v I__4014 (
            .O(N__28622),
            .I(N__28616));
    Span4Mux_h I__4013 (
            .O(N__28619),
            .I(N__28611));
    Span4Mux_v I__4012 (
            .O(N__28616),
            .I(N__28611));
    Span4Mux_v I__4011 (
            .O(N__28611),
            .I(N__28608));
    Odrv4 I__4010 (
            .O(N__28608),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    InMux I__4009 (
            .O(N__28605),
            .I(N__28601));
    InMux I__4008 (
            .O(N__28604),
            .I(N__28598));
    LocalMux I__4007 (
            .O(N__28601),
            .I(N__28595));
    LocalMux I__4006 (
            .O(N__28598),
            .I(N__28592));
    Span4Mux_h I__4005 (
            .O(N__28595),
            .I(N__28589));
    Span4Mux_h I__4004 (
            .O(N__28592),
            .I(N__28586));
    Odrv4 I__4003 (
            .O(N__28589),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ));
    Odrv4 I__4002 (
            .O(N__28586),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ));
    InMux I__4001 (
            .O(N__28581),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__4000 (
            .O(N__28578),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__3999 (
            .O(N__28575),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    CascadeMux I__3998 (
            .O(N__28572),
            .I(\pid_alt.N_90_cascade_ ));
    InMux I__3997 (
            .O(N__28569),
            .I(N__28563));
    InMux I__3996 (
            .O(N__28568),
            .I(N__28563));
    LocalMux I__3995 (
            .O(N__28563),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ));
    CascadeMux I__3994 (
            .O(N__28560),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ));
    InMux I__3993 (
            .O(N__28557),
            .I(N__28553));
    InMux I__3992 (
            .O(N__28556),
            .I(N__28550));
    LocalMux I__3991 (
            .O(N__28553),
            .I(\pid_alt.N_43 ));
    LocalMux I__3990 (
            .O(N__28550),
            .I(\pid_alt.N_43 ));
    InMux I__3989 (
            .O(N__28545),
            .I(N__28542));
    LocalMux I__3988 (
            .O(N__28542),
            .I(N__28539));
    Odrv12 I__3987 (
            .O(N__28539),
            .I(\pid_alt.N_48 ));
    InMux I__3986 (
            .O(N__28536),
            .I(N__28533));
    LocalMux I__3985 (
            .O(N__28533),
            .I(N__28530));
    Odrv12 I__3984 (
            .O(N__28530),
            .I(\pid_alt.pid_preregZ0Z_15 ));
    InMux I__3983 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__3982 (
            .O(N__28524),
            .I(N__28521));
    Span4Mux_v I__3981 (
            .O(N__28521),
            .I(N__28518));
    Odrv4 I__3980 (
            .O(N__28518),
            .I(\pid_alt.pid_preregZ0Z_23 ));
    CascadeMux I__3979 (
            .O(N__28515),
            .I(N__28512));
    InMux I__3978 (
            .O(N__28512),
            .I(N__28509));
    LocalMux I__3977 (
            .O(N__28509),
            .I(N__28506));
    Span4Mux_h I__3976 (
            .O(N__28506),
            .I(N__28503));
    Odrv4 I__3975 (
            .O(N__28503),
            .I(\pid_alt.pid_preregZ0Z_21 ));
    InMux I__3974 (
            .O(N__28500),
            .I(N__28497));
    LocalMux I__3973 (
            .O(N__28497),
            .I(N__28494));
    Odrv4 I__3972 (
            .O(N__28494),
            .I(\pid_alt.pid_preregZ0Z_18 ));
    InMux I__3971 (
            .O(N__28491),
            .I(N__28488));
    LocalMux I__3970 (
            .O(N__28488),
            .I(N__28485));
    Span4Mux_h I__3969 (
            .O(N__28485),
            .I(N__28482));
    Odrv4 I__3968 (
            .O(N__28482),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    InMux I__3967 (
            .O(N__28479),
            .I(N__28476));
    LocalMux I__3966 (
            .O(N__28476),
            .I(N__28473));
    Odrv4 I__3965 (
            .O(N__28473),
            .I(\pid_alt.pid_preregZ0Z_20 ));
    CascadeMux I__3964 (
            .O(N__28470),
            .I(N__28467));
    InMux I__3963 (
            .O(N__28467),
            .I(N__28464));
    LocalMux I__3962 (
            .O(N__28464),
            .I(N__28461));
    Odrv4 I__3961 (
            .O(N__28461),
            .I(\pid_alt.pid_preregZ0Z_17 ));
    InMux I__3960 (
            .O(N__28458),
            .I(N__28455));
    LocalMux I__3959 (
            .O(N__28455),
            .I(N__28452));
    Odrv4 I__3958 (
            .O(N__28452),
            .I(\pid_alt.pid_preregZ0Z_19 ));
    InMux I__3957 (
            .O(N__28449),
            .I(N__28446));
    LocalMux I__3956 (
            .O(N__28446),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ));
    InMux I__3955 (
            .O(N__28443),
            .I(N__28440));
    LocalMux I__3954 (
            .O(N__28440),
            .I(N__28437));
    Span4Mux_h I__3953 (
            .O(N__28437),
            .I(N__28434));
    Odrv4 I__3952 (
            .O(N__28434),
            .I(\pid_alt.pid_preregZ0Z_14 ));
    CascadeMux I__3951 (
            .O(N__28431),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ));
    InMux I__3950 (
            .O(N__28428),
            .I(N__28425));
    LocalMux I__3949 (
            .O(N__28425),
            .I(N__28422));
    Odrv4 I__3948 (
            .O(N__28422),
            .I(\pid_alt.pid_preregZ0Z_16 ));
    InMux I__3947 (
            .O(N__28419),
            .I(N__28416));
    LocalMux I__3946 (
            .O(N__28416),
            .I(N__28411));
    InMux I__3945 (
            .O(N__28415),
            .I(N__28408));
    InMux I__3944 (
            .O(N__28414),
            .I(N__28405));
    Odrv4 I__3943 (
            .O(N__28411),
            .I(\pid_alt.N_90 ));
    LocalMux I__3942 (
            .O(N__28408),
            .I(\pid_alt.N_90 ));
    LocalMux I__3941 (
            .O(N__28405),
            .I(\pid_alt.N_90 ));
    CascadeMux I__3940 (
            .O(N__28398),
            .I(\pid_alt.N_305_cascade_ ));
    CascadeMux I__3939 (
            .O(N__28395),
            .I(\pid_alt.source_pid_9_0_0_4_cascade_ ));
    InMux I__3938 (
            .O(N__28392),
            .I(N__28383));
    InMux I__3937 (
            .O(N__28391),
            .I(N__28383));
    InMux I__3936 (
            .O(N__28390),
            .I(N__28378));
    InMux I__3935 (
            .O(N__28389),
            .I(N__28378));
    InMux I__3934 (
            .O(N__28388),
            .I(N__28375));
    LocalMux I__3933 (
            .O(N__28383),
            .I(N__28372));
    LocalMux I__3932 (
            .O(N__28378),
            .I(N__28369));
    LocalMux I__3931 (
            .O(N__28375),
            .I(N__28366));
    Span4Mux_v I__3930 (
            .O(N__28372),
            .I(N__28361));
    Span4Mux_v I__3929 (
            .O(N__28369),
            .I(N__28361));
    Odrv4 I__3928 (
            .O(N__28366),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    Odrv4 I__3927 (
            .O(N__28361),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    CascadeMux I__3926 (
            .O(N__28356),
            .I(\pid_alt.N_44_cascade_ ));
    CascadeMux I__3925 (
            .O(N__28353),
            .I(N__28350));
    InMux I__3924 (
            .O(N__28350),
            .I(N__28341));
    InMux I__3923 (
            .O(N__28349),
            .I(N__28341));
    InMux I__3922 (
            .O(N__28348),
            .I(N__28341));
    LocalMux I__3921 (
            .O(N__28341),
            .I(\pid_alt.N_46 ));
    InMux I__3920 (
            .O(N__28338),
            .I(N__28332));
    InMux I__3919 (
            .O(N__28337),
            .I(N__28332));
    LocalMux I__3918 (
            .O(N__28332),
            .I(N__28329));
    Odrv4 I__3917 (
            .O(N__28329),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    CascadeMux I__3916 (
            .O(N__28326),
            .I(\pid_alt.N_46_cascade_ ));
    CascadeMux I__3915 (
            .O(N__28323),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ));
    InMux I__3914 (
            .O(N__28320),
            .I(N__28317));
    LocalMux I__3913 (
            .O(N__28317),
            .I(N__28314));
    Odrv4 I__3912 (
            .O(N__28314),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ));
    InMux I__3911 (
            .O(N__28311),
            .I(N__28308));
    LocalMux I__3910 (
            .O(N__28308),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ));
    InMux I__3909 (
            .O(N__28305),
            .I(N__28302));
    LocalMux I__3908 (
            .O(N__28302),
            .I(N__28297));
    InMux I__3907 (
            .O(N__28301),
            .I(N__28292));
    InMux I__3906 (
            .O(N__28300),
            .I(N__28292));
    Span4Mux_h I__3905 (
            .O(N__28297),
            .I(N__28289));
    LocalMux I__3904 (
            .O(N__28292),
            .I(N__28286));
    Odrv4 I__3903 (
            .O(N__28289),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    Odrv4 I__3902 (
            .O(N__28286),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    InMux I__3901 (
            .O(N__28281),
            .I(N__28277));
    CascadeMux I__3900 (
            .O(N__28280),
            .I(N__28274));
    LocalMux I__3899 (
            .O(N__28277),
            .I(N__28270));
    InMux I__3898 (
            .O(N__28274),
            .I(N__28265));
    InMux I__3897 (
            .O(N__28273),
            .I(N__28265));
    Span4Mux_v I__3896 (
            .O(N__28270),
            .I(N__28260));
    LocalMux I__3895 (
            .O(N__28265),
            .I(N__28260));
    Odrv4 I__3894 (
            .O(N__28260),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    InMux I__3893 (
            .O(N__28257),
            .I(N__28253));
    CascadeMux I__3892 (
            .O(N__28256),
            .I(N__28249));
    LocalMux I__3891 (
            .O(N__28253),
            .I(N__28246));
    InMux I__3890 (
            .O(N__28252),
            .I(N__28243));
    InMux I__3889 (
            .O(N__28249),
            .I(N__28240));
    Span4Mux_v I__3888 (
            .O(N__28246),
            .I(N__28233));
    LocalMux I__3887 (
            .O(N__28243),
            .I(N__28233));
    LocalMux I__3886 (
            .O(N__28240),
            .I(N__28233));
    Odrv4 I__3885 (
            .O(N__28233),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    InMux I__3884 (
            .O(N__28230),
            .I(N__28227));
    LocalMux I__3883 (
            .O(N__28227),
            .I(N__28222));
    InMux I__3882 (
            .O(N__28226),
            .I(N__28217));
    InMux I__3881 (
            .O(N__28225),
            .I(N__28217));
    Span4Mux_h I__3880 (
            .O(N__28222),
            .I(N__28214));
    LocalMux I__3879 (
            .O(N__28217),
            .I(N__28211));
    Odrv4 I__3878 (
            .O(N__28214),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    Odrv12 I__3877 (
            .O(N__28211),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    InMux I__3876 (
            .O(N__28206),
            .I(N__28202));
    CascadeMux I__3875 (
            .O(N__28205),
            .I(N__28199));
    LocalMux I__3874 (
            .O(N__28202),
            .I(N__28195));
    InMux I__3873 (
            .O(N__28199),
            .I(N__28190));
    InMux I__3872 (
            .O(N__28198),
            .I(N__28190));
    Span4Mux_v I__3871 (
            .O(N__28195),
            .I(N__28185));
    LocalMux I__3870 (
            .O(N__28190),
            .I(N__28185));
    Odrv4 I__3869 (
            .O(N__28185),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    CascadeMux I__3868 (
            .O(N__28182),
            .I(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ));
    InMux I__3867 (
            .O(N__28179),
            .I(N__28174));
    InMux I__3866 (
            .O(N__28178),
            .I(N__28169));
    InMux I__3865 (
            .O(N__28177),
            .I(N__28169));
    LocalMux I__3864 (
            .O(N__28174),
            .I(N__28166));
    LocalMux I__3863 (
            .O(N__28169),
            .I(N__28163));
    Span4Mux_h I__3862 (
            .O(N__28166),
            .I(N__28160));
    Span4Mux_h I__3861 (
            .O(N__28163),
            .I(N__28157));
    Odrv4 I__3860 (
            .O(N__28160),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    Odrv4 I__3859 (
            .O(N__28157),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    InMux I__3858 (
            .O(N__28152),
            .I(N__28137));
    InMux I__3857 (
            .O(N__28151),
            .I(N__28137));
    InMux I__3856 (
            .O(N__28150),
            .I(N__28137));
    InMux I__3855 (
            .O(N__28149),
            .I(N__28137));
    InMux I__3854 (
            .O(N__28148),
            .I(N__28137));
    LocalMux I__3853 (
            .O(N__28137),
            .I(\pid_alt.source_pid_9_0_tz_6 ));
    CascadeMux I__3852 (
            .O(N__28134),
            .I(N__28131));
    InMux I__3851 (
            .O(N__28131),
            .I(N__28125));
    InMux I__3850 (
            .O(N__28130),
            .I(N__28125));
    LocalMux I__3849 (
            .O(N__28125),
            .I(N__28122));
    Odrv4 I__3848 (
            .O(N__28122),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    CascadeMux I__3847 (
            .O(N__28119),
            .I(N__28115));
    InMux I__3846 (
            .O(N__28118),
            .I(N__28110));
    InMux I__3845 (
            .O(N__28115),
            .I(N__28110));
    LocalMux I__3844 (
            .O(N__28110),
            .I(N__28107));
    Odrv4 I__3843 (
            .O(N__28107),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    InMux I__3842 (
            .O(N__28104),
            .I(N__28098));
    InMux I__3841 (
            .O(N__28103),
            .I(N__28098));
    LocalMux I__3840 (
            .O(N__28098),
            .I(N__28095));
    Odrv4 I__3839 (
            .O(N__28095),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    InMux I__3838 (
            .O(N__28092),
            .I(N__28089));
    LocalMux I__3837 (
            .O(N__28089),
            .I(N__28086));
    Odrv4 I__3836 (
            .O(N__28086),
            .I(\pid_alt.m21_e_9 ));
    InMux I__3835 (
            .O(N__28083),
            .I(N__28080));
    LocalMux I__3834 (
            .O(N__28080),
            .I(\pid_alt.m21_e_10 ));
    InMux I__3833 (
            .O(N__28077),
            .I(N__28073));
    InMux I__3832 (
            .O(N__28076),
            .I(N__28070));
    LocalMux I__3831 (
            .O(N__28073),
            .I(\pid_alt.N_9_0 ));
    LocalMux I__3830 (
            .O(N__28070),
            .I(\pid_alt.N_9_0 ));
    CascadeMux I__3829 (
            .O(N__28065),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNIO7B05Z0Z_21_cascade_ ));
    CascadeMux I__3828 (
            .O(N__28062),
            .I(\pid_alt.un1_reset_1_0_i_cascade_ ));
    CascadeMux I__3827 (
            .O(N__28059),
            .I(N__28055));
    CascadeMux I__3826 (
            .O(N__28058),
            .I(N__28051));
    InMux I__3825 (
            .O(N__28055),
            .I(N__28048));
    InMux I__3824 (
            .O(N__28054),
            .I(N__28043));
    InMux I__3823 (
            .O(N__28051),
            .I(N__28043));
    LocalMux I__3822 (
            .O(N__28048),
            .I(N__28040));
    LocalMux I__3821 (
            .O(N__28043),
            .I(N__28034));
    Span4Mux_h I__3820 (
            .O(N__28040),
            .I(N__28034));
    InMux I__3819 (
            .O(N__28039),
            .I(N__28031));
    Span4Mux_v I__3818 (
            .O(N__28034),
            .I(N__28028));
    LocalMux I__3817 (
            .O(N__28031),
            .I(N__28025));
    Span4Mux_v I__3816 (
            .O(N__28028),
            .I(N__28022));
    Span12Mux_v I__3815 (
            .O(N__28025),
            .I(N__28019));
    Odrv4 I__3814 (
            .O(N__28022),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    Odrv12 I__3813 (
            .O(N__28019),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    InMux I__3812 (
            .O(N__28014),
            .I(N__28010));
    InMux I__3811 (
            .O(N__28013),
            .I(N__28007));
    LocalMux I__3810 (
            .O(N__28010),
            .I(N__28001));
    LocalMux I__3809 (
            .O(N__28007),
            .I(N__28001));
    InMux I__3808 (
            .O(N__28006),
            .I(N__27998));
    Span4Mux_v I__3807 (
            .O(N__28001),
            .I(N__27995));
    LocalMux I__3806 (
            .O(N__27998),
            .I(N__27992));
    Odrv4 I__3805 (
            .O(N__27995),
            .I(\pid_alt.error_i_acumm7lto13 ));
    Odrv4 I__3804 (
            .O(N__27992),
            .I(\pid_alt.error_i_acumm7lto13 ));
    InMux I__3803 (
            .O(N__27987),
            .I(N__27984));
    LocalMux I__3802 (
            .O(N__27984),
            .I(N__27980));
    InMux I__3801 (
            .O(N__27983),
            .I(N__27976));
    Span4Mux_v I__3800 (
            .O(N__27980),
            .I(N__27973));
    InMux I__3799 (
            .O(N__27979),
            .I(N__27970));
    LocalMux I__3798 (
            .O(N__27976),
            .I(N__27967));
    Odrv4 I__3797 (
            .O(N__27973),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14 ));
    LocalMux I__3796 (
            .O(N__27970),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14 ));
    Odrv4 I__3795 (
            .O(N__27967),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14 ));
    InMux I__3794 (
            .O(N__27960),
            .I(N__27957));
    LocalMux I__3793 (
            .O(N__27957),
            .I(N__27954));
    Odrv4 I__3792 (
            .O(N__27954),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    CEMux I__3791 (
            .O(N__27951),
            .I(N__27947));
    CEMux I__3790 (
            .O(N__27950),
            .I(N__27944));
    LocalMux I__3789 (
            .O(N__27947),
            .I(\pid_alt.N_72_i_0 ));
    LocalMux I__3788 (
            .O(N__27944),
            .I(\pid_alt.N_72_i_0 ));
    CascadeMux I__3787 (
            .O(N__27939),
            .I(\pid_alt.un1_reset_1_cascade_ ));
    CascadeMux I__3786 (
            .O(N__27936),
            .I(\pid_alt.source_pid_9_0_tz_6_cascade_ ));
    InMux I__3785 (
            .O(N__27933),
            .I(N__27929));
    InMux I__3784 (
            .O(N__27932),
            .I(N__27926));
    LocalMux I__3783 (
            .O(N__27929),
            .I(N__27922));
    LocalMux I__3782 (
            .O(N__27926),
            .I(N__27919));
    InMux I__3781 (
            .O(N__27925),
            .I(N__27916));
    Odrv4 I__3780 (
            .O(N__27922),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    Odrv4 I__3779 (
            .O(N__27919),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__3778 (
            .O(N__27916),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    CascadeMux I__3777 (
            .O(N__27909),
            .I(\pid_alt.m21_e_0_cascade_ ));
    CascadeMux I__3776 (
            .O(N__27906),
            .I(N__27901));
    CascadeMux I__3775 (
            .O(N__27905),
            .I(N__27897));
    InMux I__3774 (
            .O(N__27904),
            .I(N__27888));
    InMux I__3773 (
            .O(N__27901),
            .I(N__27888));
    InMux I__3772 (
            .O(N__27900),
            .I(N__27888));
    InMux I__3771 (
            .O(N__27897),
            .I(N__27883));
    InMux I__3770 (
            .O(N__27896),
            .I(N__27883));
    InMux I__3769 (
            .O(N__27895),
            .I(N__27880));
    LocalMux I__3768 (
            .O(N__27888),
            .I(\pid_alt.error_i_acumm7lto4 ));
    LocalMux I__3767 (
            .O(N__27883),
            .I(\pid_alt.error_i_acumm7lto4 ));
    LocalMux I__3766 (
            .O(N__27880),
            .I(\pid_alt.error_i_acumm7lto4 ));
    InMux I__3765 (
            .O(N__27873),
            .I(N__27870));
    LocalMux I__3764 (
            .O(N__27870),
            .I(\pid_alt.m35_e_3 ));
    InMux I__3763 (
            .O(N__27867),
            .I(N__27862));
    InMux I__3762 (
            .O(N__27866),
            .I(N__27857));
    InMux I__3761 (
            .O(N__27865),
            .I(N__27857));
    LocalMux I__3760 (
            .O(N__27862),
            .I(N__27854));
    LocalMux I__3759 (
            .O(N__27857),
            .I(N__27851));
    Span4Mux_v I__3758 (
            .O(N__27854),
            .I(N__27848));
    Span4Mux_v I__3757 (
            .O(N__27851),
            .I(N__27845));
    Odrv4 I__3756 (
            .O(N__27848),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    Odrv4 I__3755 (
            .O(N__27845),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    InMux I__3754 (
            .O(N__27840),
            .I(N__27837));
    LocalMux I__3753 (
            .O(N__27837),
            .I(N__27832));
    InMux I__3752 (
            .O(N__27836),
            .I(N__27827));
    InMux I__3751 (
            .O(N__27835),
            .I(N__27827));
    Odrv4 I__3750 (
            .O(N__27832),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    LocalMux I__3749 (
            .O(N__27827),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    InMux I__3748 (
            .O(N__27822),
            .I(N__27819));
    LocalMux I__3747 (
            .O(N__27819),
            .I(N__27816));
    Span4Mux_v I__3746 (
            .O(N__27816),
            .I(N__27811));
    InMux I__3745 (
            .O(N__27815),
            .I(N__27806));
    InMux I__3744 (
            .O(N__27814),
            .I(N__27806));
    Odrv4 I__3743 (
            .O(N__27811),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ));
    LocalMux I__3742 (
            .O(N__27806),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ));
    CascadeMux I__3741 (
            .O(N__27801),
            .I(N__27798));
    InMux I__3740 (
            .O(N__27798),
            .I(N__27793));
    InMux I__3739 (
            .O(N__27797),
            .I(N__27788));
    InMux I__3738 (
            .O(N__27796),
            .I(N__27788));
    LocalMux I__3737 (
            .O(N__27793),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__3736 (
            .O(N__27788),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    InMux I__3735 (
            .O(N__27783),
            .I(N__27778));
    InMux I__3734 (
            .O(N__27782),
            .I(N__27773));
    InMux I__3733 (
            .O(N__27781),
            .I(N__27773));
    LocalMux I__3732 (
            .O(N__27778),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__3731 (
            .O(N__27773),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    CascadeMux I__3730 (
            .O(N__27768),
            .I(N__27763));
    CascadeMux I__3729 (
            .O(N__27767),
            .I(N__27760));
    InMux I__3728 (
            .O(N__27766),
            .I(N__27757));
    InMux I__3727 (
            .O(N__27763),
            .I(N__27752));
    InMux I__3726 (
            .O(N__27760),
            .I(N__27752));
    LocalMux I__3725 (
            .O(N__27757),
            .I(N__27749));
    LocalMux I__3724 (
            .O(N__27752),
            .I(N__27746));
    Span4Mux_h I__3723 (
            .O(N__27749),
            .I(N__27743));
    Span4Mux_h I__3722 (
            .O(N__27746),
            .I(N__27740));
    Odrv4 I__3721 (
            .O(N__27743),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    Odrv4 I__3720 (
            .O(N__27740),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    InMux I__3719 (
            .O(N__27735),
            .I(N__27728));
    InMux I__3718 (
            .O(N__27734),
            .I(N__27728));
    InMux I__3717 (
            .O(N__27733),
            .I(N__27725));
    LocalMux I__3716 (
            .O(N__27728),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__3715 (
            .O(N__27725),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    InMux I__3714 (
            .O(N__27720),
            .I(N__27716));
    InMux I__3713 (
            .O(N__27719),
            .I(N__27713));
    LocalMux I__3712 (
            .O(N__27716),
            .I(N__27708));
    LocalMux I__3711 (
            .O(N__27713),
            .I(N__27708));
    Span4Mux_h I__3710 (
            .O(N__27708),
            .I(N__27705));
    Odrv4 I__3709 (
            .O(N__27705),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    InMux I__3708 (
            .O(N__27702),
            .I(N__27698));
    InMux I__3707 (
            .O(N__27701),
            .I(N__27695));
    LocalMux I__3706 (
            .O(N__27698),
            .I(N__27692));
    LocalMux I__3705 (
            .O(N__27695),
            .I(N__27689));
    Odrv12 I__3704 (
            .O(N__27692),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    Odrv4 I__3703 (
            .O(N__27689),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    CascadeMux I__3702 (
            .O(N__27684),
            .I(\pid_alt.m21_e_8_cascade_ ));
    InMux I__3701 (
            .O(N__27681),
            .I(N__27678));
    LocalMux I__3700 (
            .O(N__27678),
            .I(N__27673));
    InMux I__3699 (
            .O(N__27677),
            .I(N__27670));
    InMux I__3698 (
            .O(N__27676),
            .I(N__27667));
    Odrv4 I__3697 (
            .O(N__27673),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__3696 (
            .O(N__27670),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__3695 (
            .O(N__27667),
            .I(\pid_alt.error_i_acumm7lto12 ));
    InMux I__3694 (
            .O(N__27660),
            .I(N__27657));
    LocalMux I__3693 (
            .O(N__27657),
            .I(\pid_alt.m21_e_2 ));
    InMux I__3692 (
            .O(N__27654),
            .I(N__27651));
    LocalMux I__3691 (
            .O(N__27651),
            .I(N__27648));
    Span4Mux_h I__3690 (
            .O(N__27648),
            .I(N__27643));
    InMux I__3689 (
            .O(N__27647),
            .I(N__27640));
    InMux I__3688 (
            .O(N__27646),
            .I(N__27637));
    Odrv4 I__3687 (
            .O(N__27643),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    LocalMux I__3686 (
            .O(N__27640),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    LocalMux I__3685 (
            .O(N__27637),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    InMux I__3684 (
            .O(N__27630),
            .I(N__27625));
    InMux I__3683 (
            .O(N__27629),
            .I(N__27620));
    InMux I__3682 (
            .O(N__27628),
            .I(N__27620));
    LocalMux I__3681 (
            .O(N__27625),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__3680 (
            .O(N__27620),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    CEMux I__3679 (
            .O(N__27615),
            .I(N__27546));
    CEMux I__3678 (
            .O(N__27614),
            .I(N__27546));
    CEMux I__3677 (
            .O(N__27613),
            .I(N__27546));
    CEMux I__3676 (
            .O(N__27612),
            .I(N__27546));
    CEMux I__3675 (
            .O(N__27611),
            .I(N__27546));
    CEMux I__3674 (
            .O(N__27610),
            .I(N__27546));
    CEMux I__3673 (
            .O(N__27609),
            .I(N__27546));
    CEMux I__3672 (
            .O(N__27608),
            .I(N__27546));
    CEMux I__3671 (
            .O(N__27607),
            .I(N__27546));
    CEMux I__3670 (
            .O(N__27606),
            .I(N__27546));
    CEMux I__3669 (
            .O(N__27605),
            .I(N__27546));
    CEMux I__3668 (
            .O(N__27604),
            .I(N__27546));
    CEMux I__3667 (
            .O(N__27603),
            .I(N__27546));
    CEMux I__3666 (
            .O(N__27602),
            .I(N__27546));
    CEMux I__3665 (
            .O(N__27601),
            .I(N__27546));
    CEMux I__3664 (
            .O(N__27600),
            .I(N__27546));
    CEMux I__3663 (
            .O(N__27599),
            .I(N__27546));
    CEMux I__3662 (
            .O(N__27598),
            .I(N__27546));
    CEMux I__3661 (
            .O(N__27597),
            .I(N__27546));
    CEMux I__3660 (
            .O(N__27596),
            .I(N__27546));
    CEMux I__3659 (
            .O(N__27595),
            .I(N__27546));
    CEMux I__3658 (
            .O(N__27594),
            .I(N__27546));
    CEMux I__3657 (
            .O(N__27593),
            .I(N__27546));
    GlobalMux I__3656 (
            .O(N__27546),
            .I(N__27543));
    gio2CtrlBuf I__3655 (
            .O(N__27543),
            .I(\pid_alt.state_0_g_0 ));
    InMux I__3654 (
            .O(N__27540),
            .I(N__27536));
    InMux I__3653 (
            .O(N__27539),
            .I(N__27533));
    LocalMux I__3652 (
            .O(N__27536),
            .I(\Commands_frame_decoder.N_416 ));
    LocalMux I__3651 (
            .O(N__27533),
            .I(\Commands_frame_decoder.N_416 ));
    CascadeMux I__3650 (
            .O(N__27528),
            .I(\Commands_frame_decoder.N_379_cascade_ ));
    InMux I__3649 (
            .O(N__27525),
            .I(N__27517));
    InMux I__3648 (
            .O(N__27524),
            .I(N__27517));
    InMux I__3647 (
            .O(N__27523),
            .I(N__27512));
    InMux I__3646 (
            .O(N__27522),
            .I(N__27512));
    LocalMux I__3645 (
            .O(N__27517),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__3644 (
            .O(N__27512),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    InMux I__3643 (
            .O(N__27507),
            .I(N__27504));
    LocalMux I__3642 (
            .O(N__27504),
            .I(\Commands_frame_decoder.N_412 ));
    CascadeMux I__3641 (
            .O(N__27501),
            .I(N__27498));
    InMux I__3640 (
            .O(N__27498),
            .I(N__27492));
    InMux I__3639 (
            .O(N__27497),
            .I(N__27492));
    LocalMux I__3638 (
            .O(N__27492),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    CEMux I__3637 (
            .O(N__27489),
            .I(N__27485));
    CEMux I__3636 (
            .O(N__27488),
            .I(N__27480));
    LocalMux I__3635 (
            .O(N__27485),
            .I(N__27477));
    CEMux I__3634 (
            .O(N__27484),
            .I(N__27474));
    CEMux I__3633 (
            .O(N__27483),
            .I(N__27471));
    LocalMux I__3632 (
            .O(N__27480),
            .I(N__27468));
    Span4Mux_v I__3631 (
            .O(N__27477),
            .I(N__27463));
    LocalMux I__3630 (
            .O(N__27474),
            .I(N__27463));
    LocalMux I__3629 (
            .O(N__27471),
            .I(N__27460));
    Span4Mux_v I__3628 (
            .O(N__27468),
            .I(N__27457));
    Span4Mux_v I__3627 (
            .O(N__27463),
            .I(N__27454));
    Span4Mux_h I__3626 (
            .O(N__27460),
            .I(N__27451));
    Span4Mux_v I__3625 (
            .O(N__27457),
            .I(N__27448));
    Span4Mux_v I__3624 (
            .O(N__27454),
            .I(N__27445));
    Span4Mux_v I__3623 (
            .O(N__27451),
            .I(N__27442));
    Span4Mux_v I__3622 (
            .O(N__27448),
            .I(N__27439));
    Span4Mux_h I__3621 (
            .O(N__27445),
            .I(N__27436));
    Span4Mux_v I__3620 (
            .O(N__27442),
            .I(N__27433));
    Odrv4 I__3619 (
            .O(N__27439),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    Odrv4 I__3618 (
            .O(N__27436),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    Odrv4 I__3617 (
            .O(N__27433),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    InMux I__3616 (
            .O(N__27426),
            .I(N__27422));
    InMux I__3615 (
            .O(N__27425),
            .I(N__27419));
    LocalMux I__3614 (
            .O(N__27422),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    LocalMux I__3613 (
            .O(N__27419),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    InMux I__3612 (
            .O(N__27414),
            .I(N__27396));
    InMux I__3611 (
            .O(N__27413),
            .I(N__27396));
    InMux I__3610 (
            .O(N__27412),
            .I(N__27396));
    InMux I__3609 (
            .O(N__27411),
            .I(N__27396));
    InMux I__3608 (
            .O(N__27410),
            .I(N__27396));
    InMux I__3607 (
            .O(N__27409),
            .I(N__27396));
    LocalMux I__3606 (
            .O(N__27396),
            .I(N__27390));
    InMux I__3605 (
            .O(N__27395),
            .I(N__27383));
    InMux I__3604 (
            .O(N__27394),
            .I(N__27383));
    InMux I__3603 (
            .O(N__27393),
            .I(N__27383));
    Odrv4 I__3602 (
            .O(N__27390),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12 ));
    LocalMux I__3601 (
            .O(N__27383),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12 ));
    InMux I__3600 (
            .O(N__27378),
            .I(N__27374));
    InMux I__3599 (
            .O(N__27377),
            .I(N__27371));
    LocalMux I__3598 (
            .O(N__27374),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    LocalMux I__3597 (
            .O(N__27371),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    InMux I__3596 (
            .O(N__27366),
            .I(N__27363));
    LocalMux I__3595 (
            .O(N__27363),
            .I(N__27359));
    InMux I__3594 (
            .O(N__27362),
            .I(N__27356));
    Odrv4 I__3593 (
            .O(N__27359),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__3592 (
            .O(N__27356),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    CascadeMux I__3591 (
            .O(N__27351),
            .I(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ));
    CascadeMux I__3590 (
            .O(N__27348),
            .I(\Commands_frame_decoder.N_416_cascade_ ));
    InMux I__3589 (
            .O(N__27345),
            .I(N__27342));
    LocalMux I__3588 (
            .O(N__27342),
            .I(\Commands_frame_decoder.N_382 ));
    InMux I__3587 (
            .O(N__27339),
            .I(N__27336));
    LocalMux I__3586 (
            .O(N__27336),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_2_2 ));
    InMux I__3585 (
            .O(N__27333),
            .I(N__27329));
    InMux I__3584 (
            .O(N__27332),
            .I(N__27326));
    LocalMux I__3583 (
            .O(N__27329),
            .I(\Commands_frame_decoder.N_376_2 ));
    LocalMux I__3582 (
            .O(N__27326),
            .I(\Commands_frame_decoder.N_376_2 ));
    InMux I__3581 (
            .O(N__27321),
            .I(N__27318));
    LocalMux I__3580 (
            .O(N__27318),
            .I(\Commands_frame_decoder.N_377 ));
    CascadeMux I__3579 (
            .O(N__27315),
            .I(\Commands_frame_decoder.N_376_cascade_ ));
    InMux I__3578 (
            .O(N__27312),
            .I(N__27309));
    LocalMux I__3577 (
            .O(N__27309),
            .I(\Commands_frame_decoder.N_379 ));
    InMux I__3576 (
            .O(N__27306),
            .I(N__27302));
    InMux I__3575 (
            .O(N__27305),
            .I(N__27299));
    LocalMux I__3574 (
            .O(N__27302),
            .I(N__27296));
    LocalMux I__3573 (
            .O(N__27299),
            .I(N__27293));
    Span4Mux_v I__3572 (
            .O(N__27296),
            .I(N__27290));
    Span4Mux_v I__3571 (
            .O(N__27293),
            .I(N__27287));
    Odrv4 I__3570 (
            .O(N__27290),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    Odrv4 I__3569 (
            .O(N__27287),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    InMux I__3568 (
            .O(N__27282),
            .I(N__27279));
    LocalMux I__3567 (
            .O(N__27279),
            .I(N__27276));
    Span4Mux_h I__3566 (
            .O(N__27276),
            .I(N__27272));
    InMux I__3565 (
            .O(N__27275),
            .I(N__27269));
    Sp12to4 I__3564 (
            .O(N__27272),
            .I(N__27266));
    LocalMux I__3563 (
            .O(N__27269),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    Odrv12 I__3562 (
            .O(N__27266),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    InMux I__3561 (
            .O(N__27261),
            .I(N__27255));
    InMux I__3560 (
            .O(N__27260),
            .I(N__27255));
    LocalMux I__3559 (
            .O(N__27255),
            .I(N__27252));
    Span4Mux_v I__3558 (
            .O(N__27252),
            .I(N__27248));
    InMux I__3557 (
            .O(N__27251),
            .I(N__27245));
    Sp12to4 I__3556 (
            .O(N__27248),
            .I(N__27240));
    LocalMux I__3555 (
            .O(N__27245),
            .I(N__27240));
    Span12Mux_s7_h I__3554 (
            .O(N__27240),
            .I(N__27237));
    Span12Mux_v I__3553 (
            .O(N__27237),
            .I(N__27234));
    Odrv12 I__3552 (
            .O(N__27234),
            .I(\pid_alt.error_d_regZ0Z_19 ));
    InMux I__3551 (
            .O(N__27231),
            .I(N__27228));
    LocalMux I__3550 (
            .O(N__27228),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ));
    InMux I__3549 (
            .O(N__27225),
            .I(N__27222));
    LocalMux I__3548 (
            .O(N__27222),
            .I(N__27218));
    CascadeMux I__3547 (
            .O(N__27221),
            .I(N__27215));
    Span12Mux_h I__3546 (
            .O(N__27218),
            .I(N__27212));
    InMux I__3545 (
            .O(N__27215),
            .I(N__27209));
    Odrv12 I__3544 (
            .O(N__27212),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    LocalMux I__3543 (
            .O(N__27209),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    CascadeMux I__3542 (
            .O(N__27204),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ));
    InMux I__3541 (
            .O(N__27201),
            .I(N__27194));
    InMux I__3540 (
            .O(N__27200),
            .I(N__27194));
    InMux I__3539 (
            .O(N__27199),
            .I(N__27191));
    LocalMux I__3538 (
            .O(N__27194),
            .I(N__27188));
    LocalMux I__3537 (
            .O(N__27191),
            .I(N__27185));
    Span4Mux_v I__3536 (
            .O(N__27188),
            .I(N__27182));
    Odrv12 I__3535 (
            .O(N__27185),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    Odrv4 I__3534 (
            .O(N__27182),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    InMux I__3533 (
            .O(N__27177),
            .I(N__27174));
    LocalMux I__3532 (
            .O(N__27174),
            .I(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ));
    InMux I__3531 (
            .O(N__27171),
            .I(N__27165));
    InMux I__3530 (
            .O(N__27170),
            .I(N__27165));
    LocalMux I__3529 (
            .O(N__27165),
            .I(N__27162));
    Span4Mux_h I__3528 (
            .O(N__27162),
            .I(N__27159));
    Odrv4 I__3527 (
            .O(N__27159),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    InMux I__3526 (
            .O(N__27156),
            .I(N__27150));
    InMux I__3525 (
            .O(N__27155),
            .I(N__27150));
    LocalMux I__3524 (
            .O(N__27150),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    InMux I__3523 (
            .O(N__27147),
            .I(N__27138));
    InMux I__3522 (
            .O(N__27146),
            .I(N__27138));
    InMux I__3521 (
            .O(N__27145),
            .I(N__27138));
    LocalMux I__3520 (
            .O(N__27138),
            .I(N__27135));
    Span4Mux_h I__3519 (
            .O(N__27135),
            .I(N__27132));
    Sp12to4 I__3518 (
            .O(N__27132),
            .I(N__27129));
    Span12Mux_v I__3517 (
            .O(N__27129),
            .I(N__27126));
    Odrv12 I__3516 (
            .O(N__27126),
            .I(\pid_alt.error_d_regZ0Z_20 ));
    CascadeMux I__3515 (
            .O(N__27123),
            .I(N__27120));
    InMux I__3514 (
            .O(N__27120),
            .I(N__27114));
    InMux I__3513 (
            .O(N__27119),
            .I(N__27107));
    InMux I__3512 (
            .O(N__27118),
            .I(N__27107));
    InMux I__3511 (
            .O(N__27117),
            .I(N__27107));
    LocalMux I__3510 (
            .O(N__27114),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ));
    LocalMux I__3509 (
            .O(N__27107),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ));
    CascadeMux I__3508 (
            .O(N__27102),
            .I(N__27098));
    InMux I__3507 (
            .O(N__27101),
            .I(N__27095));
    InMux I__3506 (
            .O(N__27098),
            .I(N__27092));
    LocalMux I__3505 (
            .O(N__27095),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ));
    LocalMux I__3504 (
            .O(N__27092),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ));
    CascadeMux I__3503 (
            .O(N__27087),
            .I(N__27083));
    InMux I__3502 (
            .O(N__27086),
            .I(N__27076));
    InMux I__3501 (
            .O(N__27083),
            .I(N__27069));
    InMux I__3500 (
            .O(N__27082),
            .I(N__27069));
    InMux I__3499 (
            .O(N__27081),
            .I(N__27069));
    InMux I__3498 (
            .O(N__27080),
            .I(N__27064));
    InMux I__3497 (
            .O(N__27079),
            .I(N__27064));
    LocalMux I__3496 (
            .O(N__27076),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    LocalMux I__3495 (
            .O(N__27069),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    LocalMux I__3494 (
            .O(N__27064),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    CascadeMux I__3493 (
            .O(N__27057),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20_cascade_ ));
    InMux I__3492 (
            .O(N__27054),
            .I(N__27046));
    InMux I__3491 (
            .O(N__27053),
            .I(N__27043));
    InMux I__3490 (
            .O(N__27052),
            .I(N__27034));
    InMux I__3489 (
            .O(N__27051),
            .I(N__27034));
    InMux I__3488 (
            .O(N__27050),
            .I(N__27034));
    InMux I__3487 (
            .O(N__27049),
            .I(N__27034));
    LocalMux I__3486 (
            .O(N__27046),
            .I(N__27031));
    LocalMux I__3485 (
            .O(N__27043),
            .I(N__27026));
    LocalMux I__3484 (
            .O(N__27034),
            .I(N__27026));
    Span4Mux_v I__3483 (
            .O(N__27031),
            .I(N__27023));
    Odrv12 I__3482 (
            .O(N__27026),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    Odrv4 I__3481 (
            .O(N__27023),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    InMux I__3480 (
            .O(N__27018),
            .I(N__27015));
    LocalMux I__3479 (
            .O(N__27015),
            .I(\pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20 ));
    CascadeMux I__3478 (
            .O(N__27012),
            .I(N__27008));
    InMux I__3477 (
            .O(N__27011),
            .I(N__27005));
    InMux I__3476 (
            .O(N__27008),
            .I(N__27001));
    LocalMux I__3475 (
            .O(N__27005),
            .I(N__26998));
    InMux I__3474 (
            .O(N__27004),
            .I(N__26995));
    LocalMux I__3473 (
            .O(N__27001),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    Odrv4 I__3472 (
            .O(N__26998),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    LocalMux I__3471 (
            .O(N__26995),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    CascadeMux I__3470 (
            .O(N__26988),
            .I(N__26984));
    InMux I__3469 (
            .O(N__26987),
            .I(N__26979));
    InMux I__3468 (
            .O(N__26984),
            .I(N__26979));
    LocalMux I__3467 (
            .O(N__26979),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    InMux I__3466 (
            .O(N__26976),
            .I(N__26970));
    InMux I__3465 (
            .O(N__26975),
            .I(N__26970));
    LocalMux I__3464 (
            .O(N__26970),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ));
    CascadeMux I__3463 (
            .O(N__26967),
            .I(N__26964));
    InMux I__3462 (
            .O(N__26964),
            .I(N__26960));
    InMux I__3461 (
            .O(N__26963),
            .I(N__26957));
    LocalMux I__3460 (
            .O(N__26960),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    LocalMux I__3459 (
            .O(N__26957),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    InMux I__3458 (
            .O(N__26952),
            .I(N__26943));
    InMux I__3457 (
            .O(N__26951),
            .I(N__26943));
    InMux I__3456 (
            .O(N__26950),
            .I(N__26943));
    LocalMux I__3455 (
            .O(N__26943),
            .I(N__26940));
    Span4Mux_v I__3454 (
            .O(N__26940),
            .I(N__26937));
    Span4Mux_v I__3453 (
            .O(N__26937),
            .I(N__26934));
    Span4Mux_h I__3452 (
            .O(N__26934),
            .I(N__26931));
    Span4Mux_v I__3451 (
            .O(N__26931),
            .I(N__26928));
    Odrv4 I__3450 (
            .O(N__26928),
            .I(\pid_alt.error_d_regZ0Z_16 ));
    CascadeMux I__3449 (
            .O(N__26925),
            .I(N__26922));
    InMux I__3448 (
            .O(N__26922),
            .I(N__26916));
    InMux I__3447 (
            .O(N__26921),
            .I(N__26916));
    LocalMux I__3446 (
            .O(N__26916),
            .I(\pid_alt.error_d_reg_prevZ0Z_16 ));
    InMux I__3445 (
            .O(N__26913),
            .I(N__26907));
    InMux I__3444 (
            .O(N__26912),
            .I(N__26907));
    LocalMux I__3443 (
            .O(N__26907),
            .I(N__26904));
    Span4Mux_h I__3442 (
            .O(N__26904),
            .I(N__26901));
    Span4Mux_s1_h I__3441 (
            .O(N__26901),
            .I(N__26898));
    Odrv4 I__3440 (
            .O(N__26898),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    InMux I__3439 (
            .O(N__26895),
            .I(N__26892));
    LocalMux I__3438 (
            .O(N__26892),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ));
    CascadeMux I__3437 (
            .O(N__26889),
            .I(N__26885));
    InMux I__3436 (
            .O(N__26888),
            .I(N__26882));
    InMux I__3435 (
            .O(N__26885),
            .I(N__26879));
    LocalMux I__3434 (
            .O(N__26882),
            .I(N__26874));
    LocalMux I__3433 (
            .O(N__26879),
            .I(N__26874));
    Span4Mux_v I__3432 (
            .O(N__26874),
            .I(N__26871));
    Odrv4 I__3431 (
            .O(N__26871),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    CascadeMux I__3430 (
            .O(N__26868),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ));
    InMux I__3429 (
            .O(N__26865),
            .I(N__26860));
    InMux I__3428 (
            .O(N__26864),
            .I(N__26855));
    InMux I__3427 (
            .O(N__26863),
            .I(N__26855));
    LocalMux I__3426 (
            .O(N__26860),
            .I(N__26852));
    LocalMux I__3425 (
            .O(N__26855),
            .I(N__26849));
    Span4Mux_h I__3424 (
            .O(N__26852),
            .I(N__26846));
    Span4Mux_v I__3423 (
            .O(N__26849),
            .I(N__26843));
    Odrv4 I__3422 (
            .O(N__26846),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    Odrv4 I__3421 (
            .O(N__26843),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    InMux I__3420 (
            .O(N__26838),
            .I(N__26835));
    LocalMux I__3419 (
            .O(N__26835),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ));
    CascadeMux I__3418 (
            .O(N__26832),
            .I(\pid_alt.un1_pid_prereg_236_1_cascade_ ));
    InMux I__3417 (
            .O(N__26829),
            .I(N__26825));
    InMux I__3416 (
            .O(N__26828),
            .I(N__26822));
    LocalMux I__3415 (
            .O(N__26825),
            .I(N__26819));
    LocalMux I__3414 (
            .O(N__26822),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    Odrv4 I__3413 (
            .O(N__26819),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    InMux I__3412 (
            .O(N__26814),
            .I(N__26810));
    InMux I__3411 (
            .O(N__26813),
            .I(N__26807));
    LocalMux I__3410 (
            .O(N__26810),
            .I(N__26804));
    LocalMux I__3409 (
            .O(N__26807),
            .I(N__26801));
    Span4Mux_h I__3408 (
            .O(N__26804),
            .I(N__26798));
    Span4Mux_h I__3407 (
            .O(N__26801),
            .I(N__26795));
    Span4Mux_v I__3406 (
            .O(N__26798),
            .I(N__26792));
    Odrv4 I__3405 (
            .O(N__26795),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    Odrv4 I__3404 (
            .O(N__26792),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    InMux I__3403 (
            .O(N__26787),
            .I(N__26781));
    InMux I__3402 (
            .O(N__26786),
            .I(N__26781));
    LocalMux I__3401 (
            .O(N__26781),
            .I(N__26777));
    InMux I__3400 (
            .O(N__26780),
            .I(N__26774));
    Span4Mux_v I__3399 (
            .O(N__26777),
            .I(N__26769));
    LocalMux I__3398 (
            .O(N__26774),
            .I(N__26769));
    Span4Mux_v I__3397 (
            .O(N__26769),
            .I(N__26766));
    Span4Mux_v I__3396 (
            .O(N__26766),
            .I(N__26763));
    Odrv4 I__3395 (
            .O(N__26763),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    InMux I__3394 (
            .O(N__26760),
            .I(N__26754));
    InMux I__3393 (
            .O(N__26759),
            .I(N__26754));
    LocalMux I__3392 (
            .O(N__26754),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ));
    CascadeMux I__3391 (
            .O(N__26751),
            .I(N__26747));
    CascadeMux I__3390 (
            .O(N__26750),
            .I(N__26744));
    InMux I__3389 (
            .O(N__26747),
            .I(N__26741));
    InMux I__3388 (
            .O(N__26744),
            .I(N__26738));
    LocalMux I__3387 (
            .O(N__26741),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    LocalMux I__3386 (
            .O(N__26738),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    InMux I__3385 (
            .O(N__26733),
            .I(N__26724));
    InMux I__3384 (
            .O(N__26732),
            .I(N__26724));
    InMux I__3383 (
            .O(N__26731),
            .I(N__26724));
    LocalMux I__3382 (
            .O(N__26724),
            .I(N__26721));
    Span4Mux_v I__3381 (
            .O(N__26721),
            .I(N__26718));
    Span4Mux_v I__3380 (
            .O(N__26718),
            .I(N__26715));
    Odrv4 I__3379 (
            .O(N__26715),
            .I(\pid_alt.error_d_regZ0Z_7 ));
    CascadeMux I__3378 (
            .O(N__26712),
            .I(N__26709));
    InMux I__3377 (
            .O(N__26709),
            .I(N__26703));
    InMux I__3376 (
            .O(N__26708),
            .I(N__26703));
    LocalMux I__3375 (
            .O(N__26703),
            .I(\pid_alt.error_d_reg_prevZ0Z_7 ));
    InMux I__3374 (
            .O(N__26700),
            .I(N__26694));
    InMux I__3373 (
            .O(N__26699),
            .I(N__26694));
    LocalMux I__3372 (
            .O(N__26694),
            .I(N__26691));
    Span4Mux_h I__3371 (
            .O(N__26691),
            .I(N__26688));
    Odrv4 I__3370 (
            .O(N__26688),
            .I(\pid_alt.error_p_regZ0Z_7 ));
    InMux I__3369 (
            .O(N__26685),
            .I(N__26682));
    LocalMux I__3368 (
            .O(N__26682),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    InMux I__3367 (
            .O(N__26679),
            .I(N__26673));
    InMux I__3366 (
            .O(N__26678),
            .I(N__26673));
    LocalMux I__3365 (
            .O(N__26673),
            .I(N__26670));
    Span4Mux_v I__3364 (
            .O(N__26670),
            .I(N__26667));
    Odrv4 I__3363 (
            .O(N__26667),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ));
    InMux I__3362 (
            .O(N__26664),
            .I(N__26660));
    CascadeMux I__3361 (
            .O(N__26663),
            .I(N__26657));
    LocalMux I__3360 (
            .O(N__26660),
            .I(N__26654));
    InMux I__3359 (
            .O(N__26657),
            .I(N__26651));
    Span4Mux_h I__3358 (
            .O(N__26654),
            .I(N__26648));
    LocalMux I__3357 (
            .O(N__26651),
            .I(N__26645));
    Span4Mux_v I__3356 (
            .O(N__26648),
            .I(N__26642));
    Span4Mux_v I__3355 (
            .O(N__26645),
            .I(N__26639));
    Odrv4 I__3354 (
            .O(N__26642),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    Odrv4 I__3353 (
            .O(N__26639),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    CascadeMux I__3352 (
            .O(N__26634),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ));
    InMux I__3351 (
            .O(N__26631),
            .I(N__26625));
    InMux I__3350 (
            .O(N__26630),
            .I(N__26625));
    LocalMux I__3349 (
            .O(N__26625),
            .I(N__26621));
    InMux I__3348 (
            .O(N__26624),
            .I(N__26618));
    Span4Mux_v I__3347 (
            .O(N__26621),
            .I(N__26615));
    LocalMux I__3346 (
            .O(N__26618),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    Odrv4 I__3345 (
            .O(N__26615),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    InMux I__3344 (
            .O(N__26610),
            .I(N__26607));
    LocalMux I__3343 (
            .O(N__26607),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ));
    CascadeMux I__3342 (
            .O(N__26604),
            .I(N__26601));
    InMux I__3341 (
            .O(N__26601),
            .I(N__26598));
    LocalMux I__3340 (
            .O(N__26598),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ));
    InMux I__3339 (
            .O(N__26595),
            .I(N__26592));
    LocalMux I__3338 (
            .O(N__26592),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ));
    CascadeMux I__3337 (
            .O(N__26589),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ));
    InMux I__3336 (
            .O(N__26586),
            .I(N__26581));
    InMux I__3335 (
            .O(N__26585),
            .I(N__26576));
    InMux I__3334 (
            .O(N__26584),
            .I(N__26576));
    LocalMux I__3333 (
            .O(N__26581),
            .I(N__26573));
    LocalMux I__3332 (
            .O(N__26576),
            .I(N__26570));
    Span4Mux_v I__3331 (
            .O(N__26573),
            .I(N__26565));
    Span4Mux_v I__3330 (
            .O(N__26570),
            .I(N__26565));
    Odrv4 I__3329 (
            .O(N__26565),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    CascadeMux I__3328 (
            .O(N__26562),
            .I(N__26558));
    CascadeMux I__3327 (
            .O(N__26561),
            .I(N__26555));
    InMux I__3326 (
            .O(N__26558),
            .I(N__26552));
    InMux I__3325 (
            .O(N__26555),
            .I(N__26549));
    LocalMux I__3324 (
            .O(N__26552),
            .I(N__26546));
    LocalMux I__3323 (
            .O(N__26549),
            .I(N__26543));
    Odrv4 I__3322 (
            .O(N__26546),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    Odrv4 I__3321 (
            .O(N__26543),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    InMux I__3320 (
            .O(N__26538),
            .I(N__26535));
    LocalMux I__3319 (
            .O(N__26535),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ));
    CascadeMux I__3318 (
            .O(N__26532),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ));
    InMux I__3317 (
            .O(N__26529),
            .I(N__26526));
    LocalMux I__3316 (
            .O(N__26526),
            .I(N__26521));
    InMux I__3315 (
            .O(N__26525),
            .I(N__26516));
    InMux I__3314 (
            .O(N__26524),
            .I(N__26516));
    Span4Mux_v I__3313 (
            .O(N__26521),
            .I(N__26511));
    LocalMux I__3312 (
            .O(N__26516),
            .I(N__26511));
    Odrv4 I__3311 (
            .O(N__26511),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    InMux I__3310 (
            .O(N__26508),
            .I(N__26502));
    InMux I__3309 (
            .O(N__26507),
            .I(N__26502));
    LocalMux I__3308 (
            .O(N__26502),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ));
    InMux I__3307 (
            .O(N__26499),
            .I(N__26493));
    InMux I__3306 (
            .O(N__26498),
            .I(N__26493));
    LocalMux I__3305 (
            .O(N__26493),
            .I(N__26490));
    Span4Mux_v I__3304 (
            .O(N__26490),
            .I(N__26487));
    Span4Mux_h I__3303 (
            .O(N__26487),
            .I(N__26484));
    Odrv4 I__3302 (
            .O(N__26484),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    InMux I__3301 (
            .O(N__26481),
            .I(N__26475));
    InMux I__3300 (
            .O(N__26480),
            .I(N__26475));
    LocalMux I__3299 (
            .O(N__26475),
            .I(N__26472));
    Span4Mux_v I__3298 (
            .O(N__26472),
            .I(N__26469));
    Odrv4 I__3297 (
            .O(N__26469),
            .I(\pid_alt.error_d_reg_prevZ0Z_14 ));
    InMux I__3296 (
            .O(N__26466),
            .I(N__26463));
    LocalMux I__3295 (
            .O(N__26463),
            .I(N__26458));
    InMux I__3294 (
            .O(N__26462),
            .I(N__26455));
    InMux I__3293 (
            .O(N__26461),
            .I(N__26452));
    Sp12to4 I__3292 (
            .O(N__26458),
            .I(N__26445));
    LocalMux I__3291 (
            .O(N__26455),
            .I(N__26445));
    LocalMux I__3290 (
            .O(N__26452),
            .I(N__26445));
    Span12Mux_v I__3289 (
            .O(N__26445),
            .I(N__26442));
    Odrv12 I__3288 (
            .O(N__26442),
            .I(\pid_alt.error_d_regZ0Z_14 ));
    InMux I__3287 (
            .O(N__26439),
            .I(N__26435));
    CascadeMux I__3286 (
            .O(N__26438),
            .I(N__26432));
    LocalMux I__3285 (
            .O(N__26435),
            .I(N__26429));
    InMux I__3284 (
            .O(N__26432),
            .I(N__26426));
    Odrv4 I__3283 (
            .O(N__26429),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    LocalMux I__3282 (
            .O(N__26426),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    CascadeMux I__3281 (
            .O(N__26421),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ));
    InMux I__3280 (
            .O(N__26418),
            .I(N__26415));
    LocalMux I__3279 (
            .O(N__26415),
            .I(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ));
    InMux I__3278 (
            .O(N__26412),
            .I(N__26409));
    LocalMux I__3277 (
            .O(N__26409),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ));
    InMux I__3276 (
            .O(N__26406),
            .I(N__26400));
    InMux I__3275 (
            .O(N__26405),
            .I(N__26400));
    LocalMux I__3274 (
            .O(N__26400),
            .I(N__26397));
    Span4Mux_v I__3273 (
            .O(N__26397),
            .I(N__26394));
    Odrv4 I__3272 (
            .O(N__26394),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ));
    InMux I__3271 (
            .O(N__26391),
            .I(N__26388));
    LocalMux I__3270 (
            .O(N__26388),
            .I(N__26383));
    InMux I__3269 (
            .O(N__26387),
            .I(N__26378));
    InMux I__3268 (
            .O(N__26386),
            .I(N__26378));
    Span4Mux_v I__3267 (
            .O(N__26383),
            .I(N__26373));
    LocalMux I__3266 (
            .O(N__26378),
            .I(N__26373));
    Odrv4 I__3265 (
            .O(N__26373),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    CascadeMux I__3264 (
            .O(N__26370),
            .I(N__26367));
    InMux I__3263 (
            .O(N__26367),
            .I(N__26363));
    CascadeMux I__3262 (
            .O(N__26366),
            .I(N__26360));
    LocalMux I__3261 (
            .O(N__26363),
            .I(N__26357));
    InMux I__3260 (
            .O(N__26360),
            .I(N__26354));
    Span4Mux_h I__3259 (
            .O(N__26357),
            .I(N__26351));
    LocalMux I__3258 (
            .O(N__26354),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    Odrv4 I__3257 (
            .O(N__26351),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    InMux I__3256 (
            .O(N__26346),
            .I(N__26343));
    LocalMux I__3255 (
            .O(N__26343),
            .I(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ));
    InMux I__3254 (
            .O(N__26340),
            .I(N__26337));
    LocalMux I__3253 (
            .O(N__26337),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ));
    CascadeMux I__3252 (
            .O(N__26334),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ));
    InMux I__3251 (
            .O(N__26331),
            .I(N__26327));
    CascadeMux I__3250 (
            .O(N__26330),
            .I(N__26324));
    LocalMux I__3249 (
            .O(N__26327),
            .I(N__26321));
    InMux I__3248 (
            .O(N__26324),
            .I(N__26318));
    Odrv4 I__3247 (
            .O(N__26321),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    LocalMux I__3246 (
            .O(N__26318),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    InMux I__3245 (
            .O(N__26313),
            .I(N__26310));
    LocalMux I__3244 (
            .O(N__26310),
            .I(N__26306));
    InMux I__3243 (
            .O(N__26309),
            .I(N__26303));
    Span4Mux_v I__3242 (
            .O(N__26306),
            .I(N__26300));
    LocalMux I__3241 (
            .O(N__26303),
            .I(N__26297));
    Span4Mux_h I__3240 (
            .O(N__26300),
            .I(N__26294));
    Span4Mux_v I__3239 (
            .O(N__26297),
            .I(N__26291));
    Odrv4 I__3238 (
            .O(N__26294),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    Odrv4 I__3237 (
            .O(N__26291),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    InMux I__3236 (
            .O(N__26286),
            .I(N__26283));
    LocalMux I__3235 (
            .O(N__26283),
            .I(N__26279));
    InMux I__3234 (
            .O(N__26282),
            .I(N__26276));
    Odrv12 I__3233 (
            .O(N__26279),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    LocalMux I__3232 (
            .O(N__26276),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    InMux I__3231 (
            .O(N__26271),
            .I(N__26266));
    InMux I__3230 (
            .O(N__26270),
            .I(N__26261));
    InMux I__3229 (
            .O(N__26269),
            .I(N__26261));
    LocalMux I__3228 (
            .O(N__26266),
            .I(N__26258));
    LocalMux I__3227 (
            .O(N__26261),
            .I(N__26255));
    Span4Mux_v I__3226 (
            .O(N__26258),
            .I(N__26252));
    Span4Mux_v I__3225 (
            .O(N__26255),
            .I(N__26249));
    Span4Mux_v I__3224 (
            .O(N__26252),
            .I(N__26246));
    Span4Mux_v I__3223 (
            .O(N__26249),
            .I(N__26243));
    Span4Mux_v I__3222 (
            .O(N__26246),
            .I(N__26240));
    Span4Mux_v I__3221 (
            .O(N__26243),
            .I(N__26237));
    Odrv4 I__3220 (
            .O(N__26240),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    Odrv4 I__3219 (
            .O(N__26237),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    InMux I__3218 (
            .O(N__26232),
            .I(N__26229));
    LocalMux I__3217 (
            .O(N__26229),
            .I(N__26226));
    Odrv4 I__3216 (
            .O(N__26226),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    CascadeMux I__3215 (
            .O(N__26223),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_ ));
    InMux I__3214 (
            .O(N__26220),
            .I(N__26217));
    LocalMux I__3213 (
            .O(N__26217),
            .I(N__26214));
    Odrv4 I__3212 (
            .O(N__26214),
            .I(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ));
    InMux I__3211 (
            .O(N__26211),
            .I(N__26207));
    InMux I__3210 (
            .O(N__26210),
            .I(N__26204));
    LocalMux I__3209 (
            .O(N__26207),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ));
    LocalMux I__3208 (
            .O(N__26204),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ));
    InMux I__3207 (
            .O(N__26199),
            .I(N__26196));
    LocalMux I__3206 (
            .O(N__26196),
            .I(N__26193));
    Span12Mux_s4_h I__3205 (
            .O(N__26193),
            .I(N__26190));
    Odrv12 I__3204 (
            .O(N__26190),
            .I(drone_altitude_i_11));
    CascadeMux I__3203 (
            .O(N__26187),
            .I(N__26184));
    InMux I__3202 (
            .O(N__26184),
            .I(N__26180));
    InMux I__3201 (
            .O(N__26183),
            .I(N__26177));
    LocalMux I__3200 (
            .O(N__26180),
            .I(N__26174));
    LocalMux I__3199 (
            .O(N__26177),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    Odrv4 I__3198 (
            .O(N__26174),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    InMux I__3197 (
            .O(N__26169),
            .I(N__26164));
    InMux I__3196 (
            .O(N__26168),
            .I(N__26159));
    InMux I__3195 (
            .O(N__26167),
            .I(N__26159));
    LocalMux I__3194 (
            .O(N__26164),
            .I(N__26154));
    LocalMux I__3193 (
            .O(N__26159),
            .I(N__26154));
    Span4Mux_v I__3192 (
            .O(N__26154),
            .I(N__26151));
    Odrv4 I__3191 (
            .O(N__26151),
            .I(\pid_alt.error_d_regZ0Z_9 ));
    CascadeMux I__3190 (
            .O(N__26148),
            .I(N__26145));
    InMux I__3189 (
            .O(N__26145),
            .I(N__26139));
    InMux I__3188 (
            .O(N__26144),
            .I(N__26139));
    LocalMux I__3187 (
            .O(N__26139),
            .I(N__26136));
    Odrv4 I__3186 (
            .O(N__26136),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    InMux I__3185 (
            .O(N__26133),
            .I(N__26127));
    InMux I__3184 (
            .O(N__26132),
            .I(N__26127));
    LocalMux I__3183 (
            .O(N__26127),
            .I(N__26124));
    Span4Mux_h I__3182 (
            .O(N__26124),
            .I(N__26121));
    Span4Mux_v I__3181 (
            .O(N__26121),
            .I(N__26118));
    Odrv4 I__3180 (
            .O(N__26118),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    InMux I__3179 (
            .O(N__26115),
            .I(N__26112));
    LocalMux I__3178 (
            .O(N__26112),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ));
    InMux I__3177 (
            .O(N__26109),
            .I(N__26103));
    InMux I__3176 (
            .O(N__26108),
            .I(N__26103));
    LocalMux I__3175 (
            .O(N__26103),
            .I(N__26100));
    Span4Mux_v I__3174 (
            .O(N__26100),
            .I(N__26097));
    Odrv4 I__3173 (
            .O(N__26097),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ));
    CascadeMux I__3172 (
            .O(N__26094),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ));
    InMux I__3171 (
            .O(N__26091),
            .I(N__26088));
    LocalMux I__3170 (
            .O(N__26088),
            .I(N__26085));
    Odrv4 I__3169 (
            .O(N__26085),
            .I(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ));
    InMux I__3168 (
            .O(N__26082),
            .I(N__26079));
    LocalMux I__3167 (
            .O(N__26079),
            .I(N__26076));
    Span4Mux_v I__3166 (
            .O(N__26076),
            .I(N__26073));
    Odrv4 I__3165 (
            .O(N__26073),
            .I(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ));
    CascadeMux I__3164 (
            .O(N__26070),
            .I(N__26067));
    InMux I__3163 (
            .O(N__26067),
            .I(N__26063));
    InMux I__3162 (
            .O(N__26066),
            .I(N__26060));
    LocalMux I__3161 (
            .O(N__26063),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    LocalMux I__3160 (
            .O(N__26060),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    CascadeMux I__3159 (
            .O(N__26055),
            .I(N__26052));
    InMux I__3158 (
            .O(N__26052),
            .I(N__26048));
    InMux I__3157 (
            .O(N__26051),
            .I(N__26045));
    LocalMux I__3156 (
            .O(N__26048),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    LocalMux I__3155 (
            .O(N__26045),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    InMux I__3154 (
            .O(N__26040),
            .I(N__26036));
    InMux I__3153 (
            .O(N__26039),
            .I(N__26033));
    LocalMux I__3152 (
            .O(N__26036),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    LocalMux I__3151 (
            .O(N__26033),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    CascadeMux I__3150 (
            .O(N__26028),
            .I(N__26025));
    InMux I__3149 (
            .O(N__26025),
            .I(N__26021));
    InMux I__3148 (
            .O(N__26024),
            .I(N__26018));
    LocalMux I__3147 (
            .O(N__26021),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    LocalMux I__3146 (
            .O(N__26018),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    CascadeMux I__3145 (
            .O(N__26013),
            .I(N__26010));
    InMux I__3144 (
            .O(N__26010),
            .I(N__26006));
    InMux I__3143 (
            .O(N__26009),
            .I(N__26003));
    LocalMux I__3142 (
            .O(N__26006),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    LocalMux I__3141 (
            .O(N__26003),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    InMux I__3140 (
            .O(N__25998),
            .I(N__25994));
    InMux I__3139 (
            .O(N__25997),
            .I(N__25991));
    LocalMux I__3138 (
            .O(N__25994),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    LocalMux I__3137 (
            .O(N__25991),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    InMux I__3136 (
            .O(N__25986),
            .I(N__25983));
    LocalMux I__3135 (
            .O(N__25983),
            .I(N__25980));
    Odrv4 I__3134 (
            .O(N__25980),
            .I(\pid_alt.m35_e_2 ));
    CascadeMux I__3133 (
            .O(N__25977),
            .I(N__25974));
    InMux I__3132 (
            .O(N__25974),
            .I(N__25970));
    InMux I__3131 (
            .O(N__25973),
            .I(N__25967));
    LocalMux I__3130 (
            .O(N__25970),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    LocalMux I__3129 (
            .O(N__25967),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    InMux I__3128 (
            .O(N__25962),
            .I(N__25959));
    LocalMux I__3127 (
            .O(N__25959),
            .I(N__25956));
    Span4Mux_v I__3126 (
            .O(N__25956),
            .I(N__25953));
    Odrv4 I__3125 (
            .O(N__25953),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ));
    InMux I__3124 (
            .O(N__25950),
            .I(N__25947));
    LocalMux I__3123 (
            .O(N__25947),
            .I(N__25943));
    InMux I__3122 (
            .O(N__25946),
            .I(N__25940));
    Span4Mux_v I__3121 (
            .O(N__25943),
            .I(N__25937));
    LocalMux I__3120 (
            .O(N__25940),
            .I(N__25934));
    Span4Mux_h I__3119 (
            .O(N__25937),
            .I(N__25931));
    Span4Mux_v I__3118 (
            .O(N__25934),
            .I(N__25928));
    Odrv4 I__3117 (
            .O(N__25931),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ));
    Odrv4 I__3116 (
            .O(N__25928),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ));
    InMux I__3115 (
            .O(N__25923),
            .I(N__25919));
    InMux I__3114 (
            .O(N__25922),
            .I(N__25915));
    LocalMux I__3113 (
            .O(N__25919),
            .I(N__25912));
    InMux I__3112 (
            .O(N__25918),
            .I(N__25909));
    LocalMux I__3111 (
            .O(N__25915),
            .I(N__25906));
    Odrv4 I__3110 (
            .O(N__25912),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    LocalMux I__3109 (
            .O(N__25909),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    Odrv4 I__3108 (
            .O(N__25906),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    CascadeMux I__3107 (
            .O(N__25899),
            .I(N__25895));
    CascadeMux I__3106 (
            .O(N__25898),
            .I(N__25892));
    InMux I__3105 (
            .O(N__25895),
            .I(N__25889));
    InMux I__3104 (
            .O(N__25892),
            .I(N__25886));
    LocalMux I__3103 (
            .O(N__25889),
            .I(N__25883));
    LocalMux I__3102 (
            .O(N__25886),
            .I(N__25880));
    Span4Mux_v I__3101 (
            .O(N__25883),
            .I(N__25877));
    Span4Mux_h I__3100 (
            .O(N__25880),
            .I(N__25874));
    Odrv4 I__3099 (
            .O(N__25877),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ));
    Odrv4 I__3098 (
            .O(N__25874),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ));
    InMux I__3097 (
            .O(N__25869),
            .I(N__25865));
    CascadeMux I__3096 (
            .O(N__25868),
            .I(N__25862));
    LocalMux I__3095 (
            .O(N__25865),
            .I(N__25858));
    InMux I__3094 (
            .O(N__25862),
            .I(N__25855));
    InMux I__3093 (
            .O(N__25861),
            .I(N__25852));
    Span12Mux_s3_h I__3092 (
            .O(N__25858),
            .I(N__25847));
    LocalMux I__3091 (
            .O(N__25855),
            .I(N__25847));
    LocalMux I__3090 (
            .O(N__25852),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    Odrv12 I__3089 (
            .O(N__25847),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    InMux I__3088 (
            .O(N__25842),
            .I(N__25839));
    LocalMux I__3087 (
            .O(N__25839),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    CascadeMux I__3086 (
            .O(N__25836),
            .I(N__25833));
    InMux I__3085 (
            .O(N__25833),
            .I(N__25830));
    LocalMux I__3084 (
            .O(N__25830),
            .I(N__25827));
    Odrv4 I__3083 (
            .O(N__25827),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    CascadeMux I__3082 (
            .O(N__25824),
            .I(\pid_alt.N_9_0_cascade_ ));
    CascadeMux I__3081 (
            .O(N__25821),
            .I(\pid_alt.N_62_mux_cascade_ ));
    InMux I__3080 (
            .O(N__25818),
            .I(N__25815));
    LocalMux I__3079 (
            .O(N__25815),
            .I(N__25811));
    InMux I__3078 (
            .O(N__25814),
            .I(N__25808));
    Odrv4 I__3077 (
            .O(N__25811),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    LocalMux I__3076 (
            .O(N__25808),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    InMux I__3075 (
            .O(N__25803),
            .I(N__25800));
    LocalMux I__3074 (
            .O(N__25800),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    CascadeMux I__3073 (
            .O(N__25797),
            .I(N__25793));
    CascadeMux I__3072 (
            .O(N__25796),
            .I(N__25789));
    InMux I__3071 (
            .O(N__25793),
            .I(N__25779));
    InMux I__3070 (
            .O(N__25792),
            .I(N__25779));
    InMux I__3069 (
            .O(N__25789),
            .I(N__25779));
    InMux I__3068 (
            .O(N__25788),
            .I(N__25779));
    LocalMux I__3067 (
            .O(N__25779),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNIEPGB3Z0Z_5 ));
    InMux I__3066 (
            .O(N__25776),
            .I(N__25773));
    LocalMux I__3065 (
            .O(N__25773),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    InMux I__3064 (
            .O(N__25770),
            .I(N__25767));
    LocalMux I__3063 (
            .O(N__25767),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    InMux I__3062 (
            .O(N__25764),
            .I(N__25761));
    LocalMux I__3061 (
            .O(N__25761),
            .I(\pid_alt.error_i_acumm_preregZ0Z_17 ));
    InMux I__3060 (
            .O(N__25758),
            .I(N__25755));
    LocalMux I__3059 (
            .O(N__25755),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    InMux I__3058 (
            .O(N__25752),
            .I(N__25749));
    LocalMux I__3057 (
            .O(N__25749),
            .I(\pid_alt.error_i_acumm_preregZ0Z_15 ));
    InMux I__3056 (
            .O(N__25746),
            .I(N__25741));
    InMux I__3055 (
            .O(N__25745),
            .I(N__25736));
    InMux I__3054 (
            .O(N__25744),
            .I(N__25736));
    LocalMux I__3053 (
            .O(N__25741),
            .I(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ));
    LocalMux I__3052 (
            .O(N__25736),
            .I(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ));
    CascadeMux I__3051 (
            .O(N__25731),
            .I(N__25728));
    InMux I__3050 (
            .O(N__25728),
            .I(N__25723));
    InMux I__3049 (
            .O(N__25727),
            .I(N__25720));
    InMux I__3048 (
            .O(N__25726),
            .I(N__25717));
    LocalMux I__3047 (
            .O(N__25723),
            .I(N__25714));
    LocalMux I__3046 (
            .O(N__25720),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    LocalMux I__3045 (
            .O(N__25717),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    Odrv4 I__3044 (
            .O(N__25714),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    InMux I__3043 (
            .O(N__25707),
            .I(N__25702));
    InMux I__3042 (
            .O(N__25706),
            .I(N__25697));
    InMux I__3041 (
            .O(N__25705),
            .I(N__25697));
    LocalMux I__3040 (
            .O(N__25702),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    LocalMux I__3039 (
            .O(N__25697),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    InMux I__3038 (
            .O(N__25692),
            .I(N__25689));
    LocalMux I__3037 (
            .O(N__25689),
            .I(N__25686));
    Span4Mux_v I__3036 (
            .O(N__25686),
            .I(N__25683));
    Odrv4 I__3035 (
            .O(N__25683),
            .I(alt_kp_2));
    InMux I__3034 (
            .O(N__25680),
            .I(N__25677));
    LocalMux I__3033 (
            .O(N__25677),
            .I(N__25674));
    Span4Mux_s3_h I__3032 (
            .O(N__25674),
            .I(N__25671));
    Odrv4 I__3031 (
            .O(N__25671),
            .I(alt_kp_5));
    InMux I__3030 (
            .O(N__25668),
            .I(N__25664));
    CascadeMux I__3029 (
            .O(N__25667),
            .I(N__25661));
    LocalMux I__3028 (
            .O(N__25664),
            .I(N__25658));
    InMux I__3027 (
            .O(N__25661),
            .I(N__25655));
    Span4Mux_h I__3026 (
            .O(N__25658),
            .I(N__25652));
    LocalMux I__3025 (
            .O(N__25655),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    Odrv4 I__3024 (
            .O(N__25652),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    CascadeMux I__3023 (
            .O(N__25647),
            .I(N__25644));
    InMux I__3022 (
            .O(N__25644),
            .I(N__25640));
    InMux I__3021 (
            .O(N__25643),
            .I(N__25637));
    LocalMux I__3020 (
            .O(N__25640),
            .I(N__25634));
    LocalMux I__3019 (
            .O(N__25637),
            .I(N__25631));
    Span4Mux_v I__3018 (
            .O(N__25634),
            .I(N__25628));
    Odrv4 I__3017 (
            .O(N__25631),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    Odrv4 I__3016 (
            .O(N__25628),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    InMux I__3015 (
            .O(N__25623),
            .I(N__25620));
    LocalMux I__3014 (
            .O(N__25620),
            .I(\pid_alt.error_i_acumm_preregZ0Z_18 ));
    CascadeMux I__3013 (
            .O(N__25617),
            .I(N__25614));
    InMux I__3012 (
            .O(N__25614),
            .I(N__25611));
    LocalMux I__3011 (
            .O(N__25611),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    InMux I__3010 (
            .O(N__25608),
            .I(N__25605));
    LocalMux I__3009 (
            .O(N__25605),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    CascadeMux I__3008 (
            .O(N__25602),
            .I(\pid_alt.m7_e_4_cascade_ ));
    InMux I__3007 (
            .O(N__25599),
            .I(N__25595));
    InMux I__3006 (
            .O(N__25598),
            .I(N__25592));
    LocalMux I__3005 (
            .O(N__25595),
            .I(N__25589));
    LocalMux I__3004 (
            .O(N__25592),
            .I(N__25586));
    Span4Mux_h I__3003 (
            .O(N__25589),
            .I(N__25583));
    Span4Mux_v I__3002 (
            .O(N__25586),
            .I(N__25580));
    Odrv4 I__3001 (
            .O(N__25583),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    Odrv4 I__3000 (
            .O(N__25580),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    InMux I__2999 (
            .O(N__25575),
            .I(N__25569));
    InMux I__2998 (
            .O(N__25574),
            .I(N__25569));
    LocalMux I__2997 (
            .O(N__25569),
            .I(N__25566));
    Span4Mux_h I__2996 (
            .O(N__25566),
            .I(N__25562));
    InMux I__2995 (
            .O(N__25565),
            .I(N__25559));
    Span4Mux_v I__2994 (
            .O(N__25562),
            .I(N__25556));
    LocalMux I__2993 (
            .O(N__25559),
            .I(N__25553));
    Sp12to4 I__2992 (
            .O(N__25556),
            .I(N__25548));
    Span12Mux_s5_h I__2991 (
            .O(N__25553),
            .I(N__25548));
    Span12Mux_v I__2990 (
            .O(N__25548),
            .I(N__25545));
    Odrv12 I__2989 (
            .O(N__25545),
            .I(\pid_alt.error_d_regZ0Z_13 ));
    InMux I__2988 (
            .O(N__25542),
            .I(N__25539));
    LocalMux I__2987 (
            .O(N__25539),
            .I(N__25535));
    InMux I__2986 (
            .O(N__25538),
            .I(N__25532));
    Span4Mux_s3_h I__2985 (
            .O(N__25535),
            .I(N__25529));
    LocalMux I__2984 (
            .O(N__25532),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    Odrv4 I__2983 (
            .O(N__25529),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    InMux I__2982 (
            .O(N__25524),
            .I(N__25521));
    LocalMux I__2981 (
            .O(N__25521),
            .I(N__25518));
    Odrv4 I__2980 (
            .O(N__25518),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20 ));
    CascadeMux I__2979 (
            .O(N__25515),
            .I(N__25512));
    InMux I__2978 (
            .O(N__25512),
            .I(N__25509));
    LocalMux I__2977 (
            .O(N__25509),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20 ));
    CascadeMux I__2976 (
            .O(N__25506),
            .I(N__25503));
    InMux I__2975 (
            .O(N__25503),
            .I(N__25499));
    InMux I__2974 (
            .O(N__25502),
            .I(N__25496));
    LocalMux I__2973 (
            .O(N__25499),
            .I(N__25493));
    LocalMux I__2972 (
            .O(N__25496),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ));
    Odrv4 I__2971 (
            .O(N__25493),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ));
    InMux I__2970 (
            .O(N__25488),
            .I(N__25485));
    LocalMux I__2969 (
            .O(N__25485),
            .I(\dron_frame_decoder_1.drone_altitude_10 ));
    InMux I__2968 (
            .O(N__25482),
            .I(\pid_alt.un1_pid_prereg_0_cry_15 ));
    InMux I__2967 (
            .O(N__25479),
            .I(\pid_alt.un1_pid_prereg_0_cry_16 ));
    InMux I__2966 (
            .O(N__25476),
            .I(N__25473));
    LocalMux I__2965 (
            .O(N__25473),
            .I(N__25470));
    Odrv4 I__2964 (
            .O(N__25470),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ));
    InMux I__2963 (
            .O(N__25467),
            .I(\pid_alt.un1_pid_prereg_0_cry_17 ));
    InMux I__2962 (
            .O(N__25464),
            .I(N__25461));
    LocalMux I__2961 (
            .O(N__25461),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ));
    CascadeMux I__2960 (
            .O(N__25458),
            .I(N__25454));
    CascadeMux I__2959 (
            .O(N__25457),
            .I(N__25451));
    InMux I__2958 (
            .O(N__25454),
            .I(N__25448));
    InMux I__2957 (
            .O(N__25451),
            .I(N__25445));
    LocalMux I__2956 (
            .O(N__25448),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    LocalMux I__2955 (
            .O(N__25445),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    InMux I__2954 (
            .O(N__25440),
            .I(\pid_alt.un1_pid_prereg_0_cry_18 ));
    InMux I__2953 (
            .O(N__25437),
            .I(\pid_alt.un1_pid_prereg_0_cry_19 ));
    InMux I__2952 (
            .O(N__25434),
            .I(\pid_alt.un1_pid_prereg_0_cry_20 ));
    InMux I__2951 (
            .O(N__25431),
            .I(\pid_alt.un1_pid_prereg_0_cry_21 ));
    InMux I__2950 (
            .O(N__25428),
            .I(bfn_3_20_0_));
    InMux I__2949 (
            .O(N__25425),
            .I(\pid_alt.un1_pid_prereg_0_cry_23 ));
    InMux I__2948 (
            .O(N__25422),
            .I(bfn_3_18_0_));
    InMux I__2947 (
            .O(N__25419),
            .I(\pid_alt.un1_pid_prereg_0_cry_7 ));
    InMux I__2946 (
            .O(N__25416),
            .I(\pid_alt.un1_pid_prereg_0_cry_8 ));
    InMux I__2945 (
            .O(N__25413),
            .I(\pid_alt.un1_pid_prereg_0_cry_9 ));
    InMux I__2944 (
            .O(N__25410),
            .I(N__25407));
    LocalMux I__2943 (
            .O(N__25407),
            .I(N__25404));
    Odrv4 I__2942 (
            .O(N__25404),
            .I(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ));
    CascadeMux I__2941 (
            .O(N__25401),
            .I(N__25397));
    CascadeMux I__2940 (
            .O(N__25400),
            .I(N__25394));
    InMux I__2939 (
            .O(N__25397),
            .I(N__25391));
    InMux I__2938 (
            .O(N__25394),
            .I(N__25388));
    LocalMux I__2937 (
            .O(N__25391),
            .I(N__25385));
    LocalMux I__2936 (
            .O(N__25388),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    Odrv4 I__2935 (
            .O(N__25385),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    InMux I__2934 (
            .O(N__25380),
            .I(\pid_alt.un1_pid_prereg_0_cry_10 ));
    InMux I__2933 (
            .O(N__25377),
            .I(N__25374));
    LocalMux I__2932 (
            .O(N__25374),
            .I(\pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ));
    CascadeMux I__2931 (
            .O(N__25371),
            .I(N__25368));
    InMux I__2930 (
            .O(N__25368),
            .I(N__25364));
    InMux I__2929 (
            .O(N__25367),
            .I(N__25361));
    LocalMux I__2928 (
            .O(N__25364),
            .I(N__25358));
    LocalMux I__2927 (
            .O(N__25361),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ));
    Odrv4 I__2926 (
            .O(N__25358),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ));
    InMux I__2925 (
            .O(N__25353),
            .I(\pid_alt.un1_pid_prereg_0_cry_11 ));
    InMux I__2924 (
            .O(N__25350),
            .I(N__25347));
    LocalMux I__2923 (
            .O(N__25347),
            .I(\pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ));
    InMux I__2922 (
            .O(N__25344),
            .I(\pid_alt.un1_pid_prereg_0_cry_12 ));
    InMux I__2921 (
            .O(N__25341),
            .I(\pid_alt.un1_pid_prereg_0_cry_13 ));
    InMux I__2920 (
            .O(N__25338),
            .I(bfn_3_19_0_));
    InMux I__2919 (
            .O(N__25335),
            .I(N__25332));
    LocalMux I__2918 (
            .O(N__25332),
            .I(N__25329));
    Odrv4 I__2917 (
            .O(N__25329),
            .I(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ));
    CascadeMux I__2916 (
            .O(N__25326),
            .I(N__25323));
    InMux I__2915 (
            .O(N__25323),
            .I(N__25320));
    LocalMux I__2914 (
            .O(N__25320),
            .I(N__25316));
    InMux I__2913 (
            .O(N__25319),
            .I(N__25313));
    Span4Mux_v I__2912 (
            .O(N__25316),
            .I(N__25310));
    LocalMux I__2911 (
            .O(N__25313),
            .I(\pid_alt.un1_pid_prereg_0 ));
    Odrv4 I__2910 (
            .O(N__25310),
            .I(\pid_alt.un1_pid_prereg_0 ));
    InMux I__2909 (
            .O(N__25305),
            .I(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__2908 (
            .O(N__25302),
            .I(N__25299));
    LocalMux I__2907 (
            .O(N__25299),
            .I(N__25296));
    Span4Mux_v I__2906 (
            .O(N__25296),
            .I(N__25293));
    Odrv4 I__2905 (
            .O(N__25293),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1 ));
    CascadeMux I__2904 (
            .O(N__25290),
            .I(N__25286));
    InMux I__2903 (
            .O(N__25289),
            .I(N__25283));
    InMux I__2902 (
            .O(N__25286),
            .I(N__25280));
    LocalMux I__2901 (
            .O(N__25283),
            .I(N__25275));
    LocalMux I__2900 (
            .O(N__25280),
            .I(N__25275));
    Odrv12 I__2899 (
            .O(N__25275),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    InMux I__2898 (
            .O(N__25272),
            .I(\pid_alt.un1_pid_prereg_0_cry_0 ));
    InMux I__2897 (
            .O(N__25269),
            .I(N__25266));
    LocalMux I__2896 (
            .O(N__25266),
            .I(N__25263));
    Odrv4 I__2895 (
            .O(N__25263),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1 ));
    InMux I__2894 (
            .O(N__25260),
            .I(\pid_alt.un1_pid_prereg_0_cry_1 ));
    InMux I__2893 (
            .O(N__25257),
            .I(N__25254));
    LocalMux I__2892 (
            .O(N__25254),
            .I(N__25251));
    Span4Mux_v I__2891 (
            .O(N__25251),
            .I(N__25248));
    Odrv4 I__2890 (
            .O(N__25248),
            .I(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ));
    InMux I__2889 (
            .O(N__25245),
            .I(\pid_alt.un1_pid_prereg_0_cry_2 ));
    CascadeMux I__2888 (
            .O(N__25242),
            .I(N__25239));
    InMux I__2887 (
            .O(N__25239),
            .I(N__25235));
    InMux I__2886 (
            .O(N__25238),
            .I(N__25232));
    LocalMux I__2885 (
            .O(N__25235),
            .I(N__25229));
    LocalMux I__2884 (
            .O(N__25232),
            .I(N__25226));
    Span4Mux_v I__2883 (
            .O(N__25229),
            .I(N__25221));
    Span4Mux_v I__2882 (
            .O(N__25226),
            .I(N__25221));
    Odrv4 I__2881 (
            .O(N__25221),
            .I(\pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3 ));
    CascadeMux I__2880 (
            .O(N__25218),
            .I(N__25215));
    InMux I__2879 (
            .O(N__25215),
            .I(N__25212));
    LocalMux I__2878 (
            .O(N__25212),
            .I(N__25209));
    Odrv12 I__2877 (
            .O(N__25209),
            .I(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ));
    InMux I__2876 (
            .O(N__25206),
            .I(\pid_alt.un1_pid_prereg_0_cry_3 ));
    InMux I__2875 (
            .O(N__25203),
            .I(N__25200));
    LocalMux I__2874 (
            .O(N__25200),
            .I(N__25197));
    Odrv12 I__2873 (
            .O(N__25197),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ));
    CascadeMux I__2872 (
            .O(N__25194),
            .I(N__25191));
    InMux I__2871 (
            .O(N__25191),
            .I(N__25188));
    LocalMux I__2870 (
            .O(N__25188),
            .I(N__25184));
    InMux I__2869 (
            .O(N__25187),
            .I(N__25181));
    Span4Mux_v I__2868 (
            .O(N__25184),
            .I(N__25178));
    LocalMux I__2867 (
            .O(N__25181),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    Odrv4 I__2866 (
            .O(N__25178),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    InMux I__2865 (
            .O(N__25173),
            .I(\pid_alt.un1_pid_prereg_0_cry_4 ));
    InMux I__2864 (
            .O(N__25170),
            .I(N__25167));
    LocalMux I__2863 (
            .O(N__25167),
            .I(N__25164));
    Span4Mux_v I__2862 (
            .O(N__25164),
            .I(N__25161));
    Odrv4 I__2861 (
            .O(N__25161),
            .I(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ));
    CascadeMux I__2860 (
            .O(N__25158),
            .I(N__25154));
    CascadeMux I__2859 (
            .O(N__25157),
            .I(N__25151));
    InMux I__2858 (
            .O(N__25154),
            .I(N__25148));
    InMux I__2857 (
            .O(N__25151),
            .I(N__25145));
    LocalMux I__2856 (
            .O(N__25148),
            .I(N__25142));
    LocalMux I__2855 (
            .O(N__25145),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    Odrv12 I__2854 (
            .O(N__25142),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    InMux I__2853 (
            .O(N__25137),
            .I(\pid_alt.un1_pid_prereg_0_cry_5 ));
    InMux I__2852 (
            .O(N__25134),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__2851 (
            .O(N__25131),
            .I(N__25128));
    LocalMux I__2850 (
            .O(N__25128),
            .I(N__25125));
    Span4Mux_v I__2849 (
            .O(N__25125),
            .I(N__25122));
    Span4Mux_v I__2848 (
            .O(N__25122),
            .I(N__25119));
    Odrv4 I__2847 (
            .O(N__25119),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    InMux I__2846 (
            .O(N__25116),
            .I(bfn_3_16_0_));
    InMux I__2845 (
            .O(N__25113),
            .I(N__25110));
    LocalMux I__2844 (
            .O(N__25110),
            .I(N__25107));
    Span4Mux_v I__2843 (
            .O(N__25107),
            .I(N__25104));
    Span4Mux_v I__2842 (
            .O(N__25104),
            .I(N__25101));
    Odrv4 I__2841 (
            .O(N__25101),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    InMux I__2840 (
            .O(N__25098),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__2839 (
            .O(N__25095),
            .I(N__25092));
    LocalMux I__2838 (
            .O(N__25092),
            .I(N__25089));
    Span4Mux_v I__2837 (
            .O(N__25089),
            .I(N__25086));
    Span4Mux_v I__2836 (
            .O(N__25086),
            .I(N__25083));
    Odrv4 I__2835 (
            .O(N__25083),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    InMux I__2834 (
            .O(N__25080),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__2833 (
            .O(N__25077),
            .I(N__25074));
    LocalMux I__2832 (
            .O(N__25074),
            .I(N__25071));
    Span4Mux_v I__2831 (
            .O(N__25071),
            .I(N__25068));
    Span4Mux_v I__2830 (
            .O(N__25068),
            .I(N__25065));
    Odrv4 I__2829 (
            .O(N__25065),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    InMux I__2828 (
            .O(N__25062),
            .I(N__25057));
    InMux I__2827 (
            .O(N__25061),
            .I(N__25052));
    InMux I__2826 (
            .O(N__25060),
            .I(N__25052));
    LocalMux I__2825 (
            .O(N__25057),
            .I(N__25049));
    LocalMux I__2824 (
            .O(N__25052),
            .I(N__25046));
    Span4Mux_h I__2823 (
            .O(N__25049),
            .I(N__25043));
    Span4Mux_v I__2822 (
            .O(N__25046),
            .I(N__25040));
    Odrv4 I__2821 (
            .O(N__25043),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    Odrv4 I__2820 (
            .O(N__25040),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    InMux I__2819 (
            .O(N__25035),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__2818 (
            .O(N__25032),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__2817 (
            .O(N__25029),
            .I(N__25023));
    InMux I__2816 (
            .O(N__25028),
            .I(N__25023));
    LocalMux I__2815 (
            .O(N__25023),
            .I(N__25020));
    Span4Mux_h I__2814 (
            .O(N__25020),
            .I(N__25017));
    Span4Mux_v I__2813 (
            .O(N__25017),
            .I(N__25014));
    Odrv4 I__2812 (
            .O(N__25014),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    InMux I__2811 (
            .O(N__25011),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__2810 (
            .O(N__25008),
            .I(N__25005));
    LocalMux I__2809 (
            .O(N__25005),
            .I(N__25002));
    Span4Mux_h I__2808 (
            .O(N__25002),
            .I(N__24999));
    Odrv4 I__2807 (
            .O(N__24999),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ));
    InMux I__2806 (
            .O(N__24996),
            .I(N__24992));
    InMux I__2805 (
            .O(N__24995),
            .I(N__24989));
    LocalMux I__2804 (
            .O(N__24992),
            .I(N__24986));
    LocalMux I__2803 (
            .O(N__24989),
            .I(N__24982));
    Span4Mux_v I__2802 (
            .O(N__24986),
            .I(N__24979));
    InMux I__2801 (
            .O(N__24985),
            .I(N__24976));
    Odrv12 I__2800 (
            .O(N__24982),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    Odrv4 I__2799 (
            .O(N__24979),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    LocalMux I__2798 (
            .O(N__24976),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    CascadeMux I__2797 (
            .O(N__24969),
            .I(N__24966));
    InMux I__2796 (
            .O(N__24966),
            .I(N__24963));
    LocalMux I__2795 (
            .O(N__24963),
            .I(N__24960));
    Span4Mux_v I__2794 (
            .O(N__24960),
            .I(N__24957));
    Odrv4 I__2793 (
            .O(N__24957),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    InMux I__2792 (
            .O(N__24954),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6 ));
    CascadeMux I__2791 (
            .O(N__24951),
            .I(N__24948));
    InMux I__2790 (
            .O(N__24948),
            .I(N__24945));
    LocalMux I__2789 (
            .O(N__24945),
            .I(N__24942));
    Span4Mux_v I__2788 (
            .O(N__24942),
            .I(N__24939));
    Odrv4 I__2787 (
            .O(N__24939),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    InMux I__2786 (
            .O(N__24936),
            .I(bfn_3_15_0_));
    CascadeMux I__2785 (
            .O(N__24933),
            .I(N__24930));
    InMux I__2784 (
            .O(N__24930),
            .I(N__24927));
    LocalMux I__2783 (
            .O(N__24927),
            .I(N__24924));
    Span4Mux_v I__2782 (
            .O(N__24924),
            .I(N__24921));
    Odrv4 I__2781 (
            .O(N__24921),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    InMux I__2780 (
            .O(N__24918),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8 ));
    CascadeMux I__2779 (
            .O(N__24915),
            .I(N__24912));
    InMux I__2778 (
            .O(N__24912),
            .I(N__24909));
    LocalMux I__2777 (
            .O(N__24909),
            .I(N__24906));
    Span4Mux_v I__2776 (
            .O(N__24906),
            .I(N__24903));
    Span4Mux_v I__2775 (
            .O(N__24903),
            .I(N__24900));
    Odrv4 I__2774 (
            .O(N__24900),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    InMux I__2773 (
            .O(N__24897),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9 ));
    CascadeMux I__2772 (
            .O(N__24894),
            .I(N__24891));
    InMux I__2771 (
            .O(N__24891),
            .I(N__24888));
    LocalMux I__2770 (
            .O(N__24888),
            .I(N__24885));
    Odrv12 I__2769 (
            .O(N__24885),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    InMux I__2768 (
            .O(N__24882),
            .I(N__24873));
    InMux I__2767 (
            .O(N__24881),
            .I(N__24873));
    InMux I__2766 (
            .O(N__24880),
            .I(N__24873));
    LocalMux I__2765 (
            .O(N__24873),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    InMux I__2764 (
            .O(N__24870),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_10 ));
    CascadeMux I__2763 (
            .O(N__24867),
            .I(N__24864));
    InMux I__2762 (
            .O(N__24864),
            .I(N__24861));
    LocalMux I__2761 (
            .O(N__24861),
            .I(N__24858));
    Span4Mux_v I__2760 (
            .O(N__24858),
            .I(N__24855));
    Odrv4 I__2759 (
            .O(N__24855),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    InMux I__2758 (
            .O(N__24852),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_11 ));
    CascadeMux I__2757 (
            .O(N__24849),
            .I(N__24846));
    InMux I__2756 (
            .O(N__24846),
            .I(N__24843));
    LocalMux I__2755 (
            .O(N__24843),
            .I(N__24840));
    Span4Mux_h I__2754 (
            .O(N__24840),
            .I(N__24837));
    Span4Mux_v I__2753 (
            .O(N__24837),
            .I(N__24834));
    Odrv4 I__2752 (
            .O(N__24834),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    InMux I__2751 (
            .O(N__24831),
            .I(N__24826));
    InMux I__2750 (
            .O(N__24830),
            .I(N__24821));
    InMux I__2749 (
            .O(N__24829),
            .I(N__24821));
    LocalMux I__2748 (
            .O(N__24826),
            .I(N__24818));
    LocalMux I__2747 (
            .O(N__24821),
            .I(N__24815));
    Odrv4 I__2746 (
            .O(N__24818),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    Odrv4 I__2745 (
            .O(N__24815),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    InMux I__2744 (
            .O(N__24810),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__2743 (
            .O(N__24807),
            .I(N__24804));
    LocalMux I__2742 (
            .O(N__24804),
            .I(N__24801));
    Span4Mux_v I__2741 (
            .O(N__24801),
            .I(N__24798));
    Odrv4 I__2740 (
            .O(N__24798),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    InMux I__2739 (
            .O(N__24795),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_13 ));
    CascadeMux I__2738 (
            .O(N__24792),
            .I(N__24789));
    InMux I__2737 (
            .O(N__24789),
            .I(N__24786));
    LocalMux I__2736 (
            .O(N__24786),
            .I(N__24783));
    Span4Mux_v I__2735 (
            .O(N__24783),
            .I(N__24780));
    Odrv4 I__2734 (
            .O(N__24780),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    InMux I__2733 (
            .O(N__24777),
            .I(N__24774));
    LocalMux I__2732 (
            .O(N__24774),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ));
    InMux I__2731 (
            .O(N__24771),
            .I(N__24765));
    InMux I__2730 (
            .O(N__24770),
            .I(N__24765));
    LocalMux I__2729 (
            .O(N__24765),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ));
    InMux I__2728 (
            .O(N__24762),
            .I(N__24759));
    LocalMux I__2727 (
            .O(N__24759),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    InMux I__2726 (
            .O(N__24756),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_0 ));
    CascadeMux I__2725 (
            .O(N__24753),
            .I(N__24750));
    InMux I__2724 (
            .O(N__24750),
            .I(N__24747));
    LocalMux I__2723 (
            .O(N__24747),
            .I(N__24744));
    Span4Mux_v I__2722 (
            .O(N__24744),
            .I(N__24741));
    Odrv4 I__2721 (
            .O(N__24741),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    InMux I__2720 (
            .O(N__24738),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_1 ));
    CascadeMux I__2719 (
            .O(N__24735),
            .I(N__24732));
    InMux I__2718 (
            .O(N__24732),
            .I(N__24729));
    LocalMux I__2717 (
            .O(N__24729),
            .I(N__24726));
    Odrv12 I__2716 (
            .O(N__24726),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    InMux I__2715 (
            .O(N__24723),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_2 ));
    CascadeMux I__2714 (
            .O(N__24720),
            .I(N__24717));
    InMux I__2713 (
            .O(N__24717),
            .I(N__24714));
    LocalMux I__2712 (
            .O(N__24714),
            .I(N__24711));
    Span4Mux_h I__2711 (
            .O(N__24711),
            .I(N__24708));
    Span4Mux_v I__2710 (
            .O(N__24708),
            .I(N__24705));
    Odrv4 I__2709 (
            .O(N__24705),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    InMux I__2708 (
            .O(N__24702),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_3 ));
    CascadeMux I__2707 (
            .O(N__24699),
            .I(N__24696));
    InMux I__2706 (
            .O(N__24696),
            .I(N__24693));
    LocalMux I__2705 (
            .O(N__24693),
            .I(N__24690));
    Span4Mux_v I__2704 (
            .O(N__24690),
            .I(N__24687));
    Odrv4 I__2703 (
            .O(N__24687),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    InMux I__2702 (
            .O(N__24684),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_4 ));
    CascadeMux I__2701 (
            .O(N__24681),
            .I(N__24678));
    InMux I__2700 (
            .O(N__24678),
            .I(N__24675));
    LocalMux I__2699 (
            .O(N__24675),
            .I(N__24672));
    Span4Mux_v I__2698 (
            .O(N__24672),
            .I(N__24669));
    Odrv4 I__2697 (
            .O(N__24669),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    InMux I__2696 (
            .O(N__24666),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5 ));
    InMux I__2695 (
            .O(N__24663),
            .I(N__24658));
    InMux I__2694 (
            .O(N__24662),
            .I(N__24655));
    InMux I__2693 (
            .O(N__24661),
            .I(N__24652));
    LocalMux I__2692 (
            .O(N__24658),
            .I(N__24649));
    LocalMux I__2691 (
            .O(N__24655),
            .I(N__24646));
    LocalMux I__2690 (
            .O(N__24652),
            .I(N__24641));
    Span4Mux_h I__2689 (
            .O(N__24649),
            .I(N__24641));
    Span4Mux_v I__2688 (
            .O(N__24646),
            .I(N__24638));
    Span4Mux_v I__2687 (
            .O(N__24641),
            .I(N__24635));
    Span4Mux_v I__2686 (
            .O(N__24638),
            .I(N__24632));
    Odrv4 I__2685 (
            .O(N__24635),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    Odrv4 I__2684 (
            .O(N__24632),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    InMux I__2683 (
            .O(N__24627),
            .I(N__24622));
    InMux I__2682 (
            .O(N__24626),
            .I(N__24619));
    InMux I__2681 (
            .O(N__24625),
            .I(N__24616));
    LocalMux I__2680 (
            .O(N__24622),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    LocalMux I__2679 (
            .O(N__24619),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    LocalMux I__2678 (
            .O(N__24616),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    InMux I__2677 (
            .O(N__24609),
            .I(N__24605));
    InMux I__2676 (
            .O(N__24608),
            .I(N__24601));
    LocalMux I__2675 (
            .O(N__24605),
            .I(N__24597));
    InMux I__2674 (
            .O(N__24604),
            .I(N__24594));
    LocalMux I__2673 (
            .O(N__24601),
            .I(N__24591));
    InMux I__2672 (
            .O(N__24600),
            .I(N__24588));
    Span4Mux_h I__2671 (
            .O(N__24597),
            .I(N__24585));
    LocalMux I__2670 (
            .O(N__24594),
            .I(N__24578));
    Span4Mux_h I__2669 (
            .O(N__24591),
            .I(N__24578));
    LocalMux I__2668 (
            .O(N__24588),
            .I(N__24578));
    Span4Mux_v I__2667 (
            .O(N__24585),
            .I(N__24575));
    Span4Mux_v I__2666 (
            .O(N__24578),
            .I(N__24572));
    Odrv4 I__2665 (
            .O(N__24575),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    Odrv4 I__2664 (
            .O(N__24572),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    InMux I__2663 (
            .O(N__24567),
            .I(N__24564));
    LocalMux I__2662 (
            .O(N__24564),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ));
    CascadeMux I__2661 (
            .O(N__24561),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ));
    InMux I__2660 (
            .O(N__24558),
            .I(N__24552));
    InMux I__2659 (
            .O(N__24557),
            .I(N__24552));
    LocalMux I__2658 (
            .O(N__24552),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ));
    InMux I__2657 (
            .O(N__24549),
            .I(N__24543));
    InMux I__2656 (
            .O(N__24548),
            .I(N__24543));
    LocalMux I__2655 (
            .O(N__24543),
            .I(N__24540));
    Span4Mux_h I__2654 (
            .O(N__24540),
            .I(N__24537));
    Span4Mux_v I__2653 (
            .O(N__24537),
            .I(N__24534));
    Span4Mux_v I__2652 (
            .O(N__24534),
            .I(N__24531));
    Odrv4 I__2651 (
            .O(N__24531),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    CascadeMux I__2650 (
            .O(N__24528),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_ ));
    InMux I__2649 (
            .O(N__24525),
            .I(N__24516));
    InMux I__2648 (
            .O(N__24524),
            .I(N__24516));
    InMux I__2647 (
            .O(N__24523),
            .I(N__24516));
    LocalMux I__2646 (
            .O(N__24516),
            .I(N__24513));
    Odrv12 I__2645 (
            .O(N__24513),
            .I(\pid_alt.error_d_regZ0Z_4 ));
    CascadeMux I__2644 (
            .O(N__24510),
            .I(N__24507));
    InMux I__2643 (
            .O(N__24507),
            .I(N__24501));
    InMux I__2642 (
            .O(N__24506),
            .I(N__24501));
    LocalMux I__2641 (
            .O(N__24501),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    InMux I__2640 (
            .O(N__24498),
            .I(N__24495));
    LocalMux I__2639 (
            .O(N__24495),
            .I(N__24492));
    Span4Mux_h I__2638 (
            .O(N__24492),
            .I(N__24489));
    Odrv4 I__2637 (
            .O(N__24489),
            .I(\pid_alt.O_4_4 ));
    InMux I__2636 (
            .O(N__24486),
            .I(N__24483));
    LocalMux I__2635 (
            .O(N__24483),
            .I(N__24480));
    Span4Mux_h I__2634 (
            .O(N__24480),
            .I(N__24477));
    Odrv4 I__2633 (
            .O(N__24477),
            .I(\pid_alt.O_4_7 ));
    InMux I__2632 (
            .O(N__24474),
            .I(N__24471));
    LocalMux I__2631 (
            .O(N__24471),
            .I(N__24468));
    Span4Mux_h I__2630 (
            .O(N__24468),
            .I(N__24465));
    Odrv4 I__2629 (
            .O(N__24465),
            .I(\pid_alt.O_4_15 ));
    CEMux I__2628 (
            .O(N__24462),
            .I(N__24417));
    CEMux I__2627 (
            .O(N__24461),
            .I(N__24417));
    CEMux I__2626 (
            .O(N__24460),
            .I(N__24417));
    CEMux I__2625 (
            .O(N__24459),
            .I(N__24417));
    CEMux I__2624 (
            .O(N__24458),
            .I(N__24417));
    CEMux I__2623 (
            .O(N__24457),
            .I(N__24417));
    CEMux I__2622 (
            .O(N__24456),
            .I(N__24417));
    CEMux I__2621 (
            .O(N__24455),
            .I(N__24417));
    CEMux I__2620 (
            .O(N__24454),
            .I(N__24417));
    CEMux I__2619 (
            .O(N__24453),
            .I(N__24417));
    CEMux I__2618 (
            .O(N__24452),
            .I(N__24417));
    CEMux I__2617 (
            .O(N__24451),
            .I(N__24417));
    CEMux I__2616 (
            .O(N__24450),
            .I(N__24417));
    CEMux I__2615 (
            .O(N__24449),
            .I(N__24417));
    CEMux I__2614 (
            .O(N__24448),
            .I(N__24417));
    GlobalMux I__2613 (
            .O(N__24417),
            .I(N__24414));
    gio2CtrlBuf I__2612 (
            .O(N__24414),
            .I(\pid_alt.N_664_0_g ));
    InMux I__2611 (
            .O(N__24411),
            .I(N__24408));
    LocalMux I__2610 (
            .O(N__24408),
            .I(N__24405));
    Span4Mux_s3_h I__2609 (
            .O(N__24405),
            .I(N__24402));
    Span4Mux_v I__2608 (
            .O(N__24402),
            .I(N__24399));
    Span4Mux_v I__2607 (
            .O(N__24399),
            .I(N__24396));
    Odrv4 I__2606 (
            .O(N__24396),
            .I(\Commands_frame_decoder.source_CH1data8lt7_0 ));
    InMux I__2605 (
            .O(N__24393),
            .I(N__24384));
    InMux I__2604 (
            .O(N__24392),
            .I(N__24384));
    InMux I__2603 (
            .O(N__24391),
            .I(N__24381));
    InMux I__2602 (
            .O(N__24390),
            .I(N__24378));
    InMux I__2601 (
            .O(N__24389),
            .I(N__24375));
    LocalMux I__2600 (
            .O(N__24384),
            .I(N__24372));
    LocalMux I__2599 (
            .O(N__24381),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    LocalMux I__2598 (
            .O(N__24378),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    LocalMux I__2597 (
            .O(N__24375),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    Odrv4 I__2596 (
            .O(N__24372),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    InMux I__2595 (
            .O(N__24363),
            .I(N__24360));
    LocalMux I__2594 (
            .O(N__24360),
            .I(N__24357));
    Span4Mux_v I__2593 (
            .O(N__24357),
            .I(N__24354));
    Odrv4 I__2592 (
            .O(N__24354),
            .I(\pid_alt.O_5_9 ));
    InMux I__2591 (
            .O(N__24351),
            .I(N__24345));
    InMux I__2590 (
            .O(N__24350),
            .I(N__24345));
    LocalMux I__2589 (
            .O(N__24345),
            .I(N__24342));
    Odrv12 I__2588 (
            .O(N__24342),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    InMux I__2587 (
            .O(N__24339),
            .I(N__24336));
    LocalMux I__2586 (
            .O(N__24336),
            .I(N__24333));
    Span4Mux_h I__2585 (
            .O(N__24333),
            .I(N__24330));
    Odrv4 I__2584 (
            .O(N__24330),
            .I(\pid_alt.O_5_10 ));
    InMux I__2583 (
            .O(N__24327),
            .I(N__24321));
    InMux I__2582 (
            .O(N__24326),
            .I(N__24321));
    LocalMux I__2581 (
            .O(N__24321),
            .I(N__24318));
    Span12Mux_v I__2580 (
            .O(N__24318),
            .I(N__24315));
    Odrv12 I__2579 (
            .O(N__24315),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    InMux I__2578 (
            .O(N__24312),
            .I(N__24309));
    LocalMux I__2577 (
            .O(N__24309),
            .I(N__24306));
    Odrv4 I__2576 (
            .O(N__24306),
            .I(alt_kp_7));
    InMux I__2575 (
            .O(N__24303),
            .I(N__24300));
    LocalMux I__2574 (
            .O(N__24300),
            .I(N__24297));
    Odrv4 I__2573 (
            .O(N__24297),
            .I(alt_kp_3));
    InMux I__2572 (
            .O(N__24294),
            .I(N__24291));
    LocalMux I__2571 (
            .O(N__24291),
            .I(N__24288));
    Span4Mux_v I__2570 (
            .O(N__24288),
            .I(N__24285));
    Odrv4 I__2569 (
            .O(N__24285),
            .I(\pid_alt.O_3_8 ));
    CEMux I__2568 (
            .O(N__24282),
            .I(N__24279));
    LocalMux I__2567 (
            .O(N__24279),
            .I(N__24276));
    Span4Mux_h I__2566 (
            .O(N__24276),
            .I(N__24272));
    CEMux I__2565 (
            .O(N__24275),
            .I(N__24268));
    Span4Mux_s0_h I__2564 (
            .O(N__24272),
            .I(N__24265));
    CEMux I__2563 (
            .O(N__24271),
            .I(N__24262));
    LocalMux I__2562 (
            .O(N__24268),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    Odrv4 I__2561 (
            .O(N__24265),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    LocalMux I__2560 (
            .O(N__24262),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    InMux I__2559 (
            .O(N__24255),
            .I(N__24252));
    LocalMux I__2558 (
            .O(N__24252),
            .I(N__24249));
    Span4Mux_h I__2557 (
            .O(N__24249),
            .I(N__24246));
    Odrv4 I__2556 (
            .O(N__24246),
            .I(\pid_alt.O_3_11 ));
    InMux I__2555 (
            .O(N__24243),
            .I(N__24240));
    LocalMux I__2554 (
            .O(N__24240),
            .I(N__24237));
    Span4Mux_h I__2553 (
            .O(N__24237),
            .I(N__24234));
    Odrv4 I__2552 (
            .O(N__24234),
            .I(\pid_alt.O_3_12 ));
    InMux I__2551 (
            .O(N__24231),
            .I(N__24228));
    LocalMux I__2550 (
            .O(N__24228),
            .I(N__24225));
    Span4Mux_h I__2549 (
            .O(N__24225),
            .I(N__24222));
    Odrv4 I__2548 (
            .O(N__24222),
            .I(\pid_alt.O_3_13 ));
    CascadeMux I__2547 (
            .O(N__24219),
            .I(N__24216));
    InMux I__2546 (
            .O(N__24216),
            .I(N__24213));
    LocalMux I__2545 (
            .O(N__24213),
            .I(N__24210));
    Odrv4 I__2544 (
            .O(N__24210),
            .I(alt_command_7));
    InMux I__2543 (
            .O(N__24207),
            .I(N__24202));
    InMux I__2542 (
            .O(N__24206),
            .I(N__24199));
    InMux I__2541 (
            .O(N__24205),
            .I(N__24196));
    LocalMux I__2540 (
            .O(N__24202),
            .I(N__24193));
    LocalMux I__2539 (
            .O(N__24199),
            .I(N__24190));
    LocalMux I__2538 (
            .O(N__24196),
            .I(N__24187));
    Span12Mux_s2_h I__2537 (
            .O(N__24193),
            .I(N__24184));
    Span4Mux_s2_h I__2536 (
            .O(N__24190),
            .I(N__24181));
    Span4Mux_s2_h I__2535 (
            .O(N__24187),
            .I(N__24178));
    Span12Mux_v I__2534 (
            .O(N__24184),
            .I(N__24175));
    Span4Mux_v I__2533 (
            .O(N__24181),
            .I(N__24172));
    Span4Mux_v I__2532 (
            .O(N__24178),
            .I(N__24169));
    Odrv12 I__2531 (
            .O(N__24175),
            .I(\pid_alt.error_11 ));
    Odrv4 I__2530 (
            .O(N__24172),
            .I(\pid_alt.error_11 ));
    Odrv4 I__2529 (
            .O(N__24169),
            .I(\pid_alt.error_11 ));
    InMux I__2528 (
            .O(N__24162),
            .I(\pid_alt.error_cry_10 ));
    InMux I__2527 (
            .O(N__24159),
            .I(N__24156));
    LocalMux I__2526 (
            .O(N__24156),
            .I(N__24153));
    Span4Mux_v I__2525 (
            .O(N__24153),
            .I(N__24148));
    InMux I__2524 (
            .O(N__24152),
            .I(N__24145));
    InMux I__2523 (
            .O(N__24151),
            .I(N__24142));
    Span4Mux_v I__2522 (
            .O(N__24148),
            .I(N__24139));
    LocalMux I__2521 (
            .O(N__24145),
            .I(N__24136));
    LocalMux I__2520 (
            .O(N__24142),
            .I(N__24133));
    Span4Mux_v I__2519 (
            .O(N__24139),
            .I(N__24130));
    Span4Mux_v I__2518 (
            .O(N__24136),
            .I(N__24127));
    Span12Mux_s2_h I__2517 (
            .O(N__24133),
            .I(N__24124));
    Span4Mux_v I__2516 (
            .O(N__24130),
            .I(N__24119));
    Span4Mux_v I__2515 (
            .O(N__24127),
            .I(N__24119));
    Odrv12 I__2514 (
            .O(N__24124),
            .I(\pid_alt.error_12 ));
    Odrv4 I__2513 (
            .O(N__24119),
            .I(\pid_alt.error_12 ));
    InMux I__2512 (
            .O(N__24114),
            .I(\pid_alt.error_cry_11 ));
    InMux I__2511 (
            .O(N__24111),
            .I(N__24108));
    LocalMux I__2510 (
            .O(N__24108),
            .I(N__24104));
    InMux I__2509 (
            .O(N__24107),
            .I(N__24101));
    Span4Mux_s1_h I__2508 (
            .O(N__24104),
            .I(N__24097));
    LocalMux I__2507 (
            .O(N__24101),
            .I(N__24094));
    InMux I__2506 (
            .O(N__24100),
            .I(N__24091));
    Sp12to4 I__2505 (
            .O(N__24097),
            .I(N__24088));
    Span4Mux_s2_h I__2504 (
            .O(N__24094),
            .I(N__24085));
    LocalMux I__2503 (
            .O(N__24091),
            .I(N__24082));
    Span12Mux_v I__2502 (
            .O(N__24088),
            .I(N__24079));
    Span4Mux_v I__2501 (
            .O(N__24085),
            .I(N__24076));
    Span12Mux_s2_h I__2500 (
            .O(N__24082),
            .I(N__24073));
    Odrv12 I__2499 (
            .O(N__24079),
            .I(\pid_alt.error_13 ));
    Odrv4 I__2498 (
            .O(N__24076),
            .I(\pid_alt.error_13 ));
    Odrv12 I__2497 (
            .O(N__24073),
            .I(\pid_alt.error_13 ));
    InMux I__2496 (
            .O(N__24066),
            .I(\pid_alt.error_cry_12 ));
    InMux I__2495 (
            .O(N__24063),
            .I(N__24059));
    InMux I__2494 (
            .O(N__24062),
            .I(N__24055));
    LocalMux I__2493 (
            .O(N__24059),
            .I(N__24052));
    InMux I__2492 (
            .O(N__24058),
            .I(N__24049));
    LocalMux I__2491 (
            .O(N__24055),
            .I(N__24046));
    Span12Mux_s7_v I__2490 (
            .O(N__24052),
            .I(N__24041));
    LocalMux I__2489 (
            .O(N__24049),
            .I(N__24041));
    Span4Mux_s2_h I__2488 (
            .O(N__24046),
            .I(N__24038));
    Span12Mux_v I__2487 (
            .O(N__24041),
            .I(N__24035));
    Span4Mux_v I__2486 (
            .O(N__24038),
            .I(N__24032));
    Odrv12 I__2485 (
            .O(N__24035),
            .I(\pid_alt.error_14 ));
    Odrv4 I__2484 (
            .O(N__24032),
            .I(\pid_alt.error_14 ));
    InMux I__2483 (
            .O(N__24027),
            .I(\pid_alt.error_cry_13 ));
    InMux I__2482 (
            .O(N__24024),
            .I(\pid_alt.error_cry_14 ));
    InMux I__2481 (
            .O(N__24021),
            .I(N__24018));
    LocalMux I__2480 (
            .O(N__24018),
            .I(N__24014));
    InMux I__2479 (
            .O(N__24017),
            .I(N__24011));
    Span4Mux_v I__2478 (
            .O(N__24014),
            .I(N__24007));
    LocalMux I__2477 (
            .O(N__24011),
            .I(N__24004));
    InMux I__2476 (
            .O(N__24010),
            .I(N__24001));
    Span4Mux_v I__2475 (
            .O(N__24007),
            .I(N__23996));
    Span4Mux_s1_h I__2474 (
            .O(N__24004),
            .I(N__23996));
    LocalMux I__2473 (
            .O(N__24001),
            .I(N__23993));
    Span4Mux_v I__2472 (
            .O(N__23996),
            .I(N__23990));
    Span4Mux_s2_h I__2471 (
            .O(N__23993),
            .I(N__23987));
    Span4Mux_v I__2470 (
            .O(N__23990),
            .I(N__23984));
    Span4Mux_v I__2469 (
            .O(N__23987),
            .I(N__23981));
    Odrv4 I__2468 (
            .O(N__23984),
            .I(\pid_alt.error_15 ));
    Odrv4 I__2467 (
            .O(N__23981),
            .I(\pid_alt.error_15 ));
    InMux I__2466 (
            .O(N__23976),
            .I(N__23973));
    LocalMux I__2465 (
            .O(N__23973),
            .I(N__23970));
    Span4Mux_v I__2464 (
            .O(N__23970),
            .I(N__23967));
    Odrv4 I__2463 (
            .O(N__23967),
            .I(alt_kp_1));
    InMux I__2462 (
            .O(N__23964),
            .I(N__23961));
    LocalMux I__2461 (
            .O(N__23961),
            .I(drone_altitude_i_10));
    InMux I__2460 (
            .O(N__23958),
            .I(N__23955));
    LocalMux I__2459 (
            .O(N__23955),
            .I(N__23952));
    Span4Mux_s2_h I__2458 (
            .O(N__23952),
            .I(N__23949));
    Odrv4 I__2457 (
            .O(N__23949),
            .I(alt_kp_0));
    InMux I__2456 (
            .O(N__23946),
            .I(N__23943));
    LocalMux I__2455 (
            .O(N__23943),
            .I(N__23940));
    Span4Mux_s2_h I__2454 (
            .O(N__23940),
            .I(N__23937));
    Odrv4 I__2453 (
            .O(N__23937),
            .I(alt_kp_6));
    InMux I__2452 (
            .O(N__23934),
            .I(N__23930));
    CascadeMux I__2451 (
            .O(N__23933),
            .I(N__23927));
    LocalMux I__2450 (
            .O(N__23930),
            .I(N__23924));
    InMux I__2449 (
            .O(N__23927),
            .I(N__23921));
    Odrv12 I__2448 (
            .O(N__23924),
            .I(alt_command_0));
    LocalMux I__2447 (
            .O(N__23921),
            .I(alt_command_0));
    InMux I__2446 (
            .O(N__23916),
            .I(N__23913));
    LocalMux I__2445 (
            .O(N__23913),
            .I(N__23910));
    Span4Mux_h I__2444 (
            .O(N__23910),
            .I(N__23905));
    InMux I__2443 (
            .O(N__23909),
            .I(N__23902));
    InMux I__2442 (
            .O(N__23908),
            .I(N__23899));
    Span4Mux_v I__2441 (
            .O(N__23905),
            .I(N__23894));
    LocalMux I__2440 (
            .O(N__23902),
            .I(N__23894));
    LocalMux I__2439 (
            .O(N__23899),
            .I(N__23891));
    Span4Mux_v I__2438 (
            .O(N__23894),
            .I(N__23888));
    Span4Mux_s3_h I__2437 (
            .O(N__23891),
            .I(N__23885));
    Span4Mux_v I__2436 (
            .O(N__23888),
            .I(N__23882));
    Span4Mux_v I__2435 (
            .O(N__23885),
            .I(N__23879));
    Odrv4 I__2434 (
            .O(N__23882),
            .I(\pid_alt.error_4 ));
    Odrv4 I__2433 (
            .O(N__23879),
            .I(\pid_alt.error_4 ));
    InMux I__2432 (
            .O(N__23874),
            .I(\pid_alt.error_cry_3 ));
    CascadeMux I__2431 (
            .O(N__23871),
            .I(N__23867));
    InMux I__2430 (
            .O(N__23870),
            .I(N__23864));
    InMux I__2429 (
            .O(N__23867),
            .I(N__23861));
    LocalMux I__2428 (
            .O(N__23864),
            .I(alt_command_1));
    LocalMux I__2427 (
            .O(N__23861),
            .I(alt_command_1));
    InMux I__2426 (
            .O(N__23856),
            .I(N__23853));
    LocalMux I__2425 (
            .O(N__23853),
            .I(N__23850));
    Span4Mux_h I__2424 (
            .O(N__23850),
            .I(N__23845));
    InMux I__2423 (
            .O(N__23849),
            .I(N__23842));
    InMux I__2422 (
            .O(N__23848),
            .I(N__23839));
    Span4Mux_v I__2421 (
            .O(N__23845),
            .I(N__23834));
    LocalMux I__2420 (
            .O(N__23842),
            .I(N__23834));
    LocalMux I__2419 (
            .O(N__23839),
            .I(N__23831));
    Span4Mux_v I__2418 (
            .O(N__23834),
            .I(N__23828));
    Span4Mux_s2_h I__2417 (
            .O(N__23831),
            .I(N__23825));
    Span4Mux_v I__2416 (
            .O(N__23828),
            .I(N__23822));
    Span4Mux_v I__2415 (
            .O(N__23825),
            .I(N__23819));
    Odrv4 I__2414 (
            .O(N__23822),
            .I(\pid_alt.error_5 ));
    Odrv4 I__2413 (
            .O(N__23819),
            .I(\pid_alt.error_5 ));
    InMux I__2412 (
            .O(N__23814),
            .I(\pid_alt.error_cry_4 ));
    CascadeMux I__2411 (
            .O(N__23811),
            .I(N__23807));
    InMux I__2410 (
            .O(N__23810),
            .I(N__23804));
    InMux I__2409 (
            .O(N__23807),
            .I(N__23801));
    LocalMux I__2408 (
            .O(N__23804),
            .I(alt_command_2));
    LocalMux I__2407 (
            .O(N__23801),
            .I(alt_command_2));
    InMux I__2406 (
            .O(N__23796),
            .I(N__23791));
    InMux I__2405 (
            .O(N__23795),
            .I(N__23788));
    InMux I__2404 (
            .O(N__23794),
            .I(N__23785));
    LocalMux I__2403 (
            .O(N__23791),
            .I(N__23782));
    LocalMux I__2402 (
            .O(N__23788),
            .I(N__23779));
    LocalMux I__2401 (
            .O(N__23785),
            .I(N__23776));
    Span12Mux_s4_h I__2400 (
            .O(N__23782),
            .I(N__23773));
    Span4Mux_s2_h I__2399 (
            .O(N__23779),
            .I(N__23770));
    Span4Mux_s2_h I__2398 (
            .O(N__23776),
            .I(N__23767));
    Span12Mux_v I__2397 (
            .O(N__23773),
            .I(N__23764));
    Span4Mux_v I__2396 (
            .O(N__23770),
            .I(N__23761));
    Span4Mux_v I__2395 (
            .O(N__23767),
            .I(N__23758));
    Odrv12 I__2394 (
            .O(N__23764),
            .I(\pid_alt.error_6 ));
    Odrv4 I__2393 (
            .O(N__23761),
            .I(\pid_alt.error_6 ));
    Odrv4 I__2392 (
            .O(N__23758),
            .I(\pid_alt.error_6 ));
    InMux I__2391 (
            .O(N__23751),
            .I(\pid_alt.error_cry_5 ));
    CascadeMux I__2390 (
            .O(N__23748),
            .I(N__23744));
    InMux I__2389 (
            .O(N__23747),
            .I(N__23741));
    InMux I__2388 (
            .O(N__23744),
            .I(N__23738));
    LocalMux I__2387 (
            .O(N__23741),
            .I(alt_command_3));
    LocalMux I__2386 (
            .O(N__23738),
            .I(alt_command_3));
    InMux I__2385 (
            .O(N__23733),
            .I(N__23728));
    InMux I__2384 (
            .O(N__23732),
            .I(N__23725));
    InMux I__2383 (
            .O(N__23731),
            .I(N__23722));
    LocalMux I__2382 (
            .O(N__23728),
            .I(N__23719));
    LocalMux I__2381 (
            .O(N__23725),
            .I(N__23716));
    LocalMux I__2380 (
            .O(N__23722),
            .I(N__23713));
    Span12Mux_s3_h I__2379 (
            .O(N__23719),
            .I(N__23710));
    Span4Mux_s2_h I__2378 (
            .O(N__23716),
            .I(N__23707));
    Span4Mux_s2_h I__2377 (
            .O(N__23713),
            .I(N__23704));
    Span12Mux_v I__2376 (
            .O(N__23710),
            .I(N__23701));
    Span4Mux_v I__2375 (
            .O(N__23707),
            .I(N__23698));
    Span4Mux_v I__2374 (
            .O(N__23704),
            .I(N__23695));
    Odrv12 I__2373 (
            .O(N__23701),
            .I(\pid_alt.error_7 ));
    Odrv4 I__2372 (
            .O(N__23698),
            .I(\pid_alt.error_7 ));
    Odrv4 I__2371 (
            .O(N__23695),
            .I(\pid_alt.error_7 ));
    InMux I__2370 (
            .O(N__23688),
            .I(\pid_alt.error_cry_6 ));
    CascadeMux I__2369 (
            .O(N__23685),
            .I(N__23682));
    InMux I__2368 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__2367 (
            .O(N__23679),
            .I(alt_command_4));
    InMux I__2366 (
            .O(N__23676),
            .I(N__23673));
    LocalMux I__2365 (
            .O(N__23673),
            .I(N__23670));
    Span4Mux_v I__2364 (
            .O(N__23670),
            .I(N__23665));
    InMux I__2363 (
            .O(N__23669),
            .I(N__23662));
    InMux I__2362 (
            .O(N__23668),
            .I(N__23659));
    Span4Mux_v I__2361 (
            .O(N__23665),
            .I(N__23656));
    LocalMux I__2360 (
            .O(N__23662),
            .I(N__23653));
    LocalMux I__2359 (
            .O(N__23659),
            .I(N__23650));
    Span4Mux_v I__2358 (
            .O(N__23656),
            .I(N__23647));
    Span4Mux_s2_h I__2357 (
            .O(N__23653),
            .I(N__23644));
    Span4Mux_s3_h I__2356 (
            .O(N__23650),
            .I(N__23641));
    Span4Mux_v I__2355 (
            .O(N__23647),
            .I(N__23638));
    Span4Mux_v I__2354 (
            .O(N__23644),
            .I(N__23635));
    Span4Mux_v I__2353 (
            .O(N__23641),
            .I(N__23632));
    Odrv4 I__2352 (
            .O(N__23638),
            .I(\pid_alt.error_8 ));
    Odrv4 I__2351 (
            .O(N__23635),
            .I(\pid_alt.error_8 ));
    Odrv4 I__2350 (
            .O(N__23632),
            .I(\pid_alt.error_8 ));
    InMux I__2349 (
            .O(N__23625),
            .I(bfn_2_20_0_));
    CascadeMux I__2348 (
            .O(N__23622),
            .I(N__23619));
    InMux I__2347 (
            .O(N__23619),
            .I(N__23616));
    LocalMux I__2346 (
            .O(N__23616),
            .I(N__23613));
    Odrv4 I__2345 (
            .O(N__23613),
            .I(alt_command_5));
    InMux I__2344 (
            .O(N__23610),
            .I(N__23607));
    LocalMux I__2343 (
            .O(N__23607),
            .I(N__23602));
    InMux I__2342 (
            .O(N__23606),
            .I(N__23599));
    InMux I__2341 (
            .O(N__23605),
            .I(N__23596));
    Span4Mux_v I__2340 (
            .O(N__23602),
            .I(N__23593));
    LocalMux I__2339 (
            .O(N__23599),
            .I(N__23590));
    LocalMux I__2338 (
            .O(N__23596),
            .I(N__23587));
    Sp12to4 I__2337 (
            .O(N__23593),
            .I(N__23584));
    Span4Mux_s2_h I__2336 (
            .O(N__23590),
            .I(N__23581));
    Span4Mux_s2_h I__2335 (
            .O(N__23587),
            .I(N__23578));
    Span12Mux_s2_h I__2334 (
            .O(N__23584),
            .I(N__23575));
    Span4Mux_v I__2333 (
            .O(N__23581),
            .I(N__23572));
    Span4Mux_v I__2332 (
            .O(N__23578),
            .I(N__23569));
    Odrv12 I__2331 (
            .O(N__23575),
            .I(\pid_alt.error_9 ));
    Odrv4 I__2330 (
            .O(N__23572),
            .I(\pid_alt.error_9 ));
    Odrv4 I__2329 (
            .O(N__23569),
            .I(\pid_alt.error_9 ));
    InMux I__2328 (
            .O(N__23562),
            .I(\pid_alt.error_cry_8 ));
    CascadeMux I__2327 (
            .O(N__23559),
            .I(N__23556));
    InMux I__2326 (
            .O(N__23556),
            .I(N__23553));
    LocalMux I__2325 (
            .O(N__23553),
            .I(alt_command_6));
    InMux I__2324 (
            .O(N__23550),
            .I(N__23547));
    LocalMux I__2323 (
            .O(N__23547),
            .I(N__23544));
    Span4Mux_s2_h I__2322 (
            .O(N__23544),
            .I(N__23539));
    InMux I__2321 (
            .O(N__23543),
            .I(N__23536));
    InMux I__2320 (
            .O(N__23542),
            .I(N__23533));
    Span4Mux_v I__2319 (
            .O(N__23539),
            .I(N__23530));
    LocalMux I__2318 (
            .O(N__23536),
            .I(N__23527));
    LocalMux I__2317 (
            .O(N__23533),
            .I(N__23524));
    Span4Mux_v I__2316 (
            .O(N__23530),
            .I(N__23521));
    Span4Mux_s2_h I__2315 (
            .O(N__23527),
            .I(N__23518));
    Span4Mux_s3_h I__2314 (
            .O(N__23524),
            .I(N__23515));
    Span4Mux_v I__2313 (
            .O(N__23521),
            .I(N__23512));
    Span4Mux_v I__2312 (
            .O(N__23518),
            .I(N__23509));
    Span4Mux_v I__2311 (
            .O(N__23515),
            .I(N__23506));
    Odrv4 I__2310 (
            .O(N__23512),
            .I(\pid_alt.error_10 ));
    Odrv4 I__2309 (
            .O(N__23509),
            .I(\pid_alt.error_10 ));
    Odrv4 I__2308 (
            .O(N__23506),
            .I(\pid_alt.error_10 ));
    InMux I__2307 (
            .O(N__23499),
            .I(\pid_alt.error_cry_9 ));
    CascadeMux I__2306 (
            .O(N__23496),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ));
    InMux I__2305 (
            .O(N__23493),
            .I(N__23487));
    InMux I__2304 (
            .O(N__23492),
            .I(N__23487));
    LocalMux I__2303 (
            .O(N__23487),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ));
    InMux I__2302 (
            .O(N__23484),
            .I(N__23478));
    InMux I__2301 (
            .O(N__23483),
            .I(N__23478));
    LocalMux I__2300 (
            .O(N__23478),
            .I(N__23475));
    Span4Mux_h I__2299 (
            .O(N__23475),
            .I(N__23472));
    Odrv4 I__2298 (
            .O(N__23472),
            .I(\pid_alt.error_p_regZ0Z_18 ));
    InMux I__2297 (
            .O(N__23469),
            .I(N__23463));
    InMux I__2296 (
            .O(N__23468),
            .I(N__23463));
    LocalMux I__2295 (
            .O(N__23463),
            .I(\pid_alt.error_d_reg_prevZ0Z_18 ));
    InMux I__2294 (
            .O(N__23460),
            .I(N__23451));
    InMux I__2293 (
            .O(N__23459),
            .I(N__23451));
    InMux I__2292 (
            .O(N__23458),
            .I(N__23451));
    LocalMux I__2291 (
            .O(N__23451),
            .I(N__23448));
    Span12Mux_s8_h I__2290 (
            .O(N__23448),
            .I(N__23445));
    Span12Mux_v I__2289 (
            .O(N__23445),
            .I(N__23442));
    Odrv12 I__2288 (
            .O(N__23442),
            .I(\pid_alt.error_d_regZ0Z_18 ));
    CascadeMux I__2287 (
            .O(N__23439),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ));
    InMux I__2286 (
            .O(N__23436),
            .I(N__23433));
    LocalMux I__2285 (
            .O(N__23433),
            .I(N__23430));
    Span4Mux_s1_h I__2284 (
            .O(N__23430),
            .I(N__23426));
    InMux I__2283 (
            .O(N__23429),
            .I(N__23423));
    Span4Mux_v I__2282 (
            .O(N__23426),
            .I(N__23417));
    LocalMux I__2281 (
            .O(N__23423),
            .I(N__23417));
    InMux I__2280 (
            .O(N__23422),
            .I(N__23414));
    Span4Mux_v I__2279 (
            .O(N__23417),
            .I(N__23411));
    LocalMux I__2278 (
            .O(N__23414),
            .I(N__23408));
    Span4Mux_v I__2277 (
            .O(N__23411),
            .I(N__23403));
    Span4Mux_v I__2276 (
            .O(N__23408),
            .I(N__23403));
    Span4Mux_v I__2275 (
            .O(N__23403),
            .I(N__23400));
    Odrv4 I__2274 (
            .O(N__23400),
            .I(\pid_alt.error_1 ));
    InMux I__2273 (
            .O(N__23397),
            .I(\pid_alt.error_cry_0 ));
    InMux I__2272 (
            .O(N__23394),
            .I(N__23391));
    LocalMux I__2271 (
            .O(N__23391),
            .I(N__23388));
    Span4Mux_s1_h I__2270 (
            .O(N__23388),
            .I(N__23383));
    InMux I__2269 (
            .O(N__23387),
            .I(N__23380));
    InMux I__2268 (
            .O(N__23386),
            .I(N__23377));
    Span4Mux_v I__2267 (
            .O(N__23383),
            .I(N__23372));
    LocalMux I__2266 (
            .O(N__23380),
            .I(N__23372));
    LocalMux I__2265 (
            .O(N__23377),
            .I(N__23369));
    Span4Mux_v I__2264 (
            .O(N__23372),
            .I(N__23366));
    Span4Mux_v I__2263 (
            .O(N__23369),
            .I(N__23363));
    Span4Mux_v I__2262 (
            .O(N__23366),
            .I(N__23358));
    Span4Mux_v I__2261 (
            .O(N__23363),
            .I(N__23358));
    Odrv4 I__2260 (
            .O(N__23358),
            .I(\pid_alt.error_2 ));
    InMux I__2259 (
            .O(N__23355),
            .I(\pid_alt.error_cry_1 ));
    InMux I__2258 (
            .O(N__23352),
            .I(N__23349));
    LocalMux I__2257 (
            .O(N__23349),
            .I(N__23346));
    Span4Mux_s1_h I__2256 (
            .O(N__23346),
            .I(N__23342));
    InMux I__2255 (
            .O(N__23345),
            .I(N__23339));
    Span4Mux_v I__2254 (
            .O(N__23342),
            .I(N__23333));
    LocalMux I__2253 (
            .O(N__23339),
            .I(N__23333));
    InMux I__2252 (
            .O(N__23338),
            .I(N__23330));
    Span4Mux_v I__2251 (
            .O(N__23333),
            .I(N__23327));
    LocalMux I__2250 (
            .O(N__23330),
            .I(N__23324));
    Span4Mux_v I__2249 (
            .O(N__23327),
            .I(N__23321));
    Span4Mux_v I__2248 (
            .O(N__23324),
            .I(N__23318));
    Span4Mux_s1_h I__2247 (
            .O(N__23321),
            .I(N__23313));
    Span4Mux_v I__2246 (
            .O(N__23318),
            .I(N__23313));
    Odrv4 I__2245 (
            .O(N__23313),
            .I(\pid_alt.error_3 ));
    InMux I__2244 (
            .O(N__23310),
            .I(\pid_alt.error_cry_2 ));
    InMux I__2243 (
            .O(N__23307),
            .I(N__23304));
    LocalMux I__2242 (
            .O(N__23304),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ));
    CascadeMux I__2241 (
            .O(N__23301),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ));
    InMux I__2240 (
            .O(N__23298),
            .I(N__23292));
    InMux I__2239 (
            .O(N__23297),
            .I(N__23292));
    LocalMux I__2238 (
            .O(N__23292),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ));
    InMux I__2237 (
            .O(N__23289),
            .I(N__23280));
    InMux I__2236 (
            .O(N__23288),
            .I(N__23280));
    InMux I__2235 (
            .O(N__23287),
            .I(N__23280));
    LocalMux I__2234 (
            .O(N__23280),
            .I(N__23277));
    Span4Mux_h I__2233 (
            .O(N__23277),
            .I(N__23274));
    Sp12to4 I__2232 (
            .O(N__23274),
            .I(N__23271));
    Odrv12 I__2231 (
            .O(N__23271),
            .I(\pid_alt.error_d_regZ0Z_12 ));
    CascadeMux I__2230 (
            .O(N__23268),
            .I(N__23265));
    InMux I__2229 (
            .O(N__23265),
            .I(N__23259));
    InMux I__2228 (
            .O(N__23264),
            .I(N__23259));
    LocalMux I__2227 (
            .O(N__23259),
            .I(\pid_alt.error_d_reg_prevZ0Z_12 ));
    InMux I__2226 (
            .O(N__23256),
            .I(N__23250));
    InMux I__2225 (
            .O(N__23255),
            .I(N__23250));
    LocalMux I__2224 (
            .O(N__23250),
            .I(N__23247));
    Span4Mux_v I__2223 (
            .O(N__23247),
            .I(N__23244));
    Span4Mux_v I__2222 (
            .O(N__23244),
            .I(N__23241));
    Odrv4 I__2221 (
            .O(N__23241),
            .I(\pid_alt.error_p_regZ0Z_12 ));
    CascadeMux I__2220 (
            .O(N__23238),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ));
    InMux I__2219 (
            .O(N__23235),
            .I(N__23232));
    LocalMux I__2218 (
            .O(N__23232),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ));
    InMux I__2217 (
            .O(N__23229),
            .I(N__23225));
    InMux I__2216 (
            .O(N__23228),
            .I(N__23220));
    LocalMux I__2215 (
            .O(N__23225),
            .I(N__23217));
    InMux I__2214 (
            .O(N__23224),
            .I(N__23212));
    InMux I__2213 (
            .O(N__23223),
            .I(N__23212));
    LocalMux I__2212 (
            .O(N__23220),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    Odrv4 I__2211 (
            .O(N__23217),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    LocalMux I__2210 (
            .O(N__23212),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    CascadeMux I__2209 (
            .O(N__23205),
            .I(N__23202));
    InMux I__2208 (
            .O(N__23202),
            .I(N__23199));
    LocalMux I__2207 (
            .O(N__23199),
            .I(\pid_alt.N_1666_i ));
    InMux I__2206 (
            .O(N__23196),
            .I(N__23186));
    InMux I__2205 (
            .O(N__23195),
            .I(N__23186));
    InMux I__2204 (
            .O(N__23194),
            .I(N__23181));
    InMux I__2203 (
            .O(N__23193),
            .I(N__23181));
    InMux I__2202 (
            .O(N__23192),
            .I(N__23176));
    InMux I__2201 (
            .O(N__23191),
            .I(N__23176));
    LocalMux I__2200 (
            .O(N__23186),
            .I(N__23173));
    LocalMux I__2199 (
            .O(N__23181),
            .I(N__23166));
    LocalMux I__2198 (
            .O(N__23176),
            .I(N__23166));
    Span4Mux_s2_h I__2197 (
            .O(N__23173),
            .I(N__23166));
    Odrv4 I__2196 (
            .O(N__23166),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    CascadeMux I__2195 (
            .O(N__23163),
            .I(N__23157));
    CascadeMux I__2194 (
            .O(N__23162),
            .I(N__23153));
    InMux I__2193 (
            .O(N__23161),
            .I(N__23147));
    InMux I__2192 (
            .O(N__23160),
            .I(N__23147));
    InMux I__2191 (
            .O(N__23157),
            .I(N__23142));
    InMux I__2190 (
            .O(N__23156),
            .I(N__23142));
    InMux I__2189 (
            .O(N__23153),
            .I(N__23137));
    InMux I__2188 (
            .O(N__23152),
            .I(N__23137));
    LocalMux I__2187 (
            .O(N__23147),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    LocalMux I__2186 (
            .O(N__23142),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    LocalMux I__2185 (
            .O(N__23137),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__2184 (
            .O(N__23130),
            .I(\pid_alt.N_1666_i_cascade_ ));
    InMux I__2183 (
            .O(N__23127),
            .I(N__23121));
    InMux I__2182 (
            .O(N__23126),
            .I(N__23121));
    LocalMux I__2181 (
            .O(N__23121),
            .I(N__23115));
    InMux I__2180 (
            .O(N__23120),
            .I(N__23108));
    InMux I__2179 (
            .O(N__23119),
            .I(N__23108));
    InMux I__2178 (
            .O(N__23118),
            .I(N__23108));
    Span4Mux_v I__2177 (
            .O(N__23115),
            .I(N__23103));
    LocalMux I__2176 (
            .O(N__23108),
            .I(N__23100));
    InMux I__2175 (
            .O(N__23107),
            .I(N__23095));
    InMux I__2174 (
            .O(N__23106),
            .I(N__23095));
    Span4Mux_v I__2173 (
            .O(N__23103),
            .I(N__23092));
    Span12Mux_v I__2172 (
            .O(N__23100),
            .I(N__23087));
    LocalMux I__2171 (
            .O(N__23095),
            .I(N__23087));
    Odrv4 I__2170 (
            .O(N__23092),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    Odrv12 I__2169 (
            .O(N__23087),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    InMux I__2168 (
            .O(N__23082),
            .I(N__23079));
    LocalMux I__2167 (
            .O(N__23079),
            .I(\pid_alt.un1_pid_prereg_0_axb_2_1 ));
    InMux I__2166 (
            .O(N__23076),
            .I(N__23073));
    LocalMux I__2165 (
            .O(N__23073),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ));
    CascadeMux I__2164 (
            .O(N__23070),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ));
    InMux I__2163 (
            .O(N__23067),
            .I(N__23064));
    LocalMux I__2162 (
            .O(N__23064),
            .I(N__23060));
    InMux I__2161 (
            .O(N__23063),
            .I(N__23057));
    Span4Mux_v I__2160 (
            .O(N__23060),
            .I(N__23054));
    LocalMux I__2159 (
            .O(N__23057),
            .I(N__23051));
    Span4Mux_v I__2158 (
            .O(N__23054),
            .I(N__23046));
    Span4Mux_v I__2157 (
            .O(N__23051),
            .I(N__23046));
    Odrv4 I__2156 (
            .O(N__23046),
            .I(\pid_alt.error_p_regZ0Z_11 ));
    InMux I__2155 (
            .O(N__23043),
            .I(N__23037));
    InMux I__2154 (
            .O(N__23042),
            .I(N__23037));
    LocalMux I__2153 (
            .O(N__23037),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ));
    InMux I__2152 (
            .O(N__23034),
            .I(N__23027));
    InMux I__2151 (
            .O(N__23033),
            .I(N__23027));
    InMux I__2150 (
            .O(N__23032),
            .I(N__23024));
    LocalMux I__2149 (
            .O(N__23027),
            .I(N__23021));
    LocalMux I__2148 (
            .O(N__23024),
            .I(N__23016));
    Span4Mux_v I__2147 (
            .O(N__23021),
            .I(N__23016));
    Span4Mux_v I__2146 (
            .O(N__23016),
            .I(N__23013));
    Odrv4 I__2145 (
            .O(N__23013),
            .I(\pid_alt.error_d_regZ0Z_11 ));
    InMux I__2144 (
            .O(N__23010),
            .I(N__23007));
    LocalMux I__2143 (
            .O(N__23007),
            .I(N__23004));
    Span4Mux_s3_h I__2142 (
            .O(N__23004),
            .I(N__23000));
    InMux I__2141 (
            .O(N__23003),
            .I(N__22997));
    Odrv4 I__2140 (
            .O(N__23000),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    LocalMux I__2139 (
            .O(N__22997),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    InMux I__2138 (
            .O(N__22992),
            .I(N__22986));
    InMux I__2137 (
            .O(N__22991),
            .I(N__22986));
    LocalMux I__2136 (
            .O(N__22986),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ));
    InMux I__2135 (
            .O(N__22983),
            .I(N__22977));
    InMux I__2134 (
            .O(N__22982),
            .I(N__22977));
    LocalMux I__2133 (
            .O(N__22977),
            .I(\pid_alt.error_d_reg_prevZ0Z_5 ));
    InMux I__2132 (
            .O(N__22974),
            .I(N__22965));
    InMux I__2131 (
            .O(N__22973),
            .I(N__22965));
    InMux I__2130 (
            .O(N__22972),
            .I(N__22965));
    LocalMux I__2129 (
            .O(N__22965),
            .I(N__22962));
    Span12Mux_v I__2128 (
            .O(N__22962),
            .I(N__22959));
    Odrv12 I__2127 (
            .O(N__22959),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    InMux I__2126 (
            .O(N__22956),
            .I(N__22950));
    InMux I__2125 (
            .O(N__22955),
            .I(N__22950));
    LocalMux I__2124 (
            .O(N__22950),
            .I(N__22947));
    Odrv12 I__2123 (
            .O(N__22947),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    InMux I__2122 (
            .O(N__22944),
            .I(N__22937));
    InMux I__2121 (
            .O(N__22943),
            .I(N__22937));
    InMux I__2120 (
            .O(N__22942),
            .I(N__22934));
    LocalMux I__2119 (
            .O(N__22937),
            .I(N__22931));
    LocalMux I__2118 (
            .O(N__22934),
            .I(N__22926));
    Span4Mux_v I__2117 (
            .O(N__22931),
            .I(N__22926));
    Span4Mux_v I__2116 (
            .O(N__22926),
            .I(N__22923));
    Odrv4 I__2115 (
            .O(N__22923),
            .I(\pid_alt.error_d_regZ0Z_6 ));
    CascadeMux I__2114 (
            .O(N__22920),
            .I(N__22914));
    InMux I__2113 (
            .O(N__22919),
            .I(N__22908));
    InMux I__2112 (
            .O(N__22918),
            .I(N__22908));
    InMux I__2111 (
            .O(N__22917),
            .I(N__22903));
    InMux I__2110 (
            .O(N__22914),
            .I(N__22903));
    InMux I__2109 (
            .O(N__22913),
            .I(N__22900));
    LocalMux I__2108 (
            .O(N__22908),
            .I(N__22897));
    LocalMux I__2107 (
            .O(N__22903),
            .I(N__22894));
    LocalMux I__2106 (
            .O(N__22900),
            .I(N__22889));
    Span4Mux_s2_h I__2105 (
            .O(N__22897),
            .I(N__22889));
    Odrv4 I__2104 (
            .O(N__22894),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    Odrv4 I__2103 (
            .O(N__22889),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    InMux I__2102 (
            .O(N__22884),
            .I(N__22880));
    CascadeMux I__2101 (
            .O(N__22883),
            .I(N__22875));
    LocalMux I__2100 (
            .O(N__22880),
            .I(N__22871));
    InMux I__2099 (
            .O(N__22879),
            .I(N__22866));
    InMux I__2098 (
            .O(N__22878),
            .I(N__22866));
    InMux I__2097 (
            .O(N__22875),
            .I(N__22861));
    InMux I__2096 (
            .O(N__22874),
            .I(N__22861));
    Odrv4 I__2095 (
            .O(N__22871),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__2094 (
            .O(N__22866),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__2093 (
            .O(N__22861),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    InMux I__2092 (
            .O(N__22854),
            .I(N__22851));
    LocalMux I__2091 (
            .O(N__22851),
            .I(N__22848));
    Span4Mux_v I__2090 (
            .O(N__22848),
            .I(N__22840));
    InMux I__2089 (
            .O(N__22847),
            .I(N__22835));
    InMux I__2088 (
            .O(N__22846),
            .I(N__22835));
    InMux I__2087 (
            .O(N__22845),
            .I(N__22828));
    InMux I__2086 (
            .O(N__22844),
            .I(N__22828));
    InMux I__2085 (
            .O(N__22843),
            .I(N__22828));
    Span4Mux_v I__2084 (
            .O(N__22840),
            .I(N__22825));
    LocalMux I__2083 (
            .O(N__22835),
            .I(N__22820));
    LocalMux I__2082 (
            .O(N__22828),
            .I(N__22820));
    Odrv4 I__2081 (
            .O(N__22825),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    Odrv12 I__2080 (
            .O(N__22820),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    CascadeMux I__2079 (
            .O(N__22815),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_ ));
    InMux I__2078 (
            .O(N__22812),
            .I(N__22809));
    LocalMux I__2077 (
            .O(N__22809),
            .I(N__22806));
    Span4Mux_h I__2076 (
            .O(N__22806),
            .I(N__22803));
    Span4Mux_v I__2075 (
            .O(N__22803),
            .I(N__22800));
    Odrv4 I__2074 (
            .O(N__22800),
            .I(\pid_alt.O_5_4 ));
    CascadeMux I__2073 (
            .O(N__22797),
            .I(N__22794));
    InMux I__2072 (
            .O(N__22794),
            .I(N__22788));
    InMux I__2071 (
            .O(N__22793),
            .I(N__22788));
    LocalMux I__2070 (
            .O(N__22788),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    CascadeMux I__2069 (
            .O(N__22785),
            .I(N__22780));
    CascadeMux I__2068 (
            .O(N__22784),
            .I(N__22777));
    CascadeMux I__2067 (
            .O(N__22783),
            .I(N__22774));
    InMux I__2066 (
            .O(N__22780),
            .I(N__22764));
    InMux I__2065 (
            .O(N__22777),
            .I(N__22764));
    InMux I__2064 (
            .O(N__22774),
            .I(N__22764));
    InMux I__2063 (
            .O(N__22773),
            .I(N__22764));
    LocalMux I__2062 (
            .O(N__22764),
            .I(N__22761));
    Span4Mux_s3_h I__2061 (
            .O(N__22761),
            .I(N__22758));
    Span4Mux_v I__2060 (
            .O(N__22758),
            .I(N__22754));
    InMux I__2059 (
            .O(N__22757),
            .I(N__22751));
    Odrv4 I__2058 (
            .O(N__22754),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    LocalMux I__2057 (
            .O(N__22751),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    CascadeMux I__2056 (
            .O(N__22746),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ));
    CEMux I__2055 (
            .O(N__22743),
            .I(N__22740));
    LocalMux I__2054 (
            .O(N__22740),
            .I(N__22737));
    Span4Mux_v I__2053 (
            .O(N__22737),
            .I(N__22734));
    Span4Mux_v I__2052 (
            .O(N__22734),
            .I(N__22731));
    Odrv4 I__2051 (
            .O(N__22731),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ));
    InMux I__2050 (
            .O(N__22728),
            .I(N__22725));
    LocalMux I__2049 (
            .O(N__22725),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ));
    InMux I__2048 (
            .O(N__22722),
            .I(N__22719));
    LocalMux I__2047 (
            .O(N__22719),
            .I(N__22716));
    Span4Mux_h I__2046 (
            .O(N__22716),
            .I(N__22713));
    Odrv4 I__2045 (
            .O(N__22713),
            .I(\pid_alt.O_4_5 ));
    InMux I__2044 (
            .O(N__22710),
            .I(N__22707));
    LocalMux I__2043 (
            .O(N__22707),
            .I(N__22704));
    Span4Mux_v I__2042 (
            .O(N__22704),
            .I(N__22701));
    Span4Mux_v I__2041 (
            .O(N__22701),
            .I(N__22698));
    Odrv4 I__2040 (
            .O(N__22698),
            .I(\pid_alt.O_3_4 ));
    InMux I__2039 (
            .O(N__22695),
            .I(N__22692));
    LocalMux I__2038 (
            .O(N__22692),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ));
    CascadeMux I__2037 (
            .O(N__22689),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ));
    InMux I__2036 (
            .O(N__22686),
            .I(N__22683));
    LocalMux I__2035 (
            .O(N__22683),
            .I(N__22680));
    Odrv4 I__2034 (
            .O(N__22680),
            .I(alt_kd_6));
    InMux I__2033 (
            .O(N__22677),
            .I(N__22674));
    LocalMux I__2032 (
            .O(N__22674),
            .I(N__22671));
    Odrv4 I__2031 (
            .O(N__22671),
            .I(alt_kd_4));
    InMux I__2030 (
            .O(N__22668),
            .I(N__22665));
    LocalMux I__2029 (
            .O(N__22665),
            .I(N__22662));
    Span4Mux_v I__2028 (
            .O(N__22662),
            .I(N__22659));
    Odrv4 I__2027 (
            .O(N__22659),
            .I(alt_kd_3));
    InMux I__2026 (
            .O(N__22656),
            .I(N__22653));
    LocalMux I__2025 (
            .O(N__22653),
            .I(N__22650));
    Span4Mux_s2_h I__2024 (
            .O(N__22650),
            .I(N__22647));
    Odrv4 I__2023 (
            .O(N__22647),
            .I(alt_kd_0));
    InMux I__2022 (
            .O(N__22644),
            .I(N__22641));
    LocalMux I__2021 (
            .O(N__22641),
            .I(N__22638));
    Span4Mux_s3_h I__2020 (
            .O(N__22638),
            .I(N__22635));
    Odrv4 I__2019 (
            .O(N__22635),
            .I(alt_ki_0));
    InMux I__2018 (
            .O(N__22632),
            .I(N__22629));
    LocalMux I__2017 (
            .O(N__22629),
            .I(N__22626));
    Span4Mux_v I__2016 (
            .O(N__22626),
            .I(N__22623));
    Odrv4 I__2015 (
            .O(N__22623),
            .I(alt_ki_2));
    CEMux I__2014 (
            .O(N__22620),
            .I(N__22617));
    LocalMux I__2013 (
            .O(N__22617),
            .I(N__22612));
    CEMux I__2012 (
            .O(N__22616),
            .I(N__22609));
    CEMux I__2011 (
            .O(N__22615),
            .I(N__22606));
    Span4Mux_s3_h I__2010 (
            .O(N__22612),
            .I(N__22603));
    LocalMux I__2009 (
            .O(N__22609),
            .I(N__22598));
    LocalMux I__2008 (
            .O(N__22606),
            .I(N__22598));
    Odrv4 I__2007 (
            .O(N__22603),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    Odrv4 I__2006 (
            .O(N__22598),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    InMux I__2005 (
            .O(N__22593),
            .I(N__22590));
    LocalMux I__2004 (
            .O(N__22590),
            .I(N__22587));
    Span4Mux_v I__2003 (
            .O(N__22587),
            .I(N__22584));
    Odrv4 I__2002 (
            .O(N__22584),
            .I(\pid_alt.g0_4_0 ));
    InMux I__2001 (
            .O(N__22581),
            .I(N__22578));
    LocalMux I__2000 (
            .O(N__22578),
            .I(N__22575));
    Odrv4 I__1999 (
            .O(N__22575),
            .I(\pid_alt.O_5_18 ));
    InMux I__1998 (
            .O(N__22572),
            .I(N__22569));
    LocalMux I__1997 (
            .O(N__22569),
            .I(N__22566));
    Odrv4 I__1996 (
            .O(N__22566),
            .I(\pid_alt.O_5_21 ));
    InMux I__1995 (
            .O(N__22563),
            .I(N__22560));
    LocalMux I__1994 (
            .O(N__22560),
            .I(N__22557));
    Odrv4 I__1993 (
            .O(N__22557),
            .I(\pid_alt.O_5_19 ));
    InMux I__1992 (
            .O(N__22554),
            .I(N__22551));
    LocalMux I__1991 (
            .O(N__22551),
            .I(\pid_alt.O_5_14 ));
    InMux I__1990 (
            .O(N__22548),
            .I(N__22545));
    LocalMux I__1989 (
            .O(N__22545),
            .I(N__22542));
    Odrv4 I__1988 (
            .O(N__22542),
            .I(\pid_alt.O_5_23 ));
    InMux I__1987 (
            .O(N__22539),
            .I(N__22536));
    LocalMux I__1986 (
            .O(N__22536),
            .I(N__22533));
    Odrv4 I__1985 (
            .O(N__22533),
            .I(\pid_alt.O_5_16 ));
    InMux I__1984 (
            .O(N__22530),
            .I(N__22527));
    LocalMux I__1983 (
            .O(N__22527),
            .I(\pid_alt.O_5_12 ));
    InMux I__1982 (
            .O(N__22524),
            .I(N__22521));
    LocalMux I__1981 (
            .O(N__22521),
            .I(\pid_alt.O_5_13 ));
    InMux I__1980 (
            .O(N__22518),
            .I(N__22515));
    LocalMux I__1979 (
            .O(N__22515),
            .I(N__22512));
    Odrv4 I__1978 (
            .O(N__22512),
            .I(\pid_alt.O_5_24 ));
    InMux I__1977 (
            .O(N__22509),
            .I(N__22506));
    LocalMux I__1976 (
            .O(N__22506),
            .I(N__22503));
    Odrv4 I__1975 (
            .O(N__22503),
            .I(\pid_alt.O_5_7 ));
    InMux I__1974 (
            .O(N__22500),
            .I(N__22497));
    LocalMux I__1973 (
            .O(N__22497),
            .I(N__22494));
    Odrv4 I__1972 (
            .O(N__22494),
            .I(\pid_alt.O_5_8 ));
    InMux I__1971 (
            .O(N__22491),
            .I(N__22488));
    LocalMux I__1970 (
            .O(N__22488),
            .I(N__22485));
    Span4Mux_v I__1969 (
            .O(N__22485),
            .I(N__22482));
    Span4Mux_v I__1968 (
            .O(N__22482),
            .I(N__22479));
    Span4Mux_v I__1967 (
            .O(N__22479),
            .I(N__22476));
    Odrv4 I__1966 (
            .O(N__22476),
            .I(\pid_alt.O_4_8 ));
    InMux I__1965 (
            .O(N__22473),
            .I(N__22470));
    LocalMux I__1964 (
            .O(N__22470),
            .I(N__22467));
    Odrv4 I__1963 (
            .O(N__22467),
            .I(\pid_alt.O_5_11 ));
    InMux I__1962 (
            .O(N__22464),
            .I(N__22461));
    LocalMux I__1961 (
            .O(N__22461),
            .I(N__22458));
    Span4Mux_h I__1960 (
            .O(N__22458),
            .I(N__22455));
    Odrv4 I__1959 (
            .O(N__22455),
            .I(\pid_alt.O_5_22 ));
    InMux I__1958 (
            .O(N__22452),
            .I(N__22449));
    LocalMux I__1957 (
            .O(N__22449),
            .I(N__22446));
    Odrv4 I__1956 (
            .O(N__22446),
            .I(\pid_alt.O_5_15 ));
    InMux I__1955 (
            .O(N__22443),
            .I(N__22440));
    LocalMux I__1954 (
            .O(N__22440),
            .I(N__22437));
    Odrv4 I__1953 (
            .O(N__22437),
            .I(\pid_alt.O_5_17 ));
    InMux I__1952 (
            .O(N__22434),
            .I(N__22431));
    LocalMux I__1951 (
            .O(N__22431),
            .I(N__22428));
    Odrv4 I__1950 (
            .O(N__22428),
            .I(\pid_alt.O_5_20 ));
    InMux I__1949 (
            .O(N__22425),
            .I(N__22422));
    LocalMux I__1948 (
            .O(N__22422),
            .I(N__22419));
    Span4Mux_h I__1947 (
            .O(N__22419),
            .I(N__22416));
    Span4Mux_v I__1946 (
            .O(N__22416),
            .I(N__22413));
    Odrv4 I__1945 (
            .O(N__22413),
            .I(\pid_alt.O_5_5 ));
    InMux I__1944 (
            .O(N__22410),
            .I(N__22407));
    LocalMux I__1943 (
            .O(N__22407),
            .I(N__22404));
    Odrv4 I__1942 (
            .O(N__22404),
            .I(\pid_front.O_0_8 ));
    CascadeMux I__1941 (
            .O(N__22401),
            .I(\Commands_frame_decoder.source_CH1data8_cascade_ ));
    InMux I__1940 (
            .O(N__22398),
            .I(N__22389));
    InMux I__1939 (
            .O(N__22397),
            .I(N__22389));
    InMux I__1938 (
            .O(N__22396),
            .I(N__22389));
    LocalMux I__1937 (
            .O(N__22389),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    InMux I__1936 (
            .O(N__22386),
            .I(N__22383));
    LocalMux I__1935 (
            .O(N__22383),
            .I(N__22380));
    Odrv4 I__1934 (
            .O(N__22380),
            .I(\pid_front.O_0_22 ));
    InMux I__1933 (
            .O(N__22377),
            .I(N__22374));
    LocalMux I__1932 (
            .O(N__22374),
            .I(N__22371));
    Odrv4 I__1931 (
            .O(N__22371),
            .I(\pid_front.O_0_23 ));
    InMux I__1930 (
            .O(N__22368),
            .I(N__22365));
    LocalMux I__1929 (
            .O(N__22365),
            .I(N__22362));
    Odrv4 I__1928 (
            .O(N__22362),
            .I(\pid_front.O_0_24 ));
    InMux I__1927 (
            .O(N__22359),
            .I(N__22356));
    LocalMux I__1926 (
            .O(N__22356),
            .I(\pid_front.O_0_21 ));
    InMux I__1925 (
            .O(N__22353),
            .I(N__22350));
    LocalMux I__1924 (
            .O(N__22350),
            .I(\pid_front.O_0_20 ));
    InMux I__1923 (
            .O(N__22347),
            .I(N__22344));
    LocalMux I__1922 (
            .O(N__22344),
            .I(\pid_front.O_0_14 ));
    InMux I__1921 (
            .O(N__22341),
            .I(N__22338));
    LocalMux I__1920 (
            .O(N__22338),
            .I(\pid_front.O_0_10 ));
    InMux I__1919 (
            .O(N__22335),
            .I(N__22332));
    LocalMux I__1918 (
            .O(N__22332),
            .I(\pid_front.O_0_13 ));
    InMux I__1917 (
            .O(N__22329),
            .I(N__22326));
    LocalMux I__1916 (
            .O(N__22326),
            .I(N__22323));
    Span4Mux_h I__1915 (
            .O(N__22323),
            .I(N__22320));
    Span4Mux_v I__1914 (
            .O(N__22320),
            .I(N__22317));
    Odrv4 I__1913 (
            .O(N__22317),
            .I(\pid_alt.O_5_6 ));
    InMux I__1912 (
            .O(N__22314),
            .I(N__22311));
    LocalMux I__1911 (
            .O(N__22311),
            .I(\pid_alt.N_5 ));
    InMux I__1910 (
            .O(N__22308),
            .I(N__22305));
    LocalMux I__1909 (
            .O(N__22305),
            .I(\pid_alt.N_1672_0 ));
    InMux I__1908 (
            .O(N__22302),
            .I(N__22299));
    LocalMux I__1907 (
            .O(N__22299),
            .I(N__22296));
    Odrv4 I__1906 (
            .O(N__22296),
            .I(\pid_front.O_0_16 ));
    InMux I__1905 (
            .O(N__22293),
            .I(N__22290));
    LocalMux I__1904 (
            .O(N__22290),
            .I(N__22287));
    Odrv4 I__1903 (
            .O(N__22287),
            .I(\pid_front.O_0_17 ));
    InMux I__1902 (
            .O(N__22284),
            .I(N__22281));
    LocalMux I__1901 (
            .O(N__22281),
            .I(N__22278));
    Odrv4 I__1900 (
            .O(N__22278),
            .I(\pid_front.O_0_18 ));
    InMux I__1899 (
            .O(N__22275),
            .I(N__22272));
    LocalMux I__1898 (
            .O(N__22272),
            .I(N__22269));
    Odrv4 I__1897 (
            .O(N__22269),
            .I(\pid_front.O_0_19 ));
    InMux I__1896 (
            .O(N__22266),
            .I(N__22263));
    LocalMux I__1895 (
            .O(N__22263),
            .I(\pid_front.O_0_12 ));
    InMux I__1894 (
            .O(N__22260),
            .I(N__22257));
    LocalMux I__1893 (
            .O(N__22257),
            .I(\pid_front.O_0_7 ));
    InMux I__1892 (
            .O(N__22254),
            .I(N__22251));
    LocalMux I__1891 (
            .O(N__22251),
            .I(\pid_alt.N_3_1 ));
    CascadeMux I__1890 (
            .O(N__22248),
            .I(N__22245));
    InMux I__1889 (
            .O(N__22245),
            .I(N__22242));
    LocalMux I__1888 (
            .O(N__22242),
            .I(\pid_alt.N_1668_1 ));
    InMux I__1887 (
            .O(N__22239),
            .I(N__22236));
    LocalMux I__1886 (
            .O(N__22236),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2 ));
    InMux I__1885 (
            .O(N__22233),
            .I(N__22230));
    LocalMux I__1884 (
            .O(N__22230),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ));
    CascadeMux I__1883 (
            .O(N__22227),
            .I(\pid_alt.N_1674_0_cascade_ ));
    InMux I__1882 (
            .O(N__22224),
            .I(N__22221));
    LocalMux I__1881 (
            .O(N__22221),
            .I(\pid_alt.N_1666_i_0 ));
    InMux I__1880 (
            .O(N__22218),
            .I(N__22215));
    LocalMux I__1879 (
            .O(N__22215),
            .I(\pid_alt.N_3_0 ));
    CascadeMux I__1878 (
            .O(N__22212),
            .I(N__22209));
    InMux I__1877 (
            .O(N__22209),
            .I(N__22206));
    LocalMux I__1876 (
            .O(N__22206),
            .I(\pid_alt.N_1668_0 ));
    InMux I__1875 (
            .O(N__22203),
            .I(N__22200));
    LocalMux I__1874 (
            .O(N__22200),
            .I(\pid_alt.O_4_19 ));
    InMux I__1873 (
            .O(N__22197),
            .I(N__22194));
    LocalMux I__1872 (
            .O(N__22194),
            .I(\pid_alt.O_4_6 ));
    InMux I__1871 (
            .O(N__22191),
            .I(N__22188));
    LocalMux I__1870 (
            .O(N__22188),
            .I(\pid_alt.O_4_21 ));
    InMux I__1869 (
            .O(N__22185),
            .I(N__22182));
    LocalMux I__1868 (
            .O(N__22182),
            .I(\pid_alt.O_4_13 ));
    InMux I__1867 (
            .O(N__22179),
            .I(N__22176));
    LocalMux I__1866 (
            .O(N__22176),
            .I(\pid_alt.O_4_12 ));
    CascadeMux I__1865 (
            .O(N__22173),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_ ));
    InMux I__1864 (
            .O(N__22170),
            .I(N__22167));
    LocalMux I__1863 (
            .O(N__22167),
            .I(\pid_alt.N_1666_i_1 ));
    InMux I__1862 (
            .O(N__22164),
            .I(N__22161));
    LocalMux I__1861 (
            .O(N__22161),
            .I(N__22158));
    Odrv4 I__1860 (
            .O(N__22158),
            .I(\pid_alt.O_4_23 ));
    InMux I__1859 (
            .O(N__22155),
            .I(N__22152));
    LocalMux I__1858 (
            .O(N__22152),
            .I(N__22149));
    Odrv4 I__1857 (
            .O(N__22149),
            .I(\pid_alt.O_4_22 ));
    InMux I__1856 (
            .O(N__22146),
            .I(N__22143));
    LocalMux I__1855 (
            .O(N__22143),
            .I(\pid_alt.O_4_10 ));
    InMux I__1854 (
            .O(N__22140),
            .I(N__22137));
    LocalMux I__1853 (
            .O(N__22137),
            .I(\pid_alt.O_4_14 ));
    InMux I__1852 (
            .O(N__22134),
            .I(N__22131));
    LocalMux I__1851 (
            .O(N__22131),
            .I(\pid_alt.O_4_11 ));
    InMux I__1850 (
            .O(N__22128),
            .I(N__22125));
    LocalMux I__1849 (
            .O(N__22125),
            .I(N__22122));
    Odrv4 I__1848 (
            .O(N__22122),
            .I(\pid_alt.O_4_17 ));
    InMux I__1847 (
            .O(N__22119),
            .I(N__22116));
    LocalMux I__1846 (
            .O(N__22116),
            .I(\pid_alt.O_4_16 ));
    InMux I__1845 (
            .O(N__22113),
            .I(N__22110));
    LocalMux I__1844 (
            .O(N__22110),
            .I(\pid_alt.O_4_20 ));
    InMux I__1843 (
            .O(N__22107),
            .I(N__22104));
    LocalMux I__1842 (
            .O(N__22104),
            .I(\pid_alt.O_4_18 ));
    InMux I__1841 (
            .O(N__22101),
            .I(N__22098));
    LocalMux I__1840 (
            .O(N__22098),
            .I(alt_kd_5));
    InMux I__1839 (
            .O(N__22095),
            .I(N__22092));
    LocalMux I__1838 (
            .O(N__22092),
            .I(N__22089));
    Span4Mux_s2_h I__1837 (
            .O(N__22089),
            .I(N__22086));
    Odrv4 I__1836 (
            .O(N__22086),
            .I(alt_ki_6));
    InMux I__1835 (
            .O(N__22083),
            .I(N__22080));
    LocalMux I__1834 (
            .O(N__22080),
            .I(N__22077));
    Span4Mux_s2_h I__1833 (
            .O(N__22077),
            .I(N__22074));
    Odrv4 I__1832 (
            .O(N__22074),
            .I(alt_ki_7));
    InMux I__1831 (
            .O(N__22071),
            .I(N__22068));
    LocalMux I__1830 (
            .O(N__22068),
            .I(N__22065));
    Span4Mux_s2_h I__1829 (
            .O(N__22065),
            .I(N__22062));
    Odrv4 I__1828 (
            .O(N__22062),
            .I(alt_ki_1));
    InMux I__1827 (
            .O(N__22059),
            .I(N__22056));
    LocalMux I__1826 (
            .O(N__22056),
            .I(N__22053));
    Odrv4 I__1825 (
            .O(N__22053),
            .I(alt_ki_3));
    InMux I__1824 (
            .O(N__22050),
            .I(N__22047));
    LocalMux I__1823 (
            .O(N__22047),
            .I(N__22044));
    Odrv4 I__1822 (
            .O(N__22044),
            .I(alt_ki_4));
    InMux I__1821 (
            .O(N__22041),
            .I(N__22038));
    LocalMux I__1820 (
            .O(N__22038),
            .I(N__22035));
    Span4Mux_s2_h I__1819 (
            .O(N__22035),
            .I(N__22032));
    Odrv4 I__1818 (
            .O(N__22032),
            .I(alt_ki_5));
    InMux I__1817 (
            .O(N__22029),
            .I(N__22026));
    LocalMux I__1816 (
            .O(N__22026),
            .I(\pid_alt.O_4_9 ));
    InMux I__1815 (
            .O(N__22023),
            .I(N__22020));
    LocalMux I__1814 (
            .O(N__22020),
            .I(N__22017));
    Odrv4 I__1813 (
            .O(N__22017),
            .I(\pid_alt.O_4_24 ));
    InMux I__1812 (
            .O(N__22014),
            .I(N__22011));
    LocalMux I__1811 (
            .O(N__22011),
            .I(\pid_alt.O_3_21 ));
    InMux I__1810 (
            .O(N__22008),
            .I(N__22005));
    LocalMux I__1809 (
            .O(N__22005),
            .I(\pid_alt.O_3_22 ));
    InMux I__1808 (
            .O(N__22002),
            .I(N__21999));
    LocalMux I__1807 (
            .O(N__21999),
            .I(\pid_alt.O_3_23 ));
    InMux I__1806 (
            .O(N__21996),
            .I(N__21993));
    LocalMux I__1805 (
            .O(N__21993),
            .I(\pid_alt.O_3_6 ));
    InMux I__1804 (
            .O(N__21990),
            .I(N__21987));
    LocalMux I__1803 (
            .O(N__21987),
            .I(N__21984));
    Odrv4 I__1802 (
            .O(N__21984),
            .I(\pid_alt.O_3_24 ));
    InMux I__1801 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__1800 (
            .O(N__21978),
            .I(\pid_alt.O_3_7 ));
    InMux I__1799 (
            .O(N__21975),
            .I(N__21972));
    LocalMux I__1798 (
            .O(N__21972),
            .I(\pid_alt.O_3_9 ));
    InMux I__1797 (
            .O(N__21969),
            .I(N__21966));
    LocalMux I__1796 (
            .O(N__21966),
            .I(alt_kd_7));
    InMux I__1795 (
            .O(N__21963),
            .I(N__21960));
    LocalMux I__1794 (
            .O(N__21960),
            .I(alt_kd_2));
    InMux I__1793 (
            .O(N__21957),
            .I(N__21954));
    LocalMux I__1792 (
            .O(N__21954),
            .I(alt_kd_1));
    InMux I__1791 (
            .O(N__21951),
            .I(N__21948));
    LocalMux I__1790 (
            .O(N__21948),
            .I(N__21945));
    Odrv4 I__1789 (
            .O(N__21945),
            .I(\pid_alt.O_3_10 ));
    InMux I__1788 (
            .O(N__21942),
            .I(N__21939));
    LocalMux I__1787 (
            .O(N__21939),
            .I(\pid_alt.O_3_5 ));
    InMux I__1786 (
            .O(N__21936),
            .I(N__21933));
    LocalMux I__1785 (
            .O(N__21933),
            .I(\pid_alt.O_3_14 ));
    InMux I__1784 (
            .O(N__21930),
            .I(N__21927));
    LocalMux I__1783 (
            .O(N__21927),
            .I(\pid_alt.O_3_15 ));
    InMux I__1782 (
            .O(N__21924),
            .I(N__21921));
    LocalMux I__1781 (
            .O(N__21921),
            .I(N__21918));
    Odrv4 I__1780 (
            .O(N__21918),
            .I(\pid_alt.O_3_16 ));
    InMux I__1779 (
            .O(N__21915),
            .I(N__21912));
    LocalMux I__1778 (
            .O(N__21912),
            .I(N__21909));
    Odrv4 I__1777 (
            .O(N__21909),
            .I(\pid_alt.O_3_17 ));
    InMux I__1776 (
            .O(N__21906),
            .I(N__21903));
    LocalMux I__1775 (
            .O(N__21903),
            .I(N__21900));
    Odrv4 I__1774 (
            .O(N__21900),
            .I(\pid_alt.O_3_18 ));
    InMux I__1773 (
            .O(N__21897),
            .I(N__21894));
    LocalMux I__1772 (
            .O(N__21894),
            .I(N__21891));
    Odrv4 I__1771 (
            .O(N__21891),
            .I(\pid_alt.O_3_19 ));
    InMux I__1770 (
            .O(N__21888),
            .I(N__21885));
    LocalMux I__1769 (
            .O(N__21885),
            .I(N__21882));
    Odrv4 I__1768 (
            .O(N__21882),
            .I(\pid_alt.O_3_20 ));
    IoInMux I__1767 (
            .O(N__21879),
            .I(N__21876));
    LocalMux I__1766 (
            .O(N__21876),
            .I(N__21873));
    IoSpan4Mux I__1765 (
            .O(N__21873),
            .I(N__21870));
    Span4Mux_s2_v I__1764 (
            .O(N__21870),
            .I(N__21867));
    Sp12to4 I__1763 (
            .O(N__21867),
            .I(N__21864));
    Span12Mux_v I__1762 (
            .O(N__21864),
            .I(N__21861));
    Span12Mux_v I__1761 (
            .O(N__21861),
            .I(N__21858));
    Odrv12 I__1760 (
            .O(N__21858),
            .I(\Pc2drone_pll_inst.clk_system_pll ));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_2_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_20_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_2_20_0_));
    defparam IN_MUX_bfv_20_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_9_0_));
    defparam IN_MUX_bfv_20_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_10_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_cry_5 ),
            .carryinitout(bfn_20_10_0_));
    defparam IN_MUX_bfv_20_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_11_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_cry_13 ),
            .carryinitout(bfn_20_11_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_cry_5 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_12_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_23_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_cry_13 ),
            .carryinitout(bfn_12_23_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_21_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_17_0_));
    defparam IN_MUX_bfv_21_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_18_0_ (
            .carryinitin(\pid_side.error_cry_3_0 ),
            .carryinitout(bfn_21_18_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\pid_front.error_cry_3_0 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_8_6_0_));
    ICE_GB \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0  (
            .USERSIGNALTOGLOBALBUFFER(N__41964),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_419_g ));
    ICE_GB \pid_alt.state_RNICP2N1_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__47781),
            .GLOBALBUFFEROUTPUT(\pid_alt.N_664_0_g ));
    ICE_GB \Pc2drone_pll_inst.PLLOUTCORE_derived_clock_RNI5FOA  (
            .USERSIGNALTOGLOBALBUFFER(N__21879),
            .GLOBALBUFFEROUTPUT(clk_system_pll_g));
    ICE_GB \reset_module_System.reset_RNITC69_0  (
            .USERSIGNALTOGLOBALBUFFER(N__49272),
            .GLOBALBUFFEROUTPUT(N_665_g));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__44971),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB \pid_front.state_RNIPKTD_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__31203),
            .GLOBALBUFFEROUTPUT(\pid_front.state_0_g_0 ));
    ICE_GB \pid_side.state_RNIL5IF_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__35586),
            .GLOBALBUFFEROUTPUT(\pid_side.state_0_g_0 ));
    ICE_GB \pid_alt.state_RNIH1EN_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__39351),
            .GLOBALBUFFEROUTPUT(\pid_alt.state_0_g_0 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_6_LC_1_4_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_6_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21951),
            .lcout(\pid_alt.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59139),
            .ce(N__24449),
            .sr(N__58219));
    defparam \pid_alt.error_d_reg_esr_1_LC_1_5_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_1_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21942),
            .lcout(\pid_alt.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_10_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21936),
            .lcout(\pid_alt.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_11_LC_1_5_2  (
            .in0(N__21930),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_12_LC_1_5_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_5_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_12_LC_1_5_3  (
            .in0(N__21924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_13_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21915),
            .lcout(\pid_alt.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_14_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21906),
            .lcout(\pid_alt.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_15_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21897),
            .lcout(\pid_alt.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_16_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21888),
            .lcout(\pid_alt.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59152),
            .ce(N__24450),
            .sr(N__58218));
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_17_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22014),
            .lcout(\pid_alt.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59165),
            .ce(N__24451),
            .sr(N__58217));
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_18_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22008),
            .lcout(\pid_alt.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59165),
            .ce(N__24451),
            .sr(N__58217));
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_19_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22002),
            .lcout(\pid_alt.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59165),
            .ce(N__24451),
            .sr(N__58217));
    defparam \pid_alt.error_d_reg_esr_2_LC_1_6_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_2_LC_1_6_3  (
            .in0(N__21996),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59165),
            .ce(N__24451),
            .sr(N__58217));
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_20_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21990),
            .lcout(\pid_alt.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59165),
            .ce(N__24451),
            .sr(N__58217));
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_3_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21981),
            .lcout(\pid_alt.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59165),
            .ce(N__24451),
            .sr(N__58217));
    defparam \pid_alt.error_d_reg_esr_5_LC_1_6_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_5_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21975),
            .lcout(\pid_alt.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59165),
            .ce(N__24451),
            .sr(N__58217));
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_1_7_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_1_7_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_7_LC_1_7_0  (
            .in0(N__58357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55566),
            .lcout(alt_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59179),
            .ce(N__24282),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_1_7_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_1_7_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_2_LC_1_7_2  (
            .in0(N__58355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56111),
            .lcout(alt_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59179),
            .ce(N__24282),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_1_7_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_1_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_1_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__56278),
            .in2(_gnd_net_),
            .in3(N__58354),
            .lcout(alt_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59179),
            .ce(N__24282),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_1_7_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_1_7_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_5_LC_1_7_6  (
            .in0(N__58356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55899),
            .lcout(alt_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59179),
            .ce(N__24282),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_1_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_1_8_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_6_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__55732),
            .in2(_gnd_net_),
            .in3(N__58352),
            .lcout(alt_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59194),
            .ce(N__22615),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7  (
            .in0(N__58353),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55565),
            .lcout(alt_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59194),
            .ce(N__22615),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_1_9_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_1_9_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_1_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__56242),
            .in2(_gnd_net_),
            .in3(N__58346),
            .lcout(alt_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59206),
            .ce(N__22620),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_1_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_1_9_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_1_9_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_3_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__55354),
            .in2(_gnd_net_),
            .in3(N__58347),
            .lcout(alt_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59206),
            .ce(N__22620),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_1_9_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_1_9_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_1_9_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_4_LC_1_9_4  (
            .in0(N__58348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53360),
            .lcout(alt_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59206),
            .ce(N__22620),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_1_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_1_9_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_5_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__55876),
            .in2(_gnd_net_),
            .in3(N__58349),
            .lcout(alt_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59206),
            .ce(N__22620),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_5_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22029),
            .lcout(\pid_alt.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_20_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22023),
            .lcout(\pid_alt.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_19_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22164),
            .lcout(\pid_alt.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_18_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22155),
            .lcout(\pid_alt.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_6_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22146),
            .lcout(\pid_alt.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_10_LC_1_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_10_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22140),
            .lcout(\pid_alt.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_7_LC_1_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_7_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22134),
            .lcout(\pid_alt.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_13_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22128),
            .lcout(\pid_alt.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59221),
            .ce(N__24453),
            .sr(N__58215));
    defparam \pid_alt.error_i_reg_esr_12_LC_1_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_12_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22119),
            .lcout(\pid_alt.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_16_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22113),
            .lcout(\pid_alt.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_i_reg_esr_14_LC_1_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_14_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22107),
            .lcout(\pid_alt.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_15_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22203),
            .lcout(\pid_alt.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_2_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22197),
            .lcout(\pid_alt.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_17_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22191),
            .lcout(\pid_alt.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_i_reg_esr_9_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_9_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22185),
            .lcout(\pid_alt.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22179),
            .lcout(\pid_alt.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59237),
            .ce(N__24454),
            .sr(N__58213));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_12_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_12_7  (
            .in0(N__23067),
            .in1(N__23010),
            .in2(_gnd_net_),
            .in3(N__23032),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_13_0 .LUT_INIT=16'b0011000001110001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_13_0  (
            .in0(N__22170),
            .in1(N__22239),
            .in2(N__22248),
            .in3(N__22254),
            .lcout(),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_13_1  (
            .in0(N__22728),
            .in1(N__25869),
            .in2(N__22173),
            .in3(N__22233),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_13_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__23229),
            .in2(_gnd_net_),
            .in3(N__24389),
            .lcout(\pid_alt.N_1666_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_13_3  (
            .in0(N__23195),
            .in1(N__23152),
            .in2(_gnd_net_),
            .in3(N__23106),
            .lcout(\pid_alt.N_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_13_4 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_13_4  (
            .in0(N__23107),
            .in1(_gnd_net_),
            .in2(N__23162),
            .in3(N__23196),
            .lcout(\pid_alt.N_1668_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_13_5  (
            .in0(N__22918),
            .in1(N__22874),
            .in2(_gnd_net_),
            .in3(N__22843),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_13_6 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_13_6  (
            .in0(N__22844),
            .in1(_gnd_net_),
            .in2(N__22883),
            .in3(N__22919),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_2_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22845),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59270),
            .ce(N__27612),
            .sr(N__57531));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_14_0 .LUT_INIT=16'b0011000001110001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_14_0  (
            .in0(N__22224),
            .in1(N__22314),
            .in2(N__22212),
            .in3(N__22218),
            .lcout(),
            .ltout(\pid_alt.N_1674_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_14_1 .LUT_INIT=16'b1110100011010100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_14_1  (
            .in0(N__22593),
            .in1(N__22308),
            .in2(N__22227),
            .in3(N__24661),
            .lcout(\pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_14_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__23228),
            .in2(_gnd_net_),
            .in3(N__24390),
            .lcout(\pid_alt.N_1666_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_14_3  (
            .in0(N__23191),
            .in1(N__23156),
            .in2(_gnd_net_),
            .in3(N__23118),
            .lcout(\pid_alt.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_14_4 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_14_4  (
            .in0(N__23119),
            .in1(_gnd_net_),
            .in2(N__23163),
            .in3(N__23192),
            .lcout(\pid_alt.N_1668_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_14_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_14_5  (
            .in0(N__22878),
            .in1(_gnd_net_),
            .in2(N__22920),
            .in3(N__22846),
            .lcout(\pid_alt.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_14_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_14_6  (
            .in0(N__22847),
            .in1(N__22917),
            .in2(_gnd_net_),
            .in3(N__22879),
            .lcout(\pid_alt.N_1672_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_1_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_1_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_1_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23120),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59283),
            .ce(N__27609),
            .sr(N__57538));
    defparam \pid_front.error_p_reg_esr_12_LC_1_15_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_12_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_12_LC_1_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_12_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22302),
            .lcout(\pid_front.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_13_LC_1_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_13_LC_1_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_13_LC_1_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_13_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22293),
            .lcout(\pid_front.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_14_LC_1_15_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_14_LC_1_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_14_LC_1_15_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_p_reg_esr_14_LC_1_15_2  (
            .in0(N__22284),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_15_LC_1_15_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_15_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_15_LC_1_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_p_reg_esr_15_LC_1_15_3  (
            .in0(N__22275),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_8_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22266),
            .lcout(\pid_front.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_3_LC_1_15_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_3_LC_1_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_3_LC_1_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_3_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22260),
            .lcout(\pid_front.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_18_LC_1_15_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_18_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_18_LC_1_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_18_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22386),
            .lcout(\pid_front.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_19_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22377),
            .lcout(\pid_front.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59293),
            .ce(N__58537),
            .sr(N__58211));
    defparam \pid_front.error_p_reg_esr_20_LC_1_16_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_20_LC_1_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_20_LC_1_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_20_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22368),
            .lcout(\pid_front.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59303),
            .ce(N__58539),
            .sr(N__58209));
    defparam \pid_front.error_p_reg_esr_17_LC_1_16_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_17_LC_1_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_17_LC_1_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_17_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22359),
            .lcout(\pid_front.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59303),
            .ce(N__58539),
            .sr(N__58209));
    defparam \pid_front.error_p_reg_esr_16_LC_1_16_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_16_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_16_LC_1_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_16_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22353),
            .lcout(\pid_front.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59303),
            .ce(N__58539),
            .sr(N__58209));
    defparam \pid_front.error_p_reg_esr_10_LC_1_16_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_10_LC_1_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_10_LC_1_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_10_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22347),
            .lcout(\pid_front.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59303),
            .ce(N__58539),
            .sr(N__58209));
    defparam \pid_front.error_p_reg_esr_6_LC_1_16_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_6_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_6_LC_1_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_6_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22341),
            .lcout(\pid_front.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59303),
            .ce(N__58539),
            .sr(N__58209));
    defparam \pid_front.error_p_reg_esr_9_LC_1_16_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_9_LC_1_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_9_LC_1_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_9_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22335),
            .lcout(\pid_front.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59303),
            .ce(N__58539),
            .sr(N__58209));
    defparam \pid_alt.error_p_reg_esr_2_LC_1_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_2_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22329),
            .lcout(\pid_alt.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59310),
            .ce(N__24457),
            .sr(N__58208));
    defparam \pid_alt.error_p_reg_esr_1_LC_1_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_1_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22425),
            .lcout(\pid_alt.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59310),
            .ce(N__24457),
            .sr(N__58208));
    defparam \pid_front.error_p_reg_esr_4_LC_1_18_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_4_LC_1_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_4_LC_1_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_4_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22410),
            .lcout(\pid_front.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59314),
            .ce(N__58538),
            .sr(N__58207));
    defparam \Commands_frame_decoder.source_CH1data_3_LC_1_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_1_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_1_19_0 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_3_LC_1_19_0  (
            .in0(N__22398),
            .in1(N__55373),
            .in2(N__22785),
            .in3(N__23747),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59318),
            .ce(),
            .sr(N__57580));
    defparam \Commands_frame_decoder.source_CH1data_1_LC_1_19_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_1_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_1_19_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_1_LC_1_19_2  (
            .in0(N__22396),
            .in1(N__56304),
            .in2(N__22783),
            .in3(N__23870),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59318),
            .ce(),
            .sr(N__57580));
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_1_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_1_19_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_LC_1_19_4  (
            .in0(N__29166),
            .in1(N__24411),
            .in2(N__53405),
            .in3(N__55716),
            .lcout(\Commands_frame_decoder.source_CH1data8 ),
            .ltout(\Commands_frame_decoder.source_CH1data8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_0_LC_1_19_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_1_19_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_1_19_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \Commands_frame_decoder.source_CH1data_0_LC_1_19_5  (
            .in0(N__23934),
            .in1(N__56486),
            .in2(N__22401),
            .in3(N__22773),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59318),
            .ce(),
            .sr(N__57580));
    defparam \Commands_frame_decoder.source_CH1data_2_LC_1_19_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_1_19_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_1_19_6 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_2_LC_1_19_6  (
            .in0(N__22397),
            .in1(N__56139),
            .in2(N__22784),
            .in3(N__23810),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59318),
            .ce(),
            .sr(N__57580));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_1_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_1_20_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_1_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53401),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59321),
            .ce(N__22743),
            .sr(N__57589));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_1_20_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_1_20_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_1_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55927),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59321),
            .ce(N__22743),
            .sr(N__57589));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_1_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_1_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_1_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55750),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59321),
            .ce(N__22743),
            .sr(N__57589));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_1_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_1_20_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_1_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_1_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55583),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59321),
            .ce(N__22743),
            .sr(N__57589));
    defparam \pid_alt.error_p_reg_esr_3_LC_1_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_3_LC_1_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22509),
            .lcout(\pid_alt.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59326),
            .ce(N__24458),
            .sr(N__58205));
    defparam \pid_alt.error_p_reg_esr_4_LC_1_21_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_4_LC_1_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22500),
            .lcout(\pid_alt.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59326),
            .ce(N__24458),
            .sr(N__58205));
    defparam \pid_alt.error_i_reg_esr_4_LC_1_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_4_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22491),
            .lcout(\pid_alt.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59331),
            .ce(N__24459),
            .sr(N__58203));
    defparam \pid_alt.error_p_reg_esr_7_LC_1_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_22_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_7_LC_1_22_1  (
            .in0(N__22473),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59331),
            .ce(N__24459),
            .sr(N__58203));
    defparam \pid_alt.error_p_reg_esr_18_LC_1_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_18_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22464),
            .lcout(\pid_alt.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59331),
            .ce(N__24459),
            .sr(N__58203));
    defparam \pid_alt.error_p_reg_esr_11_LC_1_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_11_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22452),
            .lcout(\pid_alt.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59331),
            .ce(N__24459),
            .sr(N__58203));
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_13_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22443),
            .lcout(\pid_alt.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59331),
            .ce(N__24459),
            .sr(N__58203));
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_16_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22434),
            .lcout(\pid_alt.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59331),
            .ce(N__24459),
            .sr(N__58203));
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_14_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22581),
            .lcout(\pid_alt.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59331),
            .ce(N__24459),
            .sr(N__58203));
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_17_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22572),
            .lcout(\pid_alt.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59334),
            .ce(N__24461),
            .sr(N__58201));
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_15_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22563),
            .lcout(\pid_alt.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59334),
            .ce(N__24461),
            .sr(N__58201));
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_10_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22554),
            .lcout(\pid_alt.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59334),
            .ce(N__24461),
            .sr(N__58201));
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_19_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22548),
            .lcout(\pid_alt.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59334),
            .ce(N__24461),
            .sr(N__58201));
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_12_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22539),
            .lcout(\pid_alt.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59334),
            .ce(N__24461),
            .sr(N__58201));
    defparam \pid_alt.error_p_reg_esr_8_LC_1_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_8_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22530),
            .lcout(\pid_alt.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59334),
            .ce(N__24461),
            .sr(N__58201));
    defparam \pid_alt.error_p_reg_esr_9_LC_1_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_9_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22524),
            .lcout(\pid_alt.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59334),
            .ce(N__24461),
            .sr(N__58201));
    defparam \pid_alt.error_p_reg_esr_20_LC_1_24_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_24_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_20_LC_1_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22518),
            .lcout(\pid_alt.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59337),
            .ce(N__24462),
            .sr(N__58198));
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_6_LC_2_6_2  (
            .in0(N__58359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55731),
            .lcout(alt_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59154),
            .ce(N__24275),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_6_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_6_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_4_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__53386),
            .in2(_gnd_net_),
            .in3(N__58358),
            .lcout(alt_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59154),
            .ce(N__24275),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_3_LC_2_7_0  (
            .in0(N__58351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55355),
            .lcout(alt_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59169),
            .ce(N__24271),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_7_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_0_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__56465),
            .in2(_gnd_net_),
            .in3(N__58350),
            .lcout(alt_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59169),
            .ce(N__24271),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_2_8_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_2_8_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIQRI31_10_LC_2_8_1  (
            .in0(N__29352),
            .in1(N__31773),
            .in2(_gnd_net_),
            .in3(N__57866),
            .lcout(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_9_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_6_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22942),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59198),
            .ce(N__27615),
            .sr(N__57507));
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_10_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_0_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__56464),
            .in2(_gnd_net_),
            .in3(N__58344),
            .lcout(alt_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59210),
            .ce(N__22616),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_2_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__56125),
            .in2(_gnd_net_),
            .in3(N__58345),
            .lcout(alt_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59210),
            .ce(N__22616),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_2_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_2_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__24627),
            .in2(_gnd_net_),
            .in3(N__24604),
            .lcout(\pid_alt.g0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_3_LC_2_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_3_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_3_LC_2_12_1 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \Commands_frame_decoder.state_3_LC_2_12_1  (
            .in0(N__31741),
            .in1(N__22757),
            .in2(N__22797),
            .in3(N__31317),
            .lcout(\Commands_frame_decoder.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59242),
            .ce(),
            .sr(N__57520));
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_2_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_2_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIFJ1J_3_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__22793),
            .in2(_gnd_net_),
            .in3(N__31739),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_2_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_2_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIEI1J_2_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__25668),
            .in2(_gnd_net_),
            .in3(N__31740),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0 ),
            .ltout(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_2_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_2_12_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIBV7S_2_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22746),
            .in3(N__57854),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_12_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_12_7  (
            .in0(N__24662),
            .in1(N__24625),
            .in2(_gnd_net_),
            .in3(N__24600),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_1_LC_2_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_1_LC_2_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_1_LC_2_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_1_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22722),
            .lcout(\pid_alt.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59259),
            .ce(N__24455),
            .sr(N__58212));
    defparam \pid_alt.error_d_reg_esr_0_LC_2_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_0_LC_2_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_0_LC_2_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_0_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22710),
            .lcout(\pid_alt.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59259),
            .ce(N__24455),
            .sr(N__58212));
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_2_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_2_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_2_14_0  (
            .in0(N__22695),
            .in1(N__22991),
            .in2(N__25157),
            .in3(N__27835),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_14_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_14_1  (
            .in0(N__24351),
            .in1(N__22983),
            .in2(_gnd_net_),
            .in3(N__22973),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_14_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__22992),
            .in2(N__22689),
            .in3(N__27836),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_14_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_14_3  (
            .in0(N__24326),
            .in1(N__22955),
            .in2(_gnd_net_),
            .in3(N__22943),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_5_LC_2_14_4  (
            .in0(N__22974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59274),
            .ce(N__27606),
            .sr(N__57532));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_14_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_14_5  (
            .in0(N__24350),
            .in1(N__22982),
            .in2(_gnd_net_),
            .in3(N__22972),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_7  (
            .in0(N__24327),
            .in1(N__22956),
            .in2(_gnd_net_),
            .in3(N__22944),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_15_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_15_0  (
            .in0(N__22913),
            .in1(N__22884),
            .in2(_gnd_net_),
            .in3(N__22854),
            .lcout(),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_2_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_2_15_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__25727),
            .in2(N__22815),
            .in3(N__23082),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_15_2  (
            .in0(N__25319),
            .in1(N__23224),
            .in2(_gnd_net_),
            .in3(N__24393),
            .lcout(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_2_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_2_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_2_15_3  (
            .in0(N__23194),
            .in1(N__23161),
            .in2(N__23205),
            .in3(N__23127),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_0_LC_2_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_0_LC_2_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_0_LC_2_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_0_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22812),
            .lcout(\pid_alt.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59287),
            .ce(N__24456),
            .sr(N__58210));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_15_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__23223),
            .in2(_gnd_net_),
            .in3(N__24392),
            .lcout(\pid_alt.N_1666_i ),
            .ltout(\pid_alt.N_1666_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_2_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_2_15_7 .LUT_INIT=16'b0100001011010100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_2_15_7  (
            .in0(N__23193),
            .in1(N__23160),
            .in2(N__23130),
            .in3(N__23126),
            .lcout(\pid_alt.un1_pid_prereg_0_axb_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_2_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_2_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_2_16_0  (
            .in0(N__23042),
            .in1(N__23076),
            .in2(N__25400),
            .in3(N__24880),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_2_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_2_16_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_2_16_1  (
            .in0(N__26309),
            .in1(N__26282),
            .in2(_gnd_net_),
            .in3(N__26269),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_2_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_2_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_2_16_2  (
            .in0(N__23043),
            .in1(_gnd_net_),
            .in2(N__23070),
            .in3(N__24881),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_2_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_2_16_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_2_16_3  (
            .in0(N__23063),
            .in1(N__23003),
            .in2(_gnd_net_),
            .in3(N__23033),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_2_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_2_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_2_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_10_LC_2_16_4  (
            .in0(N__26270),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59297),
            .ce(N__27604),
            .sr(N__57546));
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_2_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_2_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_11_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23034),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59297),
            .ce(N__27604),
            .sr(N__57546));
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_11_LC_2_16_7  (
            .in0(N__24882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59297),
            .ce(N__27604),
            .sr(N__57546));
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_2_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_2_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_2_17_0  (
            .in0(N__23297),
            .in1(N__23307),
            .in2(N__25899),
            .in3(N__24829),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_2_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_2_17_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_2_17_1  (
            .in0(N__23255),
            .in1(N__23264),
            .in2(_gnd_net_),
            .in3(N__23287),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_2_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_2_17_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_2_17_2  (
            .in0(N__23298),
            .in1(_gnd_net_),
            .in2(N__23301),
            .in3(N__24830),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_2_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_2_17_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_2_17_3  (
            .in0(N__25542),
            .in1(N__25598),
            .in2(_gnd_net_),
            .in3(N__25565),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_2_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_2_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_2_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_12_LC_2_17_4  (
            .in0(N__23289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59305),
            .ce(N__27602),
            .sr(N__57556));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_2_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_2_17_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_2_17_6  (
            .in0(N__23288),
            .in1(_gnd_net_),
            .in2(N__23268),
            .in3(N__23256),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_2_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_2_17_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_2_17_7  (
            .in0(N__25922),
            .in1(N__25946),
            .in2(N__23238),
            .in3(N__25367),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_18_0  (
            .in0(N__23235),
            .in1(N__23492),
            .in2(N__25458),
            .in3(N__25060),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_18_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_18_1  (
            .in0(N__23484),
            .in1(N__23469),
            .in2(_gnd_net_),
            .in3(N__23459),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_18_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__23493),
            .in2(N__23496),
            .in3(N__25061),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_18_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_18_3  (
            .in0(N__27305),
            .in1(N__27282),
            .in2(_gnd_net_),
            .in3(N__27251),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_18_LC_2_18_4  (
            .in0(N__23460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59311),
            .ce(N__27600),
            .sr(N__57566));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_18_5  (
            .in0(N__23483),
            .in1(N__23468),
            .in2(_gnd_net_),
            .in3(N__23458),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_18_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__28605),
            .in2(N__23439),
            .in3(N__24996),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_LC_2_19_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_2_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_2_19_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_2_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_0_c_RNI1N2F_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(N__32319),
            .in2(_gnd_net_),
            .in3(N__23397),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_19_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__34848),
            .in2(_gnd_net_),
            .in3(N__23355),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_2_19_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_2_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_2_c_RNI5T4F_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__34830),
            .in2(_gnd_net_),
            .in3(N__23310),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_2_19_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_2_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKE1T_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__29658),
            .in2(N__23933),
            .in3(N__23874),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_2_19_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_2_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINI2T_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(N__29643),
            .in2(N__23871),
            .in3(N__23814),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_2_19_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_2_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQM3T_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(N__29628),
            .in2(N__23811),
            .in3(N__23751),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_2_19_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_2_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITQ4T_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(N__29754),
            .in2(N__23748),
            .in3(N__23688),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_2_20_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_2_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI9LEM_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(N__29592),
            .in2(N__23685),
            .in3(N__23625),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_2_20_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_2_20_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_2_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNICPFM_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(N__29607),
            .in2(N__23622),
            .in3(N__23562),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_20_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(N__23964),
            .in2(N__23559),
            .in3(N__23499),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_2_20_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_2_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNI0SDO_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__26199),
            .in2(N__24219),
            .in3(N__24162),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_2_20_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_2_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_11_c_RNI5JAH_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(N__29706),
            .in2(_gnd_net_),
            .in3(N__24114),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_2_20_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_2_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_12_c_RNI7MBH_LC_2_20_5  (
            .in0(_gnd_net_),
            .in1(N__29724),
            .in2(_gnd_net_),
            .in3(N__24066),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_2_20_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_2_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_13_c_RNI9PCH_LC_2_20_6  (
            .in0(_gnd_net_),
            .in1(N__29715),
            .in2(_gnd_net_),
            .in3(N__24027),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_2_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_2_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_2_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_cry_14_c_RNIBSDH_LC_2_20_7  (
            .in0(_gnd_net_),
            .in1(N__29673),
            .in2(_gnd_net_),
            .in3(N__24024),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(N__56312),
            .in2(_gnd_net_),
            .in3(N__58336),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59324),
            .ce(N__27483),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_21_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25488),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_2_22_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_2_22_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_2_22_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_0_LC_2_22_0  (
            .in0(_gnd_net_),
            .in1(N__56487),
            .in2(_gnd_net_),
            .in3(N__58334),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59329),
            .ce(N__27484),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_22_7  (
            .in0(N__58335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55723),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59329),
            .ce(N__27484),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_5_LC_2_23_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_5_LC_2_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_5_LC_2_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_5_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24363),
            .lcout(\pid_alt.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59333),
            .ce(N__24460),
            .sr(N__58200));
    defparam \pid_alt.error_p_reg_esr_6_LC_2_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_6_LC_2_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_6_LC_2_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_6_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24339),
            .lcout(\pid_alt.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59333),
            .ce(N__24460),
            .sr(N__58200));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_24_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_24_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_24_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_24_6  (
            .in0(N__58333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55581),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59336),
            .ce(N__27489),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_7  (
            .in0(_gnd_net_),
            .in1(N__55377),
            .in2(_gnd_net_),
            .in3(N__58332),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59336),
            .ce(N__27489),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_4_LC_3_5_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_4_LC_3_5_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_4_LC_3_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_4_LC_3_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24294),
            .lcout(\pid_alt.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59127),
            .ce(N__24448),
            .sr(N__58216));
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_3_7_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_3_7_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIRSI31_11_LC_3_7_2  (
            .in0(N__27004),
            .in1(N__31772),
            .in2(_gnd_net_),
            .in3(N__57860),
            .lcout(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_7_LC_3_9_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_7_LC_3_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_7_LC_3_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_7_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24255),
            .lcout(\pid_alt.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59182),
            .ce(N__24452),
            .sr(N__58214));
    defparam \pid_alt.error_d_reg_esr_8_LC_3_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_8_LC_3_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_8_LC_3_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_8_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24243),
            .lcout(\pid_alt.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59182),
            .ce(N__24452),
            .sr(N__58214));
    defparam \pid_alt.error_d_reg_esr_9_LC_3_9_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_9_LC_3_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_9_LC_3_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_9_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24231),
            .lcout(\pid_alt.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59182),
            .ce(N__24452),
            .sr(N__58214));
    defparam \pid_alt.error_i_reg_esr_0_LC_3_9_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_0_LC_3_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_0_LC_3_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_0_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24498),
            .lcout(\pid_alt.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59182),
            .ce(N__24452),
            .sr(N__58214));
    defparam \pid_alt.error_i_reg_esr_3_LC_3_9_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_3_LC_3_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_3_LC_3_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_3_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24486),
            .lcout(\pid_alt.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59182),
            .ce(N__24452),
            .sr(N__58214));
    defparam \pid_alt.error_i_reg_esr_11_LC_3_9_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_11_LC_3_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_11_LC_3_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_11_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24474),
            .lcout(\pid_alt.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59182),
            .ce(N__24452),
            .sr(N__58214));
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3  (
            .in0(N__55284),
            .in1(N__56074),
            .in2(_gnd_net_),
            .in3(N__56266),
            .lcout(\Commands_frame_decoder.source_CH1data8lt7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_3_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_3_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_3_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_14_LC_3_11_1  (
            .in0(N__26466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59211),
            .ce(N__27613),
            .sr(N__57511));
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_3_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_3_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_3_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_0_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24391),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59226),
            .ce(N__27610),
            .sr(N__57515));
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_20_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27199),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59226),
            .ce(N__27610),
            .sr(N__57515));
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_3_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_3_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_3_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_3_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24609),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59226),
            .ce(N__27610),
            .sr(N__57515));
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_3_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_3_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_3_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_18_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24995),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59226),
            .ce(N__27610),
            .sr(N__57515));
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_3_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_3_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_3_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_19_LC_3_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25062),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59226),
            .ce(N__27610),
            .sr(N__57515));
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_12_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_13_LC_3_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24831),
            .lcout(\pid_alt.error_i_acumm7lto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59226),
            .ce(N__27610),
            .sr(N__57515));
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_1_LC_3_12_6  (
            .in0(N__25289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59226),
            .ce(N__27610),
            .sr(N__57515));
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_3_13_0  (
            .in0(N__24557),
            .in1(N__24567),
            .in2(N__25242),
            .in3(N__25705),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_3_13_1  (
            .in0(N__24663),
            .in1(N__24626),
            .in2(_gnd_net_),
            .in3(N__24608),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_3_13_2  (
            .in0(N__24558),
            .in1(_gnd_net_),
            .in2(N__24561),
            .in3(N__25706),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_13_3  (
            .in0(N__24548),
            .in1(N__24506),
            .in2(_gnd_net_),
            .in3(N__24523),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_13_4 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_13_4  (
            .in0(N__24524),
            .in1(_gnd_net_),
            .in2(N__24510),
            .in3(N__24549),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_3_13_5  (
            .in0(N__25187),
            .in1(N__24770),
            .in2(N__24528),
            .in3(N__25744),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_3_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_3_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_3_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_4_LC_3_13_6  (
            .in0(N__24525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59243),
            .ce(N__27607),
            .sr(N__57521));
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_13_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_3_13_7  (
            .in0(N__24777),
            .in1(N__24771),
            .in2(_gnd_net_),
            .in3(N__25745),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__25814),
            .in2(N__25647),
            .in3(_gnd_net_),
            .lcout(\pid_alt.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__24762),
            .in2(N__25836),
            .in3(N__24756),
            .lcout(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__25776),
            .in2(N__24753),
            .in3(N__24738),
            .lcout(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__25842),
            .in2(N__24735),
            .in3(N__24723),
            .lcout(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(N__25803),
            .in2(N__24720),
            .in3(N__24702),
            .lcout(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_3_14_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_3_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(N__33366),
            .in2(N__24699),
            .in3(N__24684),
            .lcout(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__26039),
            .in2(N__24681),
            .in3(N__24666),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(N__26024),
            .in2(N__24969),
            .in3(N__24954),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__26009),
            .in2(N__24951),
            .in3(N__24936),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__25997),
            .in2(N__24933),
            .in3(N__24918),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__26066),
            .in2(N__24915),
            .in3(N__24897),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__26051),
            .in2(N__24894),
            .in3(N__24870),
            .lcout(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_3_15_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_3_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__25973),
            .in2(N__24867),
            .in3(N__24852),
            .lcout(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__27960),
            .in2(N__24849),
            .in3(N__24810),
            .lcout(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__24807),
            .in2(_gnd_net_),
            .in3(N__24795),
            .lcout(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24792),
            .in3(N__25134),
            .lcout(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__25131),
            .in2(_gnd_net_),
            .in3(N__25116),
            .lcout(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__25113),
            .in2(_gnd_net_),
            .in3(N__25098),
            .lcout(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__25095),
            .in2(_gnd_net_),
            .in3(N__25080),
            .lcout(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(N__25077),
            .in2(_gnd_net_),
            .in3(N__25035),
            .lcout(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(N__25028),
            .in2(_gnd_net_),
            .in3(N__25032),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5 .C_ON=1'b0;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5  (
            .in0(N__25029),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25011),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_3_16_6  (
            .in0(N__25008),
            .in1(N__28604),
            .in2(N__26562),
            .in3(N__24985),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_16_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_16_7  (
            .in0(N__26232),
            .in1(N__26211),
            .in2(_gnd_net_),
            .in3(N__27647),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_17_0 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__34904),
            .in2(N__34911),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_0_LC_3_17_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_0_LC_3_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_0_LC_3_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_0_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__25335),
            .in2(N__25326),
            .in3(N__25305),
            .lcout(\pid_alt.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .clk(N__59298),
            .ce(N__27601),
            .sr(N__57547));
    defparam \pid_alt.pid_prereg_esr_1_LC_3_17_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_1_LC_3_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_1_LC_3_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_1_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__25302),
            .in2(N__25290),
            .in3(N__25272),
            .lcout(\pid_alt.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .clk(N__59298),
            .ce(N__27601),
            .sr(N__57547));
    defparam \pid_alt.pid_prereg_esr_2_LC_3_17_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_2_LC_3_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_2_LC_3_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_2_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__25269),
            .in2(N__25731),
            .in3(N__25260),
            .lcout(\pid_alt.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .clk(N__59298),
            .ce(N__27601),
            .sr(N__57547));
    defparam \pid_alt.pid_prereg_esr_3_LC_3_17_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_3_LC_3_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_3_LC_3_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_3_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__25257),
            .in2(N__25868),
            .in3(N__25245),
            .lcout(\pid_alt.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .clk(N__59298),
            .ce(N__27601),
            .sr(N__57547));
    defparam \pid_alt.pid_prereg_esr_4_LC_3_17_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_4_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_4_LC_3_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_4_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__25238),
            .in2(N__25218),
            .in3(N__25206),
            .lcout(\pid_alt.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .clk(N__59298),
            .ce(N__27601),
            .sr(N__57547));
    defparam \pid_alt.pid_prereg_esr_5_LC_3_17_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_5_LC_3_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_5_LC_3_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_5_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__25203),
            .in2(N__25194),
            .in3(N__25173),
            .lcout(\pid_alt.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .clk(N__59298),
            .ce(N__27601),
            .sr(N__57547));
    defparam \pid_alt.pid_prereg_esr_6_LC_3_17_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_6_LC_3_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_6_LC_3_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_6_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__25170),
            .in2(N__25158),
            .in3(N__25137),
            .lcout(\pid_alt.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .clk(N__59298),
            .ce(N__27601),
            .sr(N__57547));
    defparam \pid_alt.pid_prereg_esr_7_LC_3_18_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_7_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_7_LC_3_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_7_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__26610),
            .in2(N__26663),
            .in3(N__25422),
            .lcout(\pid_alt.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_8_LC_3_18_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_8_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_8_LC_3_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_8_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__26346),
            .in2(N__26750),
            .in3(N__25419),
            .lcout(\pid_alt.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_9_LC_3_18_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_9_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_9_LC_3_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_9_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__26091),
            .in2(N__26330),
            .in3(N__25416),
            .lcout(\pid_alt.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_10_LC_3_18_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_10_LC_3_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_10_LC_3_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_10_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__26220),
            .in2(N__26187),
            .in3(N__25413),
            .lcout(\pid_alt.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_11_LC_3_18_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_11_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_11_LC_3_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_11_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__25410),
            .in2(N__25401),
            .in3(N__25380),
            .lcout(\pid_alt.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_12_LC_3_18_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_12_LC_3_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_12_LC_3_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_12_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__25377),
            .in2(N__25371),
            .in3(N__25353),
            .lcout(\pid_alt.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_13_LC_3_18_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_13_LC_3_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_13_LC_3_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_13_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__25350),
            .in2(N__25898),
            .in3(N__25344),
            .lcout(\pid_alt.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_14_LC_3_18_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_14_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_14_LC_3_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_14_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__26418),
            .in2(N__26438),
            .in3(N__25341),
            .lcout(\pid_alt.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .clk(N__59306),
            .ce(N__27599),
            .sr(N__57557));
    defparam \pid_alt.pid_prereg_esr_15_LC_3_19_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_15_LC_3_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_15_LC_3_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_15_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__26082),
            .in2(N__26370),
            .in3(N__25338),
            .lcout(\pid_alt.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_16_LC_3_19_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_16_LC_3_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_16_LC_3_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_16_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__26838),
            .in2(N__26889),
            .in3(N__25482),
            .lcout(\pid_alt.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_17_LC_3_19_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_17_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_17_LC_3_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_17_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__26963),
            .in2(N__26604),
            .in3(N__25479),
            .lcout(\pid_alt.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_18_LC_3_19_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_18_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_18_LC_3_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_18_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__25476),
            .in2(N__26561),
            .in3(N__25467),
            .lcout(\pid_alt.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_19_LC_3_19_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_19_LC_3_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_19_LC_3_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_19_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__25464),
            .in2(N__25457),
            .in3(N__25440),
            .lcout(\pid_alt.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_20_LC_3_19_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_20_LC_3_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_20_LC_3_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_20_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__27177),
            .in2(N__27221),
            .in3(N__25437),
            .lcout(\pid_alt.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_21_LC_3_19_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_21_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_21_LC_3_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_21_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__27018),
            .in2(N__27102),
            .in3(N__25434),
            .lcout(\pid_alt.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_22_LC_3_19_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_22_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_22_LC_3_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_22_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__25524),
            .in2(N__25506),
            .in3(N__25431),
            .lcout(\pid_alt.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .clk(N__59312),
            .ce(N__27597),
            .sr(N__57567));
    defparam \pid_alt.pid_prereg_esr_23_LC_3_20_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_23_LC_3_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_23_LC_3_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_23_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__25502),
            .in2(N__25515),
            .in3(N__25428),
            .lcout(\pid_alt.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_23 ),
            .clk(N__59317),
            .ce(N__27595),
            .sr(N__57575));
    defparam \pid_alt.pid_prereg_esr_24_LC_3_20_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_24_LC_3_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_24_LC_3_20_1 .LUT_INIT=16'b1000000101111110;
    LogicCell40 \pid_alt.pid_prereg_esr_24_LC_3_20_1  (
            .in0(N__27086),
            .in1(N__27053),
            .in2(N__27123),
            .in3(N__25425),
            .lcout(\pid_alt.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59317),
            .ce(N__27595),
            .sr(N__57575));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_21_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_21_0  (
            .in0(N__26813),
            .in1(N__26828),
            .in2(_gnd_net_),
            .in3(N__26786),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_3_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_3_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_3_21_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_8_LC_3_21_1  (
            .in0(N__26787),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59320),
            .ce(N__27593),
            .sr(N__57582));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_21_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_21_2  (
            .in0(N__25599),
            .in1(N__25538),
            .in2(_gnd_net_),
            .in3(N__25574),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_3_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_3_21_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_13_LC_3_21_3  (
            .in0(N__25575),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59320),
            .ce(N__27593),
            .sr(N__57582));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_3_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_3_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_3_21_4  (
            .in0(N__27117),
            .in1(N__27081),
            .in2(_gnd_net_),
            .in3(N__27049),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_3_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_3_21_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_3_21_5  (
            .in0(N__27051),
            .in1(_gnd_net_),
            .in2(N__27087),
            .in3(N__27119),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_3_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_3_21_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_3_21_6  (
            .in0(N__27118),
            .in1(N__27082),
            .in2(_gnd_net_),
            .in3(N__27050),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_3_21_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_3_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_3_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_21_LC_3_21_7  (
            .in0(N__27052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59320),
            .ce(N__27593),
            .sr(N__57582));
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_3_22_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_3_22_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_3_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_10_LC_3_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50394),
            .lcout(\dron_frame_decoder_1.drone_altitude_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59325),
            .ce(N__30861),
            .sr(N__57593));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_3_23_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_3_23_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_3_23_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_2_LC_3_23_4  (
            .in0(_gnd_net_),
            .in1(N__56141),
            .in2(_gnd_net_),
            .in3(N__58331),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59330),
            .ce(N__27488),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_23_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_23_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_23_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__55922),
            .in2(_gnd_net_),
            .in3(N__58330),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59330),
            .ce(N__27488),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_11_LC_4_7_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_11_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_11_LC_4_7_7 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \Commands_frame_decoder.state_11_LC_4_7_7  (
            .in0(N__31674),
            .in1(N__29351),
            .in2(N__27012),
            .in3(N__31315),
            .lcout(\Commands_frame_decoder.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59141),
            .ce(),
            .sr(N__57497));
    defparam \Commands_frame_decoder.state_2_LC_4_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_2_LC_4_9_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_2_LC_4_9_2 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \Commands_frame_decoder.state_2_LC_4_9_2  (
            .in0(N__31316),
            .in1(N__31679),
            .in2(N__25667),
            .in3(N__27345),
            .lcout(\Commands_frame_decoder.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59170),
            .ce(),
            .sr(N__57501));
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_4_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_4_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_4_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_15_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38527),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59183),
            .ce(N__27614),
            .sr(N__57503));
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_4_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_4_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_17_LC_4_11_6  (
            .in0(N__28633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59199),
            .ce(N__27611),
            .sr(N__57508));
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_11_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_0_LC_4_11_7  (
            .in0(N__25818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25643),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59199),
            .ce(N__27611),
            .sr(N__57508));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_4_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_4_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_4_12_0  (
            .in0(N__25623),
            .in1(N__25764),
            .in2(N__25617),
            .in3(N__25770),
            .lcout(),
            .ltout(\pid_alt.m7_e_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_4_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_4_12_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_4_12_1  (
            .in0(N__25608),
            .in1(N__25752),
            .in2(N__25602),
            .in3(N__25758),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNIRRP7Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_4_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_16_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26865),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59212),
            .ce(N__27608),
            .sr(N__57512));
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_4_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_4_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_17_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26586),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59212),
            .ce(N__27608),
            .sr(N__57512));
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_4_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_4_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_14_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26391),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59212),
            .ce(N__27608),
            .sr(N__57512));
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_4_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_4_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_4_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_15_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26529),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_4_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_4_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_12_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25923),
            .lcout(\pid_alt.error_i_acumm7lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_5_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25746),
            .lcout(\pid_alt.error_i_acumm7lto5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_9_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26169),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_4_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_4_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_7_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26624),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_4_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_4_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_2_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25726),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_4_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_4_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_4_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25707),
            .lcout(\pid_alt.error_i_acumm7lto4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_4_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_4_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_3_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25861),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59227),
            .ce(N__27605),
            .sr(N__57516));
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_14_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_3_LC_4_14_0  (
            .in0(N__33388),
            .in1(N__27900),
            .in2(N__25797),
            .in3(N__27378),
            .lcout(\pid_alt.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59244),
            .ce(N__27951),
            .sr(N__33338));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_14_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_14_1  (
            .in0(N__27394),
            .in1(_gnd_net_),
            .in2(N__33428),
            .in3(N__33385),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNIEPGB3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_14_2 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_1_LC_4_14_2  (
            .in0(N__33386),
            .in1(N__27720),
            .in2(N__25796),
            .in3(N__27904),
            .lcout(\pid_alt.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59244),
            .ce(N__27951),
            .sr(N__33338));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_14_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_14_3  (
            .in0(N__28039),
            .in1(N__28006),
            .in2(_gnd_net_),
            .in3(N__27983),
            .lcout(\pid_alt.N_9_0 ),
            .ltout(\pid_alt.N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_14_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_14_4  (
            .in0(N__27873),
            .in1(N__25986),
            .in2(N__25824),
            .in3(N__27393),
            .lcout(\pid_alt.N_62_mux ),
            .ltout(\pid_alt.N_62_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_14_5 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_0_LC_4_14_5  (
            .in0(N__27702),
            .in1(N__27896),
            .in2(N__25821),
            .in3(N__25788),
            .lcout(\pid_alt.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59244),
            .ce(N__27951),
            .sr(N__33338));
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_14_6 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \pid_alt.error_i_acumm_esr_4_LC_4_14_6  (
            .in0(N__33389),
            .in1(N__33424),
            .in2(N__27905),
            .in3(N__27395),
            .lcout(\pid_alt.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59244),
            .ce(N__27951),
            .sr(N__33338));
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_14_7 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \pid_alt.error_i_acumm_esr_2_LC_4_14_7  (
            .in0(N__27366),
            .in1(N__25792),
            .in2(N__27906),
            .in3(N__33387),
            .lcout(\pid_alt.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59244),
            .ce(N__27951),
            .sr(N__33338));
    defparam \pid_alt.error_i_acumm_10_LC_4_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_10_LC_4_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_10_LC_4_15_0 .LUT_INIT=16'b1101100011111010;
    LogicCell40 \pid_alt.error_i_acumm_10_LC_4_15_0  (
            .in0(N__39731),
            .in1(N__27630),
            .in2(N__26070),
            .in3(N__27409),
            .lcout(\pid_alt.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59260),
            .ce(),
            .sr(N__33331));
    defparam \pid_alt.error_i_acumm_11_LC_4_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_11_LC_4_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_11_LC_4_15_1 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \pid_alt.error_i_acumm_11_LC_4_15_1  (
            .in0(N__27410),
            .in1(N__27766),
            .in2(N__26055),
            .in3(N__39735),
            .lcout(\pid_alt.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59260),
            .ce(),
            .sr(N__33331));
    defparam \pid_alt.error_i_acumm_6_LC_4_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_6_LC_4_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_6_LC_4_15_2 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \pid_alt.error_i_acumm_6_LC_4_15_2  (
            .in0(N__26040),
            .in1(N__27735),
            .in2(N__39738),
            .in3(N__27411),
            .lcout(\pid_alt.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59260),
            .ce(),
            .sr(N__33331));
    defparam \pid_alt.error_i_acumm_7_LC_4_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_7_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_7_LC_4_15_3 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \pid_alt.error_i_acumm_7_LC_4_15_3  (
            .in0(N__27412),
            .in1(N__27933),
            .in2(N__26028),
            .in3(N__39736),
            .lcout(\pid_alt.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59260),
            .ce(),
            .sr(N__33331));
    defparam \pid_alt.error_i_acumm_8_LC_4_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_8_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_8_LC_4_15_4 .LUT_INIT=16'b1011100011111100;
    LogicCell40 \pid_alt.error_i_acumm_8_LC_4_15_4  (
            .in0(N__27783),
            .in1(N__39730),
            .in2(N__26013),
            .in3(N__27413),
            .lcout(\pid_alt.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59260),
            .ce(),
            .sr(N__33331));
    defparam \pid_alt.error_i_acumm_9_LC_4_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_9_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_9_LC_4_15_5 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \pid_alt.error_i_acumm_9_LC_4_15_5  (
            .in0(N__27414),
            .in1(N__25998),
            .in2(N__27801),
            .in3(N__39737),
            .lcout(\pid_alt.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59260),
            .ce(),
            .sr(N__33331));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(N__27932),
            .in2(_gnd_net_),
            .in3(N__27734),
            .lcout(\pid_alt.m35_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_12_LC_4_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_12_LC_4_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_12_LC_4_15_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \pid_alt.error_i_acumm_12_LC_4_15_7  (
            .in0(N__39729),
            .in1(N__27681),
            .in2(N__25977),
            .in3(N__28077),
            .lcout(\pid_alt.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59260),
            .ce(),
            .sr(N__33331));
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_4_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_4_16_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_4_16_0  (
            .in0(N__25962),
            .in1(N__25950),
            .in2(_gnd_net_),
            .in3(N__25918),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_4_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_4_16_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_4_16_1  (
            .in0(N__26313),
            .in1(N__26286),
            .in2(_gnd_net_),
            .in3(N__26271),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_4_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_4_16_2  (
            .in0(N__26183),
            .in1(N__26210),
            .in2(N__26223),
            .in3(N__27646),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_3  (
            .in0(N__26132),
            .in1(N__26144),
            .in2(_gnd_net_),
            .in3(N__26167),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_4_16_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_4_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29445),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_16_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_4_16_5  (
            .in0(N__26109),
            .in1(N__26115),
            .in2(_gnd_net_),
            .in3(N__27815),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_6  (
            .in0(N__26168),
            .in1(_gnd_net_),
            .in2(N__26148),
            .in3(N__26133),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_16_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_4_16_7  (
            .in0(N__26108),
            .in1(N__26331),
            .in2(N__26094),
            .in3(N__27814),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_17_0  (
            .in0(N__26507),
            .in1(N__26538),
            .in2(N__26366),
            .in3(N__26524),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_17_1 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_17_1  (
            .in0(N__26481),
            .in1(N__26499),
            .in2(_gnd_net_),
            .in3(N__26462),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_17_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_17_2  (
            .in0(N__26508),
            .in1(_gnd_net_),
            .in2(N__26532),
            .in3(N__26525),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_17_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_17_3  (
            .in0(N__38486),
            .in1(N__38453),
            .in2(_gnd_net_),
            .in3(N__38529),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_17_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_17_4  (
            .in0(N__26498),
            .in1(N__26480),
            .in2(_gnd_net_),
            .in3(N__26461),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_17_5  (
            .in0(N__26439),
            .in1(N__26405),
            .in2(N__26421),
            .in3(N__26386),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_17_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_17_7  (
            .in0(N__26412),
            .in1(N__26406),
            .in2(_gnd_net_),
            .in3(N__26387),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_4_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_4_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_4_18_0  (
            .in0(N__26759),
            .in1(N__26340),
            .in2(N__26751),
            .in3(N__27865),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_4_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_4_18_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_4_18_1  (
            .in0(N__26699),
            .in1(N__26708),
            .in2(_gnd_net_),
            .in3(N__26731),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_4_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_4_18_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_4_18_2  (
            .in0(N__26760),
            .in1(_gnd_net_),
            .in2(N__26334),
            .in3(N__27866),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_4_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_4_18_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_4_18_3  (
            .in0(N__26829),
            .in1(N__26814),
            .in2(_gnd_net_),
            .in3(N__26780),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_4_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_4_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_4_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_7_LC_4_18_4  (
            .in0(N__26733),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59299),
            .ce(N__27598),
            .sr(N__57548));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_4_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_4_18_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_4_18_5  (
            .in0(N__26679),
            .in1(N__26685),
            .in2(_gnd_net_),
            .in3(N__26631),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_18_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_18_6  (
            .in0(N__26732),
            .in1(_gnd_net_),
            .in2(N__26712),
            .in3(N__26700),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_4_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_4_18_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_4_18_7  (
            .in0(N__26678),
            .in1(N__26664),
            .in2(N__26634),
            .in3(N__26630),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_4_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_4_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_4_19_0  (
            .in0(N__26595),
            .in1(N__26975),
            .in2(N__26967),
            .in3(N__26584),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_4_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_4_19_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_4_19_1  (
            .in0(N__28661),
            .in1(N__28685),
            .in2(_gnd_net_),
            .in3(N__28640),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_4_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_4_19_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(N__26976),
            .in2(N__26589),
            .in3(N__26585),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_19_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_19_3  (
            .in0(N__26912),
            .in1(N__26921),
            .in2(_gnd_net_),
            .in3(N__26950),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_4_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_4_19_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_16_LC_4_19_4  (
            .in0(N__26952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59307),
            .ce(N__27596),
            .sr(N__57558));
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_4_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_4_19_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_4_19_5  (
            .in0(N__26895),
            .in1(N__38430),
            .in2(_gnd_net_),
            .in3(N__26864),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_4_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_4_19_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_4_19_6  (
            .in0(N__26951),
            .in1(_gnd_net_),
            .in2(N__26925),
            .in3(N__26913),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_4_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_4_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_4_19_7  (
            .in0(N__26888),
            .in1(N__38429),
            .in2(N__26868),
            .in3(N__26863),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_4_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_4_20_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_4_20_0  (
            .in0(N__27170),
            .in1(N__27155),
            .in2(_gnd_net_),
            .in3(N__27145),
            .lcout(\pid_alt.un1_pid_prereg_236_1 ),
            .ltout(\pid_alt.un1_pid_prereg_236_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_4_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_4_20_1 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__27231),
            .in2(N__26832),
            .in3(N__27201),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_4_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_4_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_4_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_20_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27147),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59313),
            .ce(N__27594),
            .sr(N__57568));
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_4_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_4_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_19_LC_4_20_3  (
            .in0(N__27261),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59313),
            .ce(N__27594),
            .sr(N__57568));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_4_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_4_20_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_4_20_4  (
            .in0(N__27306),
            .in1(N__27275),
            .in2(_gnd_net_),
            .in3(N__27260),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_4_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_4_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_4_20_5  (
            .in0(N__27225),
            .in1(N__27079),
            .in2(N__27204),
            .in3(N__27200),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_4_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_4_20_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_4_20_6  (
            .in0(N__27171),
            .in1(N__27156),
            .in2(_gnd_net_),
            .in3(N__27146),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_4_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_4_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_4_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_4_20_7  (
            .in0(N__27101),
            .in1(N__27080),
            .in2(N__27057),
            .in3(N__27054),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_12_LC_5_7_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_12_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_12_LC_5_7_0 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \Commands_frame_decoder.state_12_LC_5_7_0  (
            .in0(N__27011),
            .in1(N__26987),
            .in2(N__31738),
            .in3(N__31290),
            .lcout(\Commands_frame_decoder.stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59128),
            .ce(),
            .sr(N__57496));
    defparam \Commands_frame_decoder.state_13_LC_5_7_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_13_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_13_LC_5_7_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \Commands_frame_decoder.state_13_LC_5_7_7  (
            .in0(N__31291),
            .in1(N__31804),
            .in2(N__26988),
            .in3(N__31678),
            .lcout(\Commands_frame_decoder.stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59128),
            .ce(),
            .sr(N__57496));
    defparam \uart_pc.data_rdy_LC_5_8_1 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_5_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.data_rdy_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__30344),
            .in2(_gnd_net_),
            .in3(N__29292),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59142),
            .ce(),
            .sr(N__57498));
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_5_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_5_9_0 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_0_LC_5_9_0  (
            .in0(N__27332),
            .in1(N__27539),
            .in2(N__29067),
            .in3(N__27507),
            .lcout(\Commands_frame_decoder.N_377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_5_9_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_5_9_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_5_9_1  (
            .in0(N__53325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56224),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_5_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_5_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_0_LC_5_9_2  (
            .in0(N__55705),
            .in1(N__31655),
            .in2(N__27351),
            .in3(N__55332),
            .lcout(\Commands_frame_decoder.N_416 ),
            .ltout(\Commands_frame_decoder.N_416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_5_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_5_9_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_2_LC_5_9_3  (
            .in0(N__27339),
            .in1(N__55846),
            .in2(N__27348),
            .in3(N__56046),
            .lcout(\Commands_frame_decoder.N_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_5_9_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_5_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNI6QPK_1_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__31831),
            .in2(_gnd_net_),
            .in3(N__27523),
            .lcout(\Commands_frame_decoder.N_376_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_5_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_5_9_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_2_LC_5_9_6  (
            .in0(N__56433),
            .in1(N__27522),
            .in2(_gnd_net_),
            .in3(N__55521),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_0_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_5_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_5_10_1 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_0_LC_5_10_1  (
            .in0(N__31304),
            .in1(N__31726),
            .in2(N__29198),
            .in3(N__27333),
            .lcout(),
            .ltout(\Commands_frame_decoder.N_376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_0_LC_5_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_0_LC_5_10_2 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_0_LC_5_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.state_0_LC_5_10_2  (
            .in0(N__29268),
            .in1(N__27321),
            .in2(N__27315),
            .in3(N__27312),
            .lcout(\Commands_frame_decoder.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59171),
            .ce(),
            .sr(N__57502));
    defparam \Commands_frame_decoder.state_14_LC_5_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_14_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_14_LC_5_10_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_14_LC_5_10_3  (
            .in0(N__31808),
            .in1(N__29267),
            .in2(_gnd_net_),
            .in3(N__31727),
            .lcout(\Commands_frame_decoder.stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59171),
            .ce(),
            .sr(N__57502));
    defparam \Commands_frame_decoder.state_RNIOMNA5_1_LC_5_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIOMNA5_1_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIOMNA5_1_LC_5_10_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Commands_frame_decoder.state_RNIOMNA5_1_LC_5_10_4  (
            .in0(N__31725),
            .in1(N__27525),
            .in2(_gnd_net_),
            .in3(N__31303),
            .lcout(\Commands_frame_decoder.N_379 ),
            .ltout(\Commands_frame_decoder.N_379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_LC_5_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_LC_5_10_5 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \Commands_frame_decoder.state_1_LC_5_10_5  (
            .in0(N__29178),
            .in1(N__27540),
            .in2(N__27528),
            .in3(N__55549),
            .lcout(\Commands_frame_decoder.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59171),
            .ce(),
            .sr(N__57502));
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_5_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_5_10_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_2_0_LC_5_10_7  (
            .in0(N__27524),
            .in1(N__56440),
            .in2(N__56106),
            .in3(N__29159),
            .lcout(\Commands_frame_decoder.N_412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_9_LC_5_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_9_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_9_LC_5_11_0 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \Commands_frame_decoder.state_9_LC_5_11_0  (
            .in0(N__31314),
            .in1(N__27497),
            .in2(N__31774),
            .in3(N__27426),
            .lcout(\Commands_frame_decoder.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59184),
            .ce(),
            .sr(N__57504));
    defparam \Commands_frame_decoder.state_8_LC_5_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_8_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_8_LC_5_11_7 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \Commands_frame_decoder.state_8_LC_5_11_7  (
            .in0(N__29391),
            .in1(N__31728),
            .in2(N__27501),
            .in3(N__31313),
            .lcout(\Commands_frame_decoder.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59184),
            .ce(),
            .sr(N__57504));
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_5_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_5_12_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIF38S_6_LC_5_12_0  (
            .in0(N__29550),
            .in1(N__31778),
            .in2(_gnd_net_),
            .in3(N__57837),
            .lcout(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_12_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_12_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_5_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_5_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNILP1J_9_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__27425),
            .in2(_gnd_net_),
            .in3(N__31777),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_5_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_5_13_5 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_5_13_5  (
            .in0(N__28013),
            .in1(N__27677),
            .in2(N__28059),
            .in3(N__27979),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNI175BZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_5_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_5_13_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__27377),
            .in2(_gnd_net_),
            .in3(N__27362),
            .lcout(),
            .ltout(\pid_alt.m21_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_5_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_5_13_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_5_13_7  (
            .in0(N__27925),
            .in1(N__33420),
            .in2(N__27909),
            .in3(N__27895),
            .lcout(\pid_alt.m21_e_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_5_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_5_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_5_14_0  (
            .in0(N__27797),
            .in1(N__27782),
            .in2(N__27768),
            .in3(N__27629),
            .lcout(\pid_alt.m35_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_5_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_8_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27867),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59228),
            .ce(N__27603),
            .sr(N__57517));
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_5_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_6_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27840),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59228),
            .ce(N__27603),
            .sr(N__57517));
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_5_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_9_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27822),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59228),
            .ce(N__27603),
            .sr(N__57517));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_5_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_5_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_5_14_4  (
            .in0(N__27796),
            .in1(N__27781),
            .in2(N__27767),
            .in3(N__27733),
            .lcout(),
            .ltout(\pid_alt.m21_e_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEK7C2_0_LC_5_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEK7C2_0_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEK7C2_0_LC_5_14_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIEK7C2_0_LC_5_14_5  (
            .in0(N__27719),
            .in1(N__27701),
            .in2(N__27684),
            .in3(N__27660),
            .lcout(\pid_alt.m21_e_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_5_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_5_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__27628),
            .in2(_gnd_net_),
            .in3(N__27676),
            .lcout(\pid_alt.m21_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_5_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_5_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_10_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27654),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59228),
            .ce(N__27603),
            .sr(N__57517));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_5_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_5_15_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_5_15_1  (
            .in0(N__28092),
            .in1(N__28083),
            .in2(N__28058),
            .in3(N__28076),
            .lcout(),
            .ltout(\pid_alt.error_i_acumm_prereg_esr_RNIO7B05Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIAAPN5_1_LC_5_15_2 .C_ON=1'b0;
    defparam \pid_alt.state_RNIAAPN5_1_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIAAPN5_1_LC_5_15_2 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \pid_alt.state_RNIAAPN5_1_LC_5_15_2  (
            .in0(N__39720),
            .in1(_gnd_net_),
            .in2(N__28065),
            .in3(N__44979),
            .lcout(\pid_alt.un1_reset_1_0_i ),
            .ltout(\pid_alt.un1_reset_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIVV066_1_LC_5_15_3 .C_ON=1'b0;
    defparam \pid_alt.state_RNIVV066_1_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIVV066_1_LC_5_15_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_alt.state_RNIVV066_1_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28062),
            .in3(N__39721),
            .lcout(\pid_alt.N_72_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_13_LC_5_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_13_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_13_LC_5_15_5 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \pid_alt.error_i_acumm_esr_13_LC_5_15_5  (
            .in0(N__28054),
            .in1(N__28014),
            .in2(_gnd_net_),
            .in3(N__27987),
            .lcout(\pid_alt.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59245),
            .ce(N__27950),
            .sr(N__33330));
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_15_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_15_6 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_5_15_6  (
            .in0(N__39719),
            .in1(N__44978),
            .in2(N__28910),
            .in3(N__28545),
            .lcout(),
            .ltout(\pid_alt.un1_reset_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_15_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_15_7 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_5_15_7  (
            .in0(N__28320),
            .in1(N__28960),
            .in2(N__27939),
            .in3(N__28832),
            .lcout(\pid_alt.un1_reset_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_16_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_16_0 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_16_0  (
            .in0(N__28961),
            .in1(N__28899),
            .in2(N__28779),
            .in3(N__28833),
            .lcout(\pid_alt.source_pid_9_0_tz_6 ),
            .ltout(\pid_alt.source_pid_9_0_tz_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_10_LC_5_16_1 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_10_LC_5_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_10_LC_5_16_1 .LUT_INIT=16'b1110111001001110;
    LogicCell40 \pid_alt.source_pid_1_10_LC_5_16_1  (
            .in0(N__39723),
            .in1(N__34717),
            .in2(N__27936),
            .in3(N__28257),
            .lcout(throttle_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59261),
            .ce(),
            .sr(N__28708));
    defparam \pid_alt.source_pid_1_11_LC_5_16_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_11_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_11_LC_5_16_2 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_11_LC_5_16_2  (
            .in0(N__28148),
            .in1(N__39726),
            .in2(N__40045),
            .in3(N__28305),
            .lcout(throttle_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59261),
            .ce(),
            .sr(N__28708));
    defparam \pid_alt.source_pid_1_6_LC_5_16_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_6_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_6_LC_5_16_3 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_6_LC_5_16_3  (
            .in0(N__39724),
            .in1(N__28149),
            .in2(N__36124),
            .in3(N__28179),
            .lcout(throttle_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59261),
            .ce(),
            .sr(N__28708));
    defparam \pid_alt.source_pid_1_7_LC_5_16_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_7_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_7_LC_5_16_4 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_7_LC_5_16_4  (
            .in0(N__28150),
            .in1(N__39727),
            .in2(N__36215),
            .in3(N__28206),
            .lcout(throttle_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59261),
            .ce(),
            .sr(N__28708));
    defparam \pid_alt.source_pid_1_8_LC_5_16_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_8_LC_5_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_8_LC_5_16_5 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_8_LC_5_16_5  (
            .in0(N__39725),
            .in1(N__28151),
            .in2(N__35971),
            .in3(N__28230),
            .lcout(throttle_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59261),
            .ce(),
            .sr(N__28708));
    defparam \pid_alt.source_pid_1_9_LC_5_16_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_9_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_9_LC_5_16_6 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_9_LC_5_16_6  (
            .in0(N__28152),
            .in1(N__39728),
            .in2(N__36058),
            .in3(N__28281),
            .lcout(throttle_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59261),
            .ce(),
            .sr(N__28708));
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_16_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_16_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_alt.state_RNIOVDUE_1_LC_5_16_7  (
            .in0(N__39722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28699),
            .lcout(\pid_alt.N_72_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_17_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_17_0  (
            .in0(N__28103),
            .in1(N__28130),
            .in2(N__28119),
            .in3(N__28337),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_2_LC_5_17_1 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_2_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_2_LC_5_17_1 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \pid_alt.source_pid_1_esr_2_LC_5_17_1  (
            .in0(N__28835),
            .in1(N__28349),
            .in2(N__28134),
            .in3(N__28901),
            .lcout(throttle_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59275),
            .ce(N__28730),
            .sr(N__28715));
    defparam \pid_alt.source_pid_1_esr_3_LC_5_17_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_3_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_3_LC_5_17_2 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \pid_alt.source_pid_1_esr_3_LC_5_17_2  (
            .in0(N__28118),
            .in1(N__28906),
            .in2(N__28353),
            .in3(N__28837),
            .lcout(throttle_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59275),
            .ce(N__28730),
            .sr(N__28715));
    defparam \pid_alt.source_pid_1_esr_1_LC_5_17_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_1_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_1_LC_5_17_3 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_1_LC_5_17_3  (
            .in0(N__28834),
            .in1(N__28348),
            .in2(N__28911),
            .in3(N__28104),
            .lcout(throttle_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59275),
            .ce(N__28730),
            .sr(N__28715));
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_17_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_17_4 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_17_4  (
            .in0(N__28959),
            .in1(N__28774),
            .in2(_gnd_net_),
            .in3(N__28557),
            .lcout(\pid_alt.N_44 ),
            .ltout(\pid_alt.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_17_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_17_5 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_17_5  (
            .in0(N__28415),
            .in1(_gnd_net_),
            .in2(N__28356),
            .in3(N__28388),
            .lcout(\pid_alt.N_46 ),
            .ltout(\pid_alt.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_0_LC_5_17_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_0_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_0_LC_5_17_6 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \pid_alt.source_pid_1_esr_0_LC_5_17_6  (
            .in0(N__28900),
            .in1(N__28338),
            .in2(N__28326),
            .in3(N__28836),
            .lcout(throttle_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59275),
            .ce(N__28730),
            .sr(N__28715));
    defparam \pid_front.error_d_reg_esr_RNI1VUF_9_LC_5_17_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNI1VUF_9_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNI1VUF_9_LC_5_17_7 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \pid_front.error_d_reg_esr_RNI1VUF_9_LC_5_17_7  (
            .in0(N__30774),
            .in1(N__32304),
            .in2(N__56775),
            .in3(N__32271),
            .lcout(\pid_front.error_d_reg_esr_RNI1VUFZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_18_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_18_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_18_0  (
            .in0(N__28252),
            .in1(N__28311),
            .in2(N__28205),
            .in3(N__39678),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_18_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_18_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_18_1  (
            .in0(N__28390),
            .in1(N__28569),
            .in2(N__28323),
            .in3(N__28414),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_5_18_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_5_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_5_18_2  (
            .in0(N__28226),
            .in1(N__28178),
            .in2(N__28280),
            .in3(N__28301),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI8H141_10_LC_5_18_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI8H141_10_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI8H141_10_LC_5_18_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI8H141_10_LC_5_18_3  (
            .in0(N__28300),
            .in1(N__28273),
            .in2(N__28256),
            .in3(N__28225),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_5_18_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_5_18_4 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_5_18_4  (
            .in0(N__28198),
            .in1(_gnd_net_),
            .in2(N__28182),
            .in3(N__28177),
            .lcout(\pid_alt.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_18_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_18_5 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_18_5  (
            .in0(N__28764),
            .in1(N__28991),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.N_90 ),
            .ltout(\pid_alt.N_90_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_18_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_18_6  (
            .in0(N__39677),
            .in1(N__28389),
            .in2(N__28572),
            .in3(N__28941),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_18_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_18_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_18_7  (
            .in0(N__28808),
            .in1(N__28568),
            .in2(N__28560),
            .in3(N__28556),
            .lcout(\pid_alt.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_19_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_19_0  (
            .in0(N__28536),
            .in1(N__28527),
            .in2(N__28515),
            .in3(N__28500),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_19_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_19_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_19_1  (
            .in0(N__28491),
            .in1(N__28479),
            .in2(N__28470),
            .in3(N__28458),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_19_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_19_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_5_19_2  (
            .in0(N__28449),
            .in1(N__28443),
            .in2(N__28431),
            .in3(N__28428),
            .lcout(\pid_alt.N_305 ),
            .ltout(\pid_alt.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_19_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_19_3 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_19_3  (
            .in0(N__28391),
            .in1(N__28419),
            .in2(N__28398),
            .in3(N__28902),
            .lcout(),
            .ltout(\pid_alt.source_pid_9_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_4_LC_5_19_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_4_LC_5_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_4_LC_5_19_4 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \pid_alt.source_pid_1_esr_4_LC_5_19_4  (
            .in0(N__29004),
            .in1(N__28825),
            .in2(N__28395),
            .in3(N__28392),
            .lcout(throttle_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59300),
            .ce(N__28731),
            .sr(N__28716));
    defparam \pid_alt.source_pid_1_esr_5_LC_5_19_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_5_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_5_LC_5_19_5 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_5_LC_5_19_5  (
            .in0(N__28905),
            .in1(N__29003),
            .in2(N__28839),
            .in3(N__28992),
            .lcout(throttle_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59300),
            .ce(N__28731),
            .sr(N__28716));
    defparam \pid_alt.source_pid_1_esr_13_LC_5_19_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_13_LC_5_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_13_LC_5_19_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.source_pid_1_esr_13_LC_5_19_6  (
            .in0(N__28904),
            .in1(N__28824),
            .in2(_gnd_net_),
            .in3(N__28967),
            .lcout(throttle_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59300),
            .ce(N__28731),
            .sr(N__28716));
    defparam \pid_alt.source_pid_1_esr_12_LC_5_19_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_12_LC_5_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_12_LC_5_19_7 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_12_LC_5_19_7  (
            .in0(N__28968),
            .in1(N__28903),
            .in2(N__28838),
            .in3(N__28778),
            .lcout(throttle_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59300),
            .ce(N__28731),
            .sr(N__28716));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_5_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_5_20_0 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_5_20_0  (
            .in0(N__28686),
            .in1(N__28665),
            .in2(_gnd_net_),
            .in3(N__28644),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state57_i_LC_7_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state57_i_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state57_i_LC_7_6_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.un1_state57_i_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__31771),
            .in2(_gnd_net_),
            .in3(N__57851),
            .lcout(\Commands_frame_decoder.un1_state57_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_7_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_7_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_7_7_0  (
            .in0(N__29085),
            .in1(N__29036),
            .in2(N__29088),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_7_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__29136),
            .in2(_gnd_net_),
            .in3(N__28581),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_7_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__29881),
            .in2(_gnd_net_),
            .in3(N__28578),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_7_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__29919),
            .in2(_gnd_net_),
            .in3(N__28575),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_7_7_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_7_7_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_7_7_4  (
            .in0(N__29086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29037),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_7_7_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_7_7_5 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_4_LC_7_7_5  (
            .in0(N__57881),
            .in1(N__29992),
            .in2(N__29118),
            .in3(N__29049),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59108),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_7_7_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_7_7_6 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_pc.timer_Count_1_LC_7_7_6  (
            .in0(N__29043),
            .in1(N__29110),
            .in2(N__29998),
            .in3(N__57882),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59108),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_7_7_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_7_7_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_3_LC_7_7_7  (
            .in0(N__57880),
            .in1(N__29991),
            .in2(N__29117),
            .in3(N__29028),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59108),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_8_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_8_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_7_8_0  (
            .in0(N__30620),
            .in1(N__29930),
            .in2(_gnd_net_),
            .in3(N__29878),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(\uart_pc.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_4_LC_7_8_1 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_7_8_1 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \uart_pc.state_4_LC_7_8_1  (
            .in0(N__30237),
            .in1(N__29108),
            .in2(N__29022),
            .in3(N__44951),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59116),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_8_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_8_2 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_7_8_2  (
            .in0(N__29967),
            .in1(N__30029),
            .in2(N__29019),
            .in3(N__30236),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3  (
            .in0(N__29876),
            .in1(N__29134),
            .in2(N__29937),
            .in3(N__29965),
            .lcout(\uart_pc.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_7_8_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_7_8_4 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.timer_Count_2_LC_7_8_4  (
            .in0(N__29109),
            .in1(N__29010),
            .in2(N__30003),
            .in3(N__57869),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59116),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_8_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_7_8_5  (
            .in0(N__29877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29135),
            .lcout(\uart_pc.N_126_li ),
            .ltout(\uart_pc.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_8_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_8_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_7_8_6  (
            .in0(N__29966),
            .in1(N__29931),
            .in2(N__29121),
            .in3(N__57867),
            .lcout(\uart_pc.N_143 ),
            .ltout(\uart_pc.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_7_8_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_7_8_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_pc.timer_Count_0_LC_7_8_7  (
            .in0(N__57868),
            .in1(N__29999),
            .in2(N__29091),
            .in3(N__29087),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59116),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_4_LC_7_9_0 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_7_9_0 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \uart_pc.data_1_4_LC_7_9_0  (
            .in0(N__29251),
            .in1(N__30411),
            .in2(N__29228),
            .in3(N__55818),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59129),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_7_9_1 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_7_9_1 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \uart_pc.data_0_LC_7_9_1  (
            .in0(N__56388),
            .in1(N__29218),
            .in2(N__30108),
            .in3(N__29250),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59129),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_7_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_7_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_3_0_LC_7_9_2  (
            .in0(N__56001),
            .in1(N__55446),
            .in2(N__56441),
            .in3(N__55817),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_7_9_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_7_9_3 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_7_9_3  (
            .in0(N__29287),
            .in1(N__30326),
            .in2(_gnd_net_),
            .in3(N__57861),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_7_9_4 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_7_9_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \uart_pc.data_4_LC_7_9_4  (
            .in0(N__30422),
            .in1(N__29288),
            .in2(N__29052),
            .in3(N__53324),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59129),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_2_LC_7_9_5 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_7_9_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \uart_pc.data_2_LC_7_9_5  (
            .in0(N__30074),
            .in1(N__29222),
            .in2(N__56073),
            .in3(N__29253),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59129),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__29286),
            .in2(_gnd_net_),
            .in3(N__44970),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_7_9_7 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_7_9_7 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \uart_pc.data_1_LC_7_9_7  (
            .in0(N__30089),
            .in1(N__29252),
            .in2(N__29271),
            .in3(N__56220),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59129),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNISEFT5_0_LC_7_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNISEFT5_0_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNISEFT5_0_LC_7_10_0 .LUT_INIT=16'b0000100001001100;
    LogicCell40 \Commands_frame_decoder.count_RNISEFT5_0_LC_7_10_0  (
            .in0(N__31763),
            .in1(N__31840),
            .in2(N__31866),
            .in3(N__31269),
            .lcout(\Commands_frame_decoder.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_5_LC_7_10_1 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_7_10_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \uart_pc.data_5_LC_7_10_1  (
            .in0(N__29255),
            .in1(N__30392),
            .in2(N__29229),
            .in3(N__55666),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59143),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_3_LC_7_10_2 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_7_10_2 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \uart_pc.data_3_LC_7_10_2  (
            .in0(N__55280),
            .in1(N__29223),
            .in2(N__30060),
            .in3(N__29254),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59143),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_6_LC_7_10_4 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_7_10_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \uart_pc.data_6_LC_7_10_4  (
            .in0(N__30278),
            .in1(N__29256),
            .in2(N__55534),
            .in3(N__29227),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59143),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_7_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_7_10_5 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \Commands_frame_decoder.count_0_LC_7_10_5  (
            .in0(N__31841),
            .in1(N__31864),
            .in2(N__31785),
            .in3(N__57853),
            .lcout(\Commands_frame_decoder.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59143),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_10_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_1_LC_7_10_6  (
            .in0(N__56384),
            .in1(N__56016),
            .in2(N__29199),
            .in3(N__55835),
            .lcout(\Commands_frame_decoder.state_ns_0_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIEAGS_4_LC_7_10_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_7_10_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_7_10_7  (
            .in0(N__30249),
            .in1(N__29973),
            .in2(_gnd_net_),
            .in3(N__57852),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_7_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_7_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__55445),
            .in2(_gnd_net_),
            .in3(N__55845),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_7_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_7_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIHL1J_5_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__29574),
            .in2(_gnd_net_),
            .in3(N__31762),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_7_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_7_11_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIE28S_5_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29436),
            .in3(N__57864),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0  (
            .in0(N__29410),
            .in1(N__31767),
            .in2(N__29387),
            .in3(N__53349),
            .lcout(xy_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59172),
            .ce(),
            .sr(N__57509));
    defparam \Commands_frame_decoder.state_7_LC_7_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_7_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_7_LC_7_12_1 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \Commands_frame_decoder.state_7_LC_7_12_1  (
            .in0(N__31766),
            .in1(N__29383),
            .in2(N__29549),
            .in3(N__31306),
            .lcout(\Commands_frame_decoder.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59172),
            .ce(),
            .sr(N__57509));
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_7_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_7_12_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIG48S_7_LC_7_12_2  (
            .in0(N__29379),
            .in1(N__31764),
            .in2(_gnd_net_),
            .in3(N__57862),
            .lcout(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_7_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_7_12_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_RNII68S_9_LC_7_12_5  (
            .in0(N__57863),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29363),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_10_LC_7_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_10_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_10_LC_7_12_7 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \Commands_frame_decoder.state_10_LC_7_12_7  (
            .in0(N__31765),
            .in1(N__29364),
            .in2(N__29347),
            .in3(N__31305),
            .lcout(\Commands_frame_decoder.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59172),
            .ce(),
            .sr(N__57509));
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_7_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_7_13_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_7_13_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_4_LC_7_13_0  (
            .in0(N__31780),
            .in1(N__29306),
            .in2(N__29547),
            .in3(N__53350),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59185),
            .ce(),
            .sr(N__57513));
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIGK1J_4_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__29513),
            .in2(_gnd_net_),
            .in3(N__31779),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_5_LC_7_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_5_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_5_LC_7_13_2 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \Commands_frame_decoder.state_5_LC_7_13_2  (
            .in0(N__31308),
            .in1(N__29573),
            .in2(N__29577),
            .in3(N__31782),
            .lcout(\Commands_frame_decoder.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59185),
            .ce(),
            .sr(N__57513));
    defparam \Commands_frame_decoder.state_6_LC_7_13_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_6_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_6_LC_7_13_6 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \Commands_frame_decoder.state_6_LC_7_13_6  (
            .in0(N__31309),
            .in1(N__29559),
            .in2(N__29548),
            .in3(N__31783),
            .lcout(\Commands_frame_decoder.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59185),
            .ce(),
            .sr(N__57513));
    defparam \Commands_frame_decoder.state_4_LC_7_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_4_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_4_LC_7_13_7 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \Commands_frame_decoder.state_4_LC_7_13_7  (
            .in0(N__29514),
            .in1(N__31781),
            .in2(N__47946),
            .in3(N__31307),
            .lcout(\Commands_frame_decoder.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59185),
            .ce(),
            .sr(N__57513));
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNID18S_4_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__29502),
            .in2(_gnd_net_),
            .in3(N__57846),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_2_LC_7_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_2_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_2_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_2_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29496),
            .lcout(\pid_front.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59213),
            .ce(N__58507),
            .sr(N__58206));
    defparam \pid_front.error_p_reg_esr_0_LC_7_15_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_0_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_0_LC_7_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_0_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29487),
            .lcout(\pid_front.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59213),
            .ce(N__58507),
            .sr(N__58206));
    defparam \pid_front.error_p_reg_esr_5_LC_7_15_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_5_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_5_LC_7_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_5_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29475),
            .lcout(\pid_front.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59213),
            .ce(N__58507),
            .sr(N__58206));
    defparam \pid_front.error_p_reg_esr_11_LC_7_15_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_11_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_11_LC_7_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_11_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29460),
            .lcout(\pid_front.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59213),
            .ce(N__58507),
            .sr(N__58206));
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52679),
            .lcout(\dron_frame_decoder_1.drone_altitude_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59229),
            .ce(N__30854),
            .sr(N__57526));
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_16_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52361),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59229),
            .ce(N__30854),
            .sr(N__57526));
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_16_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50767),
            .lcout(\dron_frame_decoder_1.drone_altitude_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59229),
            .ce(N__30854),
            .sr(N__57526));
    defparam \dron_frame_decoder_1.state_7_LC_7_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_7_17_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_7_17_0  (
            .in0(N__32142),
            .in1(N__32170),
            .in2(_gnd_net_),
            .in3(N__34698),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59246),
            .ce(),
            .sr(N__57533));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_7_17_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_7_17_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__35810),
            .in2(_gnd_net_),
            .in3(N__35787),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_7_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_7_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30642),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_7_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_7_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30903),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_7_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_7_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30897),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_7_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_7_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29613),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_7_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_7_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30885),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_7_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_7_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30891),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_inv_LC_7_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_7_19_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_7_19_5  (
            .in0(N__42299),
            .in1(N__30655),
            .in2(_gnd_net_),
            .in3(N__29738),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_13_LC_7_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_7_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30873),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_14_LC_7_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_7_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_14_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30879),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_12_LC_7_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_7_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30867),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIM6G7_9_LC_7_21_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIM6G7_9_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIM6G7_9_LC_7_21_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIM6G7_9_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__30825),
            .in2(_gnd_net_),
            .in3(N__30787),
            .lcout(\pid_front.error_p_reg_esr_RNIM6G7Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_2 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29697),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59075),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_8_2_2 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29679),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59076),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_8_2_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29691),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59076),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_2__0__0_LC_8_2_7 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29685),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59076),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_8_5_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_8_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__29799),
            .in2(N__31164),
            .in3(N__31163),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_1_LC_8_5_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_8_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(N__29793),
            .in2(_gnd_net_),
            .in3(N__29787),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_2_LC_8_5_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_8_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__29784),
            .in2(_gnd_net_),
            .in3(N__29778),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_3_LC_8_5_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_8_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__29775),
            .in2(_gnd_net_),
            .in3(N__29769),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_4_LC_8_5_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_8_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__31053),
            .in2(_gnd_net_),
            .in3(N__29766),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_5_LC_8_5_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_8_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__31080),
            .in2(_gnd_net_),
            .in3(N__29763),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_6_LC_8_5_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_8_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__31104),
            .in2(_gnd_net_),
            .in3(N__29760),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_7_LC_8_5_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_8_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(N__31131),
            .in2(_gnd_net_),
            .in3(N__29757),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__59086),
            .ce(),
            .sr(N__29823));
    defparam \Commands_frame_decoder.WDT_8_LC_8_6_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_8_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__31092),
            .in2(_gnd_net_),
            .in3(N__29847),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \Commands_frame_decoder.WDT_9_LC_8_6_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_8_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__31067),
            .in2(_gnd_net_),
            .in3(N__29844),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \Commands_frame_decoder.WDT_10_LC_8_6_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_8_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__31407),
            .in2(_gnd_net_),
            .in3(N__29841),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \Commands_frame_decoder.WDT_11_LC_8_6_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_8_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__31118),
            .in2(_gnd_net_),
            .in3(N__29838),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \Commands_frame_decoder.WDT_12_LC_8_6_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_8_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__31419),
            .in2(_gnd_net_),
            .in3(N__29835),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \Commands_frame_decoder.WDT_13_LC_8_6_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_8_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__31335),
            .in2(_gnd_net_),
            .in3(N__29832),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \Commands_frame_decoder.WDT_14_LC_8_6_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_8_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__31359),
            .in2(_gnd_net_),
            .in3(N__29829),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \Commands_frame_decoder.WDT_15_LC_8_6_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_8_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__31377),
            .in2(_gnd_net_),
            .in3(N__29826),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59092),
            .ce(),
            .sr(N__29819));
    defparam \uart_pc.state_RNO_0_2_LC_8_7_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_8_7_0 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_8_7_0  (
            .in0(N__30144),
            .in1(N__30327),
            .in2(N__30045),
            .in3(N__57878),
            .lcout(),
            .ltout(\uart_pc.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_8_7_1 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_8_7_1 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \uart_pc.state_2_LC_8_7_1  (
            .in0(N__29936),
            .in1(N__30043),
            .in2(N__29802),
            .in3(N__29883),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59100),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_1_LC_8_7_2 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_8_7_2 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.state_1_LC_8_7_2  (
            .in0(N__30044),
            .in1(N__30329),
            .in2(N__30015),
            .in3(N__57879),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59100),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_8_7_3 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_8_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_8_7_3  (
            .in0(N__31140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59100),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_8_7_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_8_7_4 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_drone.timer_Count_3_LC_8_7_4  (
            .in0(N__31509),
            .in1(N__31484),
            .in2(N__57901),
            .in3(N__32500),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59100),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_8_7_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_8_7_5 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_8_7_5  (
            .in0(N__30328),
            .in1(N__57871),
            .in2(_gnd_net_),
            .in3(N__30011),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_8_7_6 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_8_7_6 .LUT_INIT=16'b1010111110001111;
    LogicCell40 \uart_pc.state_0_LC_8_7_6  (
            .in0(N__29972),
            .in1(N__30030),
            .in2(N__30018),
            .in3(N__29935),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59100),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_8_7_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_8_7_7 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_8_7_7  (
            .in0(N__29934),
            .in1(N__30238),
            .in2(N__30148),
            .in3(N__29882),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_8_8_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_8_8_0 .LUT_INIT=16'b0011000100010001;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_8_8_0  (
            .in0(N__30233),
            .in1(N__29968),
            .in2(N__29932),
            .in3(N__29879),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(\uart_pc.un1_state_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_8_8_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_8_8_1 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__30234),
            .in2(N__29940),
            .in3(N__30619),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_8_8_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_8_8_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_8_8_2  (
            .in0(N__30235),
            .in1(N__30149),
            .in2(N__29933),
            .in3(N__29880),
            .lcout(),
            .ltout(\uart_pc.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_8_8_3 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_8_8_3 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \uart_pc.state_3_LC_8_8_3  (
            .in0(N__30159),
            .in1(N__44950),
            .in2(N__30153),
            .in3(N__30150),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59109),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_8_8_4 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_8_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30117),
            .lcout(debug_CH2_18A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59109),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_8_8_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_8_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__31543),
            .in2(_gnd_net_),
            .in3(N__31557),
            .lcout(),
            .ltout(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_8_8_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_8_8_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \uart_drone.timer_Count_1_LC_8_8_6  (
            .in0(N__31482),
            .in1(N__57883),
            .in2(N__30111),
            .in3(N__32504),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59109),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_8_8_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_8_8_7 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \uart_drone.timer_Count_0_LC_8_8_7  (
            .in0(N__57884),
            .in1(N__31544),
            .in2(N__32505),
            .in3(N__31481),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59109),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_8_9_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_8_9_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_0_LC_8_9_0  (
            .in0(N__30591),
            .in1(N__30333),
            .in2(N__30107),
            .in3(N__30378),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.data_Aux_1_LC_8_9_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_8_9_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_pc.data_Aux_1_LC_8_9_1  (
            .in0(N__30374),
            .in1(N__30582),
            .in2(N__30090),
            .in3(N__30338),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.data_Aux_2_LC_8_9_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_8_9_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_2_LC_8_9_2  (
            .in0(N__30573),
            .in1(N__30334),
            .in2(N__30075),
            .in3(N__30379),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.data_Aux_3_LC_8_9_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_8_9_3 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \uart_pc.data_Aux_3_LC_8_9_3  (
            .in0(N__30375),
            .in1(N__30056),
            .in2(N__30441),
            .in3(N__30339),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.data_Aux_4_LC_8_9_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_8_9_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_4_LC_8_9_4  (
            .in0(N__30168),
            .in1(N__30335),
            .in2(N__30429),
            .in3(N__30380),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.data_Aux_5_LC_8_9_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_8_9_5 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \uart_pc.data_Aux_5_LC_8_9_5  (
            .in0(N__30376),
            .in1(N__30407),
            .in2(N__30636),
            .in3(N__30340),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.data_Aux_6_LC_8_9_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_8_9_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_6_LC_8_9_6  (
            .in0(N__30627),
            .in1(N__30336),
            .in2(N__30396),
            .in3(N__30381),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.data_Aux_7_LC_8_9_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_8_9_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_pc.data_Aux_7_LC_8_9_7  (
            .in0(N__30377),
            .in1(N__30337),
            .in2(N__30279),
            .in3(N__30621),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59117),
            .ce(),
            .sr(N__30264));
    defparam \uart_pc.bit_Count_0_LC_8_10_0 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_8_10_0 .LUT_INIT=16'b0000110000101100;
    LogicCell40 \uart_pc.bit_Count_0_LC_8_10_0  (
            .in0(N__30248),
            .in1(N__30527),
            .in2(N__30198),
            .in3(N__30618),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59130),
            .ce(),
            .sr(N__57505));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_8_10_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_8_10_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_8_10_1  (
            .in0(N__30526),
            .in1(N__30193),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uart_pc.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_2_LC_8_10_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_8_10_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_pc.bit_Count_2_LC_8_10_2  (
            .in0(N__30180),
            .in1(N__30564),
            .in2(N__30201),
            .in3(N__30485),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59130),
            .ce(),
            .sr(N__57505));
    defparam \uart_pc.bit_Count_1_LC_8_10_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_8_10_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_pc.bit_Count_1_LC_8_10_3  (
            .in0(N__30528),
            .in1(N__30197),
            .in2(N__30489),
            .in3(N__30179),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59130),
            .ce(),
            .sr(N__57505));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_10_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_10_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_8_10_4  (
            .in0(N__30561),
            .in1(N__30477),
            .in2(_gnd_net_),
            .in3(N__30523),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_10_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_10_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_8_10_5  (
            .in0(N__30524),
            .in1(_gnd_net_),
            .in2(N__30488),
            .in3(N__30563),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_10_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_10_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_8_10_6  (
            .in0(N__30562),
            .in1(N__30481),
            .in2(_gnd_net_),
            .in3(N__30525),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_5_LC_8_11_0 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_8_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_8_11_0  (
            .in0(N__41258),
            .in1(N__41197),
            .in2(_gnd_net_),
            .in3(N__41174),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59144),
            .ce(N__37453),
            .sr(N__57510));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_8_11_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_8_11_1 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_8_11_1  (
            .in0(N__35577),
            .in1(N__35502),
            .in2(N__35430),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_8_11_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_8_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_8_11_3  (
            .in0(N__30556),
            .in1(N__30518),
            .in2(_gnd_net_),
            .in3(N__30468),
            .lcout(\uart_pc.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_8_11_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_8_11_4 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_8_11_4  (
            .in0(N__30519),
            .in1(_gnd_net_),
            .in2(N__30486),
            .in3(N__30557),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_8_11_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_8_11_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_8_11_5  (
            .in0(N__30559),
            .in1(N__30520),
            .in2(_gnd_net_),
            .in3(N__30472),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_8_11_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_8_11_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_8_11_6  (
            .in0(N__30521),
            .in1(_gnd_net_),
            .in2(N__30487),
            .in3(N__30558),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_11_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_11_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_8_11_7  (
            .in0(N__30560),
            .in1(N__30522),
            .in2(_gnd_net_),
            .in3(N__30476),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56454),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59155),
            .ce(N__33077),
            .sr(N__57514));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_8_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_8_13_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_5_LC_8_13_2  (
            .in0(N__55709),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58343),
            .lcout(xy_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59173),
            .ce(N__31925),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_8_13_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_8_13_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_8_13_6  (
            .in0(N__55875),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58342),
            .lcout(xy_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59173),
            .ce(N__31925),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_LC_8_14_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_8_14_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_8_14_3  (
            .in0(N__32213),
            .in1(N__40979),
            .in2(_gnd_net_),
            .in3(N__47661),
            .lcout(debug_CH1_0A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59186),
            .ce(),
            .sr(N__57522));
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__32148),
            .in2(_gnd_net_),
            .in3(N__57847),
            .lcout(\dron_frame_decoder_1.N_513_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_0_LC_8_17_1 .C_ON=1'b0;
    defparam \pid_front.state_0_LC_8_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_0_LC_8_17_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.state_0_LC_8_17_1  (
            .in0(N__50480),
            .in1(N__50611),
            .in2(_gnd_net_),
            .in3(N__47677),
            .lcout(\pid_front.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59230),
            .ce(),
            .sr(N__57539));
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_8_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_8_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_8_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_0_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52259),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59247),
            .ce(N__34946),
            .sr(N__57549));
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_8_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_8_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_1_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50772),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59247),
            .ce(N__34946),
            .sr(N__57549));
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_8_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_8_18_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_8_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_4_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52576),
            .lcout(\dron_frame_decoder_1.drone_altitude_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59247),
            .ce(N__34946),
            .sr(N__57549));
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_8_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_8_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_5_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52457),
            .lcout(\dron_frame_decoder_1.drone_altitude_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59247),
            .ce(N__34946),
            .sr(N__57549));
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_8_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_8_18_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_8_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_6_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53204),
            .lcout(\dron_frame_decoder_1.drone_altitude_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59247),
            .ce(N__34946),
            .sr(N__57549));
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_8_18_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_8_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_7_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52378),
            .lcout(\dron_frame_decoder_1.drone_altitude_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59247),
            .ce(N__34946),
            .sr(N__57549));
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_8_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_8_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_8_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_8_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52273),
            .lcout(\dron_frame_decoder_1.drone_altitude_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59262),
            .ce(N__30850),
            .sr(N__57559));
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_8_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_8_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_8_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_14_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53205),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59262),
            .ce(N__30850),
            .sr(N__57559));
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_8_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_8_19_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_8_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_13_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52468),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59262),
            .ce(N__30850),
            .sr(N__57559));
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_8_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_8_19_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_8_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_12_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52590),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59262),
            .ce(N__30850),
            .sr(N__57559));
    defparam \pid_front.error_d_reg_esr_RNIDQE8_9_LC_8_20_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIDQE8_9_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIDQE8_9_LC_8_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_esr_RNIDQE8_9_LC_8_20_2  (
            .in0(N__56773),
            .in1(N__30824),
            .in2(_gnd_net_),
            .in3(N__30789),
            .lcout(\pid_front.un1_pid_prereg_80_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_9_LC_8_20_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_8_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_8_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_9_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56774),
            .lcout(\pid_front.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59276),
            .ce(N__49364),
            .sr(N__57569));
    defparam \pid_front.error_p_reg_esr_RNIM6G7_0_9_LC_8_20_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIM6G7_0_9_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIM6G7_0_9_LC_8_20_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIM6G7_0_9_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__30823),
            .in2(_gnd_net_),
            .in3(N__30788),
            .lcout(\pid_front.N_1459_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_8_20_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_8_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(N__30918),
            .in2(_gnd_net_),
            .in3(N__33245),
            .lcout(\pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_7_LC_8_21_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_7_LC_8_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_7_LC_8_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_7_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30948),
            .lcout(\pid_front.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59288),
            .ce(N__58449),
            .sr(N__58193));
    defparam \pid_front.error_p_reg_esr_RNII2G7_7_LC_8_21_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNII2G7_7_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNII2G7_7_LC_8_21_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_front.error_p_reg_esr_RNII2G7_7_LC_8_21_1  (
            .in0(N__35128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35037),
            .lcout(),
            .ltout(\pid_front.N_1451_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNINKUF_7_LC_8_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNINKUF_7_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNINKUF_7_LC_8_21_2 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_front.error_d_reg_esr_RNINKUF_7_LC_8_21_2  (
            .in0(N__59397),
            .in1(N__34983),
            .in2(N__30930),
            .in3(N__35010),
            .lcout(\pid_front.error_d_reg_esr_RNINKUFZ0Z_7 ),
            .ltout(\pid_front.error_d_reg_esr_RNINKUFZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJETV_7_LC_8_21_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJETV_7_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJETV_7_LC_8_21_3 .LUT_INIT=16'b0011001110011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJETV_7_LC_8_21_3  (
            .in0(N__35129),
            .in1(N__30924),
            .in2(N__30927),
            .in3(N__35038),
            .lcout(\pid_front.error_p_reg_esr_RNIJETVZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIANE8_8_LC_8_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIANE8_8_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIANE8_8_LC_8_21_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_d_reg_esr_RNIANE8_8_LC_8_21_4  (
            .in0(N__32267),
            .in1(_gnd_net_),
            .in2(N__32310),
            .in3(N__53911),
            .lcout(\pid_front.un1_pid_prereg_70_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK4G7_8_LC_8_21_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK4G7_8_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK4G7_8_LC_8_21_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK4G7_8_LC_8_21_7  (
            .in0(_gnd_net_),
            .in1(N__32305),
            .in2(_gnd_net_),
            .in3(N__32266),
            .lcout(\pid_front.N_1455_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI42GP4_13_LC_8_22_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI42GP4_13_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI42GP4_13_LC_8_22_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI42GP4_13_LC_8_22_0  (
            .in0(N__30961),
            .in1(N__30917),
            .in2(N__33246),
            .in3(N__31001),
            .lcout(\pid_front.error_p_reg_esr_RNI42GP4Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_8_22_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_8_22_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_8_22_1  (
            .in0(N__30987),
            .in1(N__45057),
            .in2(_gnd_net_),
            .in3(N__59466),
            .lcout(\pid_front.un1_pid_prereg_23 ),
            .ltout(\pid_front.un1_pid_prereg_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIN47A4_12_LC_8_22_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN47A4_12_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN47A4_12_LC_8_22_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN47A4_12_LC_8_22_2  (
            .in0(N__33241),
            .in1(N__33189),
            .in2(N__31041),
            .in3(N__32379),
            .lcout(\pid_front.error_p_reg_esr_RNIN47A4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIO6FT1_12_LC_8_22_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO6FT1_12_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO6FT1_12_LC_8_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO6FT1_12_LC_8_22_4  (
            .in0(_gnd_net_),
            .in1(N__33188),
            .in2(_gnd_net_),
            .in3(N__32378),
            .lcout(\pid_front.error_p_reg_esr_RNIO6FT1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBAOC2_15_LC_8_23_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBAOC2_15_LC_8_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBAOC2_15_LC_8_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBAOC2_15_LC_8_23_0  (
            .in0(_gnd_net_),
            .in1(N__33537),
            .in2(_gnd_net_),
            .in3(N__33509),
            .lcout(\pid_front.error_p_reg_esr_RNIBAOC2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_8_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_8_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_8_23_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_15_LC_8_23_1  (
            .in0(N__59360),
            .in1(_gnd_net_),
            .in2(N__31014),
            .in3(N__31035),
            .lcout(\pid_front.un1_pid_prereg_30 ),
            .ltout(\pid_front.un1_pid_prereg_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIGEGP4_14_LC_8_23_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGEGP4_14_LC_8_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGEGP4_14_LC_8_23_2 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGEGP4_14_LC_8_23_2  (
            .in0(N__30963),
            .in1(N__33536),
            .in2(N__31038),
            .in3(N__31002),
            .lcout(\pid_front.error_p_reg_esr_RNIGEGP4Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_15_LC_8_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_8_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_8_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_15_LC_8_23_3  (
            .in0(N__59361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59308),
            .ce(N__49358),
            .sr(N__57594));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_8_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_8_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_8_23_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_8_23_4  (
            .in0(N__31034),
            .in1(N__31010),
            .in2(_gnd_net_),
            .in3(N__59359),
            .lcout(\pid_front.un1_pid_prereg_29 ),
            .ltout(\pid_front.un1_pid_prereg_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI54OC2_14_LC_8_23_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI54OC2_14_LC_8_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI54OC2_14_LC_8_23_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI54OC2_14_LC_8_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30990),
            .in3(N__30962),
            .lcout(\pid_front.error_p_reg_esr_RNI54OC2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_8_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_8_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_8_23_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_14_LC_8_23_6  (
            .in0(N__30986),
            .in1(N__45056),
            .in2(_gnd_net_),
            .in3(N__59459),
            .lcout(\pid_front.un1_pid_prereg_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIPKTD_0_LC_8_27_0 .C_ON=1'b0;
    defparam \pid_front.state_RNIPKTD_0_LC_8_27_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIPKTD_0_LC_8_27_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNIPKTD_0_LC_8_27_0  (
            .in0(_gnd_net_),
            .in1(N__50493),
            .in2(_gnd_net_),
            .in3(N__57833),
            .lcout(\pid_front.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_7 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_9_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31191),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59074),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_1__0__0_LC_9_3_5 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31185),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59077),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.Q_0__0_LC_9_5_1 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_9_5_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__31176),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(debug_CH0_16A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59083),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI1NQ51_15_LC_9_5_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI1NQ51_15_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI1NQ51_15_LC_9_5_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI1NQ51_15_LC_9_5_2  (
            .in0(N__31375),
            .in1(N__31356),
            .in2(_gnd_net_),
            .in3(N__31333),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIGA2K5_LC_9_5_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIGA2K5_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIGA2K5_LC_9_5_3 .LUT_INIT=16'b0011000000110001;
    LogicCell40 \Commands_frame_decoder.preinit_RNIGA2K5_LC_9_5_3  (
            .in0(N__31357),
            .in1(N__31435),
            .in2(N__31167),
            .in3(N__31383),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_9_5_6 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_9_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31149),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59083),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI8EBE1_6_LC_9_6_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI8EBE1_6_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI8EBE1_6_LC_9_6_1 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI8EBE1_6_LC_9_6_1  (
            .in0(N__31405),
            .in1(N__31130),
            .in2(N__31119),
            .in3(N__31103),
            .lcout(\Commands_frame_decoder.WDT8lto15_N_5L7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_9_6_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_9_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNII19A1_4_LC_9_6_3  (
            .in0(N__31091),
            .in1(N__31079),
            .in2(N__31068),
            .in3(N__31052),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIAERH3_12_LC_9_6_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIAERH3_12_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIAERH3_12_LC_9_6_4 .LUT_INIT=16'b1010111011111111;
    LogicCell40 \Commands_frame_decoder.WDT_RNIAERH3_12_LC_9_6_4  (
            .in0(N__31418),
            .in1(N__31406),
            .in2(N__31392),
            .in3(N__31389),
            .lcout(\Commands_frame_decoder.WDT_RNIAERH3Z0Z_12 ),
            .ltout(\Commands_frame_decoder.WDT_RNIAERH3Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIB5MN4_15_LC_9_6_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIB5MN4_15_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIB5MN4_15_LC_9_6_5 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIB5MN4_15_LC_9_6_5  (
            .in0(N__31376),
            .in1(N__31358),
            .in2(N__31338),
            .in3(N__31334),
            .lcout(\Commands_frame_decoder.WDT8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_LC_9_6_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_9_6_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_9_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__31775),
            .in2(_gnd_net_),
            .in3(N__31436),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59087),
            .ce(),
            .sr(N__57499));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_0 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__33825),
            .in2(_gnd_net_),
            .in3(N__31457),
            .lcout(\uart_drone.N_126_li ),
            .ltout(\uart_drone.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_7_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_7_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_9_7_1  (
            .in0(N__33788),
            .in1(N__32606),
            .in2(N__31209),
            .in3(N__57856),
            .lcout(\uart_drone.N_143 ),
            .ltout(\uart_drone.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_9_7_2 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_9_7_2 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \uart_drone.state_4_LC_9_7_2  (
            .in0(N__33741),
            .in1(N__33930),
            .in2(N__31206),
            .in3(N__44928),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59093),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_9_7_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_9_7_3 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_9_7_3  (
            .in0(N__32624),
            .in1(N__33928),
            .in2(N__31524),
            .in3(N__32607),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_9_7_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_9_7_6 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_drone.timer_Count_4_LC_9_7_6  (
            .in0(N__57857),
            .in1(N__31497),
            .in2(N__32490),
            .in3(N__31485),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59093),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_9_7_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_9_7_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_9_7_7  (
            .in0(N__33929),
            .in1(N__32608),
            .in2(_gnd_net_),
            .in3(N__57855),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_9_8_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_9_8_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_9_8_0  (
            .in0(N__31539),
            .in1(N__31556),
            .in2(N__31545),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_9_8_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_9_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31458),
            .in3(N__31512),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_9_8_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_9_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33836),
            .in3(N__31503),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_9_8_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_9_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__33776),
            .in2(_gnd_net_),
            .in3(N__31500),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_9_8_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_9_8_5 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_drone.timer_Count_2_LC_9_8_5  (
            .in0(N__31491),
            .in1(N__31483),
            .in2(N__57903),
            .in3(N__32491),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59101),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_8_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_8_6 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_9_8_6  (
            .in0(N__33821),
            .in1(N__31453),
            .in2(N__33789),
            .in3(N__32602),
            .lcout(\uart_drone.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_rdy_LC_9_9_4 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_9_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.data_rdy_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__32897),
            .in2(_gnd_net_),
            .in3(N__31885),
            .lcout(uart_drone_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59110),
            .ce(),
            .sr(N__57506));
    defparam \Commands_frame_decoder.source_data_valid_LC_9_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_9_9_7 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_9_9_7  (
            .in0(N__31818),
            .in1(N__31776),
            .in2(N__41009),
            .in3(N__31440),
            .lcout(debug_CH3_20A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59110),
            .ce(),
            .sr(N__57506));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_10_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_10_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_9_10_2  (
            .in0(N__32864),
            .in1(N__31886),
            .in2(_gnd_net_),
            .in3(N__57859),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_10_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_10_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_9_10_3  (
            .in0(N__31887),
            .in1(_gnd_net_),
            .in2(N__31869),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_rdyc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__31865),
            .in2(_gnd_net_),
            .in3(N__31845),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_esr_3_LC_9_11_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_9_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_3_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32643),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59131),
            .ce(N__32997),
            .sr(N__32985));
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_9_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_9_12_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNITUI31_13_LC_9_12_0  (
            .in0(N__31812),
            .in1(N__31784),
            .in2(_gnd_net_),
            .in3(N__57832),
            .lcout(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_9_12_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_9_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_9_12_6  (
            .in0(N__32955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40943),
            .lcout(\dron_frame_decoder_1.N_224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_1_LC_9_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_9_13_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_9_13_2  (
            .in0(N__34678),
            .in1(N__32945),
            .in2(N__31569),
            .in3(N__31578),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59156),
            .ce(),
            .sr(N__57523));
    defparam \dron_frame_decoder_1.state_ns_0_a3_0_1_1_LC_9_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_a3_0_1_1_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_a3_0_1_1_LC_9_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_a3_0_1_1_LC_9_13_3  (
            .in0(N__53184),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52541),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_a3_0_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_9_13_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_9_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_9_13_4  (
            .in0(N__52649),
            .in1(N__31909),
            .in2(N__31581),
            .in3(N__50749),
            .lcout(\dron_frame_decoder_1.N_220 ),
            .ltout(\dron_frame_decoder_1.N_220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_9_13_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_9_13_5 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_9_13_5  (
            .in0(N__33060),
            .in1(N__31893),
            .in2(N__31572),
            .in3(N__31565),
            .lcout(),
            .ltout(\dron_frame_decoder_1.N_198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_0_LC_9_13_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_9_13_6 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_9_13_6 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_9_13_6  (
            .in0(N__34679),
            .in1(N__32121),
            .in2(N__32124),
            .in3(N__31913),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59156),
            .ce(),
            .sr(N__57523));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_7  (
            .in0(N__40968),
            .in1(N__32941),
            .in2(N__31914),
            .in3(N__32214),
            .lcout(\dron_frame_decoder_1.N_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_0_LC_9_14_0  (
            .in0(N__56466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58337),
            .lcout(xy_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59174),
            .ce(N__31932),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_1_LC_9_14_1  (
            .in0(N__58338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56271),
            .lcout(xy_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59174),
            .ce(N__31932),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_2_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__56110),
            .in2(_gnd_net_),
            .in3(N__58339),
            .lcout(xy_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59174),
            .ce(N__31932),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_3_LC_9_14_3  (
            .in0(N__58340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55342),
            .lcout(xy_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59174),
            .ce(N__31932),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_6_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__55548),
            .in2(_gnd_net_),
            .in3(N__58341),
            .lcout(xy_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59174),
            .ce(N__31932),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_9_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_9_14_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \dron_frame_decoder_1.state_RNO_2_0_LC_9_14_7  (
            .in0(N__32206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31908),
            .lcout(\dron_frame_decoder_1.state_ns_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_6_LC_9_15_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_9_15_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_9_15_6  (
            .in0(N__32212),
            .in1(N__40980),
            .in2(N__32178),
            .in3(N__34694),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59187),
            .ce(),
            .sr(N__57534));
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_9_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_9_16_1 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \dron_frame_decoder_1.state_RNI0TLI1_4_LC_9_16_1  (
            .in0(N__32208),
            .in1(N__33144),
            .in2(N__57900),
            .in3(N__33108),
            .lcout(\dron_frame_decoder_1.N_521_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_16_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_16_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_9_16_3  (
            .in0(N__32207),
            .in1(N__33107),
            .in2(N__32177),
            .in3(N__33143),
            .lcout(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__33109),
            .in2(_gnd_net_),
            .in3(N__40981),
            .lcout(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ),
            .ltout(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_9_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_9_17_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \dron_frame_decoder_1.state_RNI36DT_4_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32133),
            .in3(N__57850),
            .lcout(\dron_frame_decoder_1.N_505_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI4KF7_0_0_LC_9_17_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI4KF7_0_0_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI4KF7_0_0_LC_9_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI4KF7_0_0_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__38386),
            .in2(_gnd_net_),
            .in3(N__38352),
            .lcout(\pid_front.un1_pid_prereg_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_8_LC_9_18_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_9_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_8_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53915),
            .lcout(\pid_front.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59231),
            .ce(N__49370),
            .sr(N__57560));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_9_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_9_19_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__32130),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_9_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_9_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50768),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59248),
            .ce(N__53117),
            .sr(N__57570));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_9_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50384),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59248),
            .ce(N__53117),
            .sr(N__57570));
    defparam \pid_alt.error_axb_1_LC_9_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_9_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_1_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32325),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNITOTV_8_LC_9_20_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITOTV_8_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITOTV_8_LC_9_20_6 .LUT_INIT=16'b0100101101001011;
    LogicCell40 \pid_front.error_p_reg_esr_RNITOTV_8_LC_9_20_6  (
            .in0(N__32309),
            .in1(N__32262),
            .in2(N__32235),
            .in3(N__36488),
            .lcout(\pid_front.error_p_reg_esr_RNITOTVZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNISPUF_8_LC_9_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNISPUF_8_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNISPUF_8_LC_9_21_4 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \pid_front.error_d_reg_esr_RNISPUF_8_LC_9_21_4  (
            .in0(N__32226),
            .in1(N__35039),
            .in2(N__53916),
            .in3(N__35130),
            .lcout(\pid_front.error_d_reg_esr_RNISPUFZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI57KP4_18_LC_9_21_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI57KP4_18_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI57KP4_18_LC_9_21_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI57KP4_18_LC_9_21_7  (
            .in0(N__32403),
            .in1(N__32421),
            .in2(N__42636),
            .in3(N__33293),
            .lcout(\pid_front.error_p_reg_esr_RNI57KP4Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIO6FT1_0_12_LC_9_22_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO6FT1_0_12_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO6FT1_0_12_LC_9_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO6FT1_0_12_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__33182),
            .in2(_gnd_net_),
            .in3(N__32377),
            .lcout(\pid_front.error_p_reg_esr_RNIO6FT1_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_22_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_22_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_22_4  (
            .in0(N__33968),
            .in1(N__46850),
            .in2(_gnd_net_),
            .in3(N__56815),
            .lcout(\pid_front.error_p_reg_esr_RNI8NB61Z0Z_11 ),
            .ltout(\pid_front.error_p_reg_esr_RNI8NB61Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIBO6A4_12_LC_9_22_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIBO6A4_12_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIBO6A4_12_LC_9_22_5 .LUT_INIT=16'b1011001010110010;
    LogicCell40 \pid_front.error_d_reg_esr_RNIBO6A4_12_LC_9_22_5  (
            .in0(N__53853),
            .in1(N__32388),
            .in2(N__32220),
            .in3(N__36983),
            .lcout(\pid_front.error_d_reg_esr_RNIBO6A4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_9_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_9_23_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_19_LC_9_23_1  (
            .in0(N__32441),
            .in1(N__32450),
            .in2(_gnd_net_),
            .in3(N__59527),
            .lcout(\pid_front.un1_pid_prereg_57 ),
            .ltout(\pid_front.un1_pid_prereg_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8ARC2_19_LC_9_23_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8ARC2_19_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8ARC2_19_LC_9_23_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8ARC2_19_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32217),
            .in3(N__42628),
            .lcout(\pid_front.error_p_reg_esr_RNI8ARC2Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_19_LC_9_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_9_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_19_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59529),
            .lcout(\pid_front.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59301),
            .ce(N__49360),
            .sr(N__57601));
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_9_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_9_23_4 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_18_LC_9_23_4  (
            .in0(N__33276),
            .in1(_gnd_net_),
            .in2(N__49404),
            .in3(N__59572),
            .lcout(\pid_front.un1_pid_prereg_48 ),
            .ltout(\pid_front.un1_pid_prereg_48_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIKJHP4_17_LC_9_23_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKJHP4_17_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKJHP4_17_LC_9_23_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKJHP4_17_LC_9_23_5  (
            .in0(N__33621),
            .in1(N__33609),
            .in2(N__32457),
            .in3(N__32417),
            .lcout(\pid_front.error_p_reg_esr_RNIKJHP4Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_9_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_9_23_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_9_23_6  (
            .in0(N__59528),
            .in1(_gnd_net_),
            .in2(N__32454),
            .in3(N__32442),
            .lcout(\pid_front.un1_pid_prereg_56 ),
            .ltout(\pid_front.un1_pid_prereg_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNITSOC2_18_LC_9_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITSOC2_18_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITSOC2_18_LC_9_23_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNITSOC2_18_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32406),
            .in3(N__32399),
            .lcout(\pid_front.error_p_reg_esr_RNITSOC2Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIA93N_0_12_LC_9_24_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIA93N_0_12_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIA93N_0_12_LC_9_24_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIA93N_0_12_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__32347),
            .in2(_gnd_net_),
            .in3(N__32359),
            .lcout(\pid_front.N_1471_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_12_LC_9_24_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_9_24_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_9_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_12_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53849),
            .lcout(\pid_front.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59309),
            .ce(N__49359),
            .sr(N__57609));
    defparam \pid_front.error_p_reg_esr_RNIA93N_12_LC_9_24_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIA93N_12_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIA93N_12_LC_9_24_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIA93N_12_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__32348),
            .in2(_gnd_net_),
            .in3(N__32360),
            .lcout(\pid_front.error_p_reg_esr_RNIA93NZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBQB61_12_LC_9_24_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBQB61_12_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBQB61_12_LC_9_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBQB61_12_LC_9_24_4  (
            .in0(N__32361),
            .in1(N__53848),
            .in2(_gnd_net_),
            .in3(N__32349),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_107_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI1E6A4_12_LC_9_24_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI1E6A4_12_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI1E6A4_12_LC_9_24_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI1E6A4_12_LC_9_24_5  (
            .in0(N__35676),
            .in1(N__35661),
            .in2(N__32328),
            .in3(N__32544),
            .lcout(\pid_front.error_p_reg_esr_RNI1E6A4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_3_LC_10_5_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_10_5_0 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_10_5_0  (
            .in0(N__33852),
            .in1(N__33911),
            .in2(N__33797),
            .in3(N__32525),
            .lcout(),
            .ltout(\uart_drone.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_10_5_1 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_10_5_1 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_drone.state_3_LC_10_5_1  (
            .in0(N__32526),
            .in1(N__33734),
            .in2(N__32535),
            .in3(N__44966),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59078),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI62411_4_LC_10_5_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_10_5_3 .LUT_INIT=16'b0100010100000101;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_10_5_3  (
            .in0(N__32610),
            .in1(N__33790),
            .in2(N__33919),
            .in3(N__33851),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(\uart_drone.un1_state_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI63LK2_3_LC_10_5_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_5_4 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_10_5_4  (
            .in0(_gnd_net_),
            .in1(N__33910),
            .in2(N__32532),
            .in3(N__35615),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_10_6_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_10_6_0 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_10_6_0  (
            .in0(N__32519),
            .in1(N__32860),
            .in2(N__32568),
            .in3(N__57876),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_10_6_1 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_10_6_1 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_drone.state_2_LC_10_6_1  (
            .in0(N__32567),
            .in1(N__33787),
            .in2(N__32529),
            .in3(N__33859),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59081),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_10_6_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_10_6_3 .LUT_INIT=16'b0011111100101010;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_10_6_3  (
            .in0(N__33912),
            .in1(N__33785),
            .in2(N__33861),
            .in3(N__32518),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_6_4 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_6_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__33874),
            .in2(_gnd_net_),
            .in3(N__35407),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_10_6_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_10_6_5 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_10_6_5  (
            .in0(N__57875),
            .in1(N__32576),
            .in2(_gnd_net_),
            .in3(N__32859),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_10_6_6 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_10_6_6 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_drone.state_0_LC_10_6_6  (
            .in0(N__33786),
            .in1(N__32625),
            .in2(N__32613),
            .in3(N__32609),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59081),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_10_6_7 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_10_6_7 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_drone.state_1_LC_10_6_7  (
            .in0(N__57877),
            .in1(N__32566),
            .in2(N__32888),
            .in3(N__32577),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59081),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_10_7_0 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_10_7_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_10_7_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \reset_module_System.count_2_LC_10_7_0  (
            .in0(N__32688),
            .in1(N__32676),
            .in2(N__34266),
            .in3(N__33669),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59084),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_10_7_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_10_7_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_10_7_2  (
            .in0(N__35538),
            .in1(N__35465),
            .in2(_gnd_net_),
            .in3(N__35406),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_10_7_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_10_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_10_7_3  (
            .in0(N__34022),
            .in1(N__34037),
            .in2(N__34008),
            .in3(N__34067),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_10_7_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_10_7_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_10_7_4  (
            .in0(N__34053),
            .in1(N__33660),
            .in2(N__34092),
            .in3(N__33681),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(\reset_module_System.reset6_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_10_7_5 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_10_7_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_10_7_5 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_10_7_5  (
            .in0(N__33704),
            .in1(N__34261),
            .in2(N__32550),
            .in3(N__32686),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59084),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_10_7_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_10_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__33703),
            .in2(_gnd_net_),
            .in3(N__33723),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_10_7_7 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_10_7_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_10_7_7  (
            .in0(N__32675),
            .in1(N__34262),
            .in2(N__32547),
            .in3(N__32687),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59084),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_10_8_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_10_8_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_10_8_0  (
            .in0(N__35486),
            .in1(N__35560),
            .in2(_gnd_net_),
            .in3(N__35421),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIR9N6_1_LC_10_8_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIR9N6_1_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIR9N6_1_LC_10_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIR9N6_1_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__33644),
            .in2(_gnd_net_),
            .in3(N__33721),
            .lcout(),
            .ltout(\reset_module_System.reset6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIA72I1_16_LC_10_8_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIA72I1_16_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIA72I1_16_LC_10_8_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \reset_module_System.count_RNIA72I1_16_LC_10_8_2  (
            .in0(N__34109),
            .in1(N__34127),
            .in2(N__32700),
            .in3(N__32697),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIMJ304_12_LC_10_8_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIMJ304_12_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIMJ304_12_LC_10_8_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIMJ304_12_LC_10_8_3  (
            .in0(N__33984),
            .in1(N__33702),
            .in2(N__32691),
            .in3(N__34194),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_10_8_4 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_10_8_4 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \reset_module_System.reset_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__32674),
            .in2(N__32661),
            .in3(N__34250),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59089),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_10_8_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_10_8_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_10_8_5  (
            .in0(N__35420),
            .in1(_gnd_net_),
            .in2(N__35572),
            .in3(N__35487),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_0_LC_10_9_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_10_9_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_0_LC_10_9_0  (
            .in0(N__32658),
            .in1(N__32889),
            .in2(N__32778),
            .in3(N__32820),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_Aux_1_LC_10_9_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_10_9_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_1_LC_10_9_1  (
            .in0(N__32894),
            .in1(N__34320),
            .in2(N__32763),
            .in3(N__32816),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_Aux_2_LC_10_9_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_10_9_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_2_LC_10_9_2  (
            .in0(N__32652),
            .in1(N__32890),
            .in2(N__32748),
            .in3(N__32821),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_Aux_3_LC_10_9_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_10_9_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_3_LC_10_9_3  (
            .in0(N__32895),
            .in1(N__35349),
            .in2(N__32642),
            .in3(N__32817),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_Aux_4_LC_10_9_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_10_9_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_4_LC_10_9_4  (
            .in0(N__32964),
            .in1(N__32891),
            .in2(N__32718),
            .in3(N__32822),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_Aux_5_LC_10_9_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_10_9_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_5_LC_10_9_5  (
            .in0(N__32896),
            .in1(N__32925),
            .in2(N__32733),
            .in3(N__32818),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_Aux_6_LC_10_9_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_10_9_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_6_LC_10_9_6  (
            .in0(N__32913),
            .in1(N__32892),
            .in2(N__33027),
            .in3(N__32823),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_Aux_7_LC_10_9_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_10_9_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_10_9_7  (
            .in0(N__32893),
            .in1(N__32819),
            .in2(N__33012),
            .in3(N__35616),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59095),
            .ce(),
            .sr(N__32790));
    defparam \uart_drone.data_esr_0_LC_10_10_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_10_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32777),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59103),
            .ce(N__32996),
            .sr(N__32981));
    defparam \uart_drone.data_esr_1_LC_10_10_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_10_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32762),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59103),
            .ce(N__32996),
            .sr(N__32981));
    defparam \uart_drone.data_esr_2_LC_10_10_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_10_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32747),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59103),
            .ce(N__32996),
            .sr(N__32981));
    defparam \uart_drone.data_esr_5_LC_10_10_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_5_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32732),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59103),
            .ce(N__32996),
            .sr(N__32981));
    defparam \uart_drone.data_esr_4_LC_10_10_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_10_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32714),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59103),
            .ce(N__32996),
            .sr(N__32981));
    defparam \uart_drone.data_esr_6_LC_10_10_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_10_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33026),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59103),
            .ce(N__32996),
            .sr(N__32981));
    defparam \uart_drone.data_esr_7_LC_10_10_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33011),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59103),
            .ce(N__32996),
            .sr(N__32981));
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_10_11_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_10_11_0 .LUT_INIT=16'b0000001100010011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_10_11_0  (
            .in0(N__34464),
            .in1(N__40944),
            .in2(N__34560),
            .in3(N__34580),
            .lcout(\dron_frame_decoder_1.N_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_10_11_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_10_11_1 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_10_11_1  (
            .in0(N__34579),
            .in1(N__34555),
            .in2(_gnd_net_),
            .in3(N__34463),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_10_11_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_10_11_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_10_11_4  (
            .in0(N__35422),
            .in1(N__35576),
            .in2(_gnd_net_),
            .in3(N__35498),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_11_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_10_11_5  (
            .in0(N__52426),
            .in1(N__52247),
            .in2(N__52347),
            .in3(N__50336),
            .lcout(\dron_frame_decoder_1.N_263_5 ),
            .ltout(\dron_frame_decoder_1.N_263_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_10_11_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_10_11_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_3_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__40945),
            .in2(N__32949),
            .in3(N__32946),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_10_11_7 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_10_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.source_data_1_esr_ctle_14_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__41008),
            .in2(_gnd_net_),
            .in3(N__57849),
            .lcout(\scaler_4.debug_CH3_20A_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_10_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_10_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_10_12_0  (
            .in0(N__56105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59119),
            .ce(N__33081),
            .sr(N__57518));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_10_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56270),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59119),
            .ce(N__33081),
            .sr(N__57518));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_10_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55730),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59119),
            .ce(N__33081),
            .sr(N__57518));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_10_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_10_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_10_12_3  (
            .in0(N__55343),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59119),
            .ce(N__33081),
            .sr(N__57518));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_10_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_10_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53370),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59119),
            .ce(N__33081),
            .sr(N__57518));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_10_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_10_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55898),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59119),
            .ce(N__33081),
            .sr(N__57518));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_10_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_10_12_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55541),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59119),
            .ce(N__33081),
            .sr(N__57518));
    defparam \dron_frame_decoder_1.state_ns_i_a2_0_4_0_LC_10_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_0_4_0_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_0_4_0_LC_10_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_0_4_0_LC_10_13_0  (
            .in0(N__50731),
            .in1(N__53185),
            .in2(N__52663),
            .in3(N__52542),
            .lcout(\dron_frame_decoder_1.N_219_4 ),
            .ltout(\dron_frame_decoder_1.N_219_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_3_LC_10_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_10_13_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_10_13_1  (
            .in0(N__34366),
            .in1(N__34677),
            .in2(N__33051),
            .in3(N__33048),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59132),
            .ce(),
            .sr(N__57524));
    defparam \ppm_encoder_1.rudder_esr_5_LC_10_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_10_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33039),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59146),
            .ce(N__46763),
            .sr(N__57527));
    defparam \pid_front.error_p_reg_esr_1_LC_10_15_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_1_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_1_LC_10_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_1_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33153),
            .lcout(\pid_front.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59158),
            .ce(N__58503),
            .sr(N__58197));
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_10_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_10_16_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \dron_frame_decoder_1.state_RNI7Q6K_5_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__40964),
            .in2(_gnd_net_),
            .in3(N__33129),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_5_LC_10_16_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_10_16_4 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_10_16_4  (
            .in0(N__34693),
            .in1(_gnd_net_),
            .in2(N__33135),
            .in3(N__36174),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59175),
            .ce(),
            .sr(N__57540));
    defparam \dron_frame_decoder_1.state_4_LC_10_16_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_10_16_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_10_16_5  (
            .in0(N__40970),
            .in1(N__33131),
            .in2(N__33117),
            .in3(N__34692),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59175),
            .ce(),
            .sr(N__57540));
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_10_16_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_10_16_7 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \dron_frame_decoder_1.state_RNI1H181_5_LC_10_16_7  (
            .in0(N__40969),
            .in1(N__33130),
            .in2(N__33116),
            .in3(N__57848),
            .lcout(\dron_frame_decoder_1.N_497_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_16_LC_10_17_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_10_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_16_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56727),
            .lcout(\pid_front.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59189),
            .ce(N__49371),
            .sr(N__57550));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33087),
            .lcout(drone_H_disp_side_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_10_LC_10_19_0 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_10_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_10_LC_10_19_0 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_front.source_pid_1_10_LC_10_19_0  (
            .in0(N__50605),
            .in1(N__35271),
            .in2(N__37915),
            .in3(N__36378),
            .lcout(front_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59214),
            .ce(),
            .sr(N__35189));
    defparam \pid_front.source_pid_1_11_LC_10_19_1 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_11_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_11_LC_10_19_1 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_front.source_pid_1_11_LC_10_19_1  (
            .in0(N__35272),
            .in1(N__50608),
            .in2(N__37873),
            .in3(N__37062),
            .lcout(front_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59214),
            .ce(),
            .sr(N__35189));
    defparam \pid_front.source_pid_1_6_LC_10_19_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_6_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_6_LC_10_19_2 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_front.source_pid_1_6_LC_10_19_2  (
            .in0(N__50606),
            .in1(N__35273),
            .in2(N__37681),
            .in3(N__36633),
            .lcout(front_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59214),
            .ce(),
            .sr(N__35189));
    defparam \pid_front.source_pid_1_7_LC_10_19_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_7_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_7_LC_10_19_3 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_front.source_pid_1_7_LC_10_19_3  (
            .in0(N__35274),
            .in1(N__50609),
            .in2(N__40291),
            .in3(N__36585),
            .lcout(front_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59214),
            .ce(),
            .sr(N__35189));
    defparam \pid_front.source_pid_1_8_LC_10_19_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_8_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_8_LC_10_19_4 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_front.source_pid_1_8_LC_10_19_4  (
            .in0(N__50607),
            .in1(N__35275),
            .in2(N__37993),
            .in3(N__36525),
            .lcout(front_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59214),
            .ce(),
            .sr(N__35189));
    defparam \pid_front.source_pid_1_9_LC_10_19_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_9_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_9_LC_10_19_5 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_front.source_pid_1_9_LC_10_19_5  (
            .in0(N__35276),
            .in1(N__50610),
            .in2(N__37954),
            .in3(N__36459),
            .lcout(front_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59214),
            .ce(),
            .sr(N__35189));
    defparam \pid_front.pid_prereg_esr_RNI6DCJ3_13_LC_10_20_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI6DCJ3_13_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI6DCJ3_13_LC_10_20_0 .LUT_INIT=16'b1010101011111010;
    LogicCell40 \pid_front.pid_prereg_esr_RNI6DCJ3_13_LC_10_20_0  (
            .in0(N__37141),
            .in1(_gnd_net_),
            .in2(N__35331),
            .in3(N__36956),
            .lcout(\pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13 ),
            .ltout(\pid_front.pid_prereg_esr_RNI6DCJ3Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNICUKFA_6_LC_10_20_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNICUKFA_6_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNICUKFA_6_LC_10_20_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNICUKFA_6_LC_10_20_1  (
            .in0(N__35085),
            .in1(N__35076),
            .in2(N__33171),
            .in3(N__33630),
            .lcout(),
            .ltout(\pid_front.pid_prereg_esr_RNICUKFAZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIC8N8C_5_LC_10_20_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIC8N8C_5_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIC8N8C_5_LC_10_20_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIC8N8C_5_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__33441),
            .in2(N__33168),
            .in3(N__33162),
            .lcout(\pid_front.un1_reset_0_i ),
            .ltout(\pid_front.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI9HEDC_1_LC_10_20_3 .C_ON=1'b0;
    defparam \pid_front.state_RNI9HEDC_1_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI9HEDC_1_LC_10_20_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_front.state_RNI9HEDC_1_LC_10_20_3  (
            .in0(N__50624),
            .in1(_gnd_net_),
            .in2(N__33165),
            .in3(_gnd_net_),
            .lcout(\pid_front.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIKVDO_23_LC_10_20_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIKVDO_23_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIKVDO_23_LC_10_20_4 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIKVDO_23_LC_10_20_4  (
            .in0(N__37142),
            .in1(N__50622),
            .in2(_gnd_net_),
            .in3(N__57831),
            .lcout(\pid_front.un1_reset_0_i_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI86GE_2_LC_10_20_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI86GE_2_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI86GE_2_LC_10_20_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNI86GE_2_LC_10_20_5  (
            .in0(N__36336),
            .in1(N__49427),
            .in2(N__36780),
            .in3(N__50441),
            .lcout(),
            .ltout(\pid_front.m32_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNICAK01_5_LC_10_20_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNICAK01_5_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNICAK01_5_LC_10_20_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNICAK01_5_LC_10_20_6  (
            .in0(N__36678),
            .in1(N__50623),
            .in2(N__33156),
            .in3(N__44984),
            .lcout(\pid_front.un1_reset_0_i_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_5_LC_10_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_5_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_5_LC_10_21_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \pid_alt.error_i_acumm_5_LC_10_21_0  (
            .in0(N__33356),
            .in1(N__39675),
            .in2(N__33435),
            .in3(N__33402),
            .lcout(\pid_alt.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59249),
            .ce(),
            .sr(N__33342));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_10_21_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_10_21_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_10_21_1  (
            .in0(N__33581),
            .in1(N__33554),
            .in2(_gnd_net_),
            .in3(N__56723),
            .lcout(\pid_front.un1_pid_prereg_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIOUOP4_19_LC_10_21_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIOUOP4_19_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIOUOP4_19_LC_10_21_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIOUOP4_19_LC_10_21_3  (
            .in0(N__42562),
            .in1(N__42635),
            .in2(N__33300),
            .in3(N__42634),
            .lcout(\pid_front.error_p_reg_esr_RNIOUOP4Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI09RP4_20_LC_10_21_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI09RP4_20_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI09RP4_20_LC_10_21_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI09RP4_20_LC_10_21_4  (
            .in0(N__42566),
            .in1(N__42633),
            .in2(N__42567),
            .in3(N__42632),
            .lcout(\pid_front.error_p_reg_esr_RNI09RP4Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_10_21_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_10_21_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_10_21_7  (
            .in0(N__33272),
            .in1(N__49400),
            .in2(_gnd_net_),
            .in3(N__59574),
            .lcout(\pid_front.un1_pid_prereg_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_10_22_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_10_22_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_13_LC_10_22_1  (
            .in0(N__33219),
            .in1(N__56849),
            .in2(_gnd_net_),
            .in3(N__33198),
            .lcout(\pid_front.un1_pid_prereg_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_13_LC_10_22_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_10_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_10_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_13_LC_10_22_2  (
            .in0(N__56850),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59264),
            .ce(N__49363),
            .sr(N__57595));
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_22_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_22_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_22_3  (
            .in0(N__33218),
            .in1(N__56848),
            .in2(_gnd_net_),
            .in3(N__33197),
            .lcout(\pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI6FQ75_23_LC_10_22_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI6FQ75_23_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI6FQ75_23_LC_10_22_7 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \pid_front.pid_prereg_esr_RNI6FQ75_23_LC_10_22_7  (
            .in0(N__37140),
            .in1(N__36732),
            .in2(N__35094),
            .in3(N__35318),
            .lcout(\pid_front.pid_prereg_esr_RNI6FQ75Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNINMOC2_17_LC_10_23_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNINMOC2_17_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNINMOC2_17_LC_10_23_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNINMOC2_17_LC_10_23_0  (
            .in0(N__33604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33620),
            .lcout(\pid_front.error_p_reg_esr_RNINMOC2Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_10_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_10_23_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_10_23_1  (
            .in0(N__56672),
            .in1(_gnd_net_),
            .in2(N__33477),
            .in3(N__33498),
            .lcout(\pid_front.un1_pid_prereg_42 ),
            .ltout(\pid_front.un1_pid_prereg_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI87HP4_16_LC_10_23_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI87HP4_16_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI87HP4_16_LC_10_23_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI87HP4_16_LC_10_23_2  (
            .in0(N__33605),
            .in1(N__33453),
            .in2(N__33585),
            .in3(N__33465),
            .lcout(\pid_front.error_p_reg_esr_RNI87HP4Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_17_LC_10_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_10_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_17_LC_10_23_3  (
            .in0(N__56673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59277),
            .ce(N__49361),
            .sr(N__57602));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_10_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_10_23_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_16_LC_10_23_4  (
            .in0(N__33582),
            .in1(N__33558),
            .in2(_gnd_net_),
            .in3(N__56710),
            .lcout(\pid_front.un1_pid_prereg_36 ),
            .ltout(\pid_front.un1_pid_prereg_36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNISQGP4_15_LC_10_23_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNISQGP4_15_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNISQGP4_15_LC_10_23_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNISQGP4_15_LC_10_23_5  (
            .in0(N__33464),
            .in1(N__33535),
            .in2(N__33516),
            .in3(N__33513),
            .lcout(\pid_front.error_p_reg_esr_RNISQGP4Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_10_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_10_23_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_10_23_6  (
            .in0(N__33497),
            .in1(N__33473),
            .in2(_gnd_net_),
            .in3(N__56671),
            .lcout(\pid_front.un1_pid_prereg_41 ),
            .ltout(\pid_front.un1_pid_prereg_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIHGOC2_16_LC_10_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIHGOC2_16_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIHGOC2_16_LC_10_23_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIHGOC2_16_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33456),
            .in3(N__33452),
            .lcout(\pid_front.error_p_reg_esr_RNIHGOC2Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_10_24_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_10_24_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_10_24_0  (
            .in0(N__33969),
            .in1(N__46851),
            .in2(_gnd_net_),
            .in3(N__56823),
            .lcout(\pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_1_LC_11_6_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_11_6_2 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uart_drone.bit_Count_1_LC_11_6_2  (
            .in0(N__35483),
            .in1(N__35408),
            .in2(N__33882),
            .in3(N__33944),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59079),
            .ce(),
            .sr(N__57500));
    defparam \uart_drone.bit_Count_2_LC_11_6_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_11_6_5 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uart_drone.bit_Count_2_LC_11_6_5  (
            .in0(N__33945),
            .in1(N__33936),
            .in2(N__35571),
            .in3(N__35484),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59079),
            .ce(),
            .sr(N__57500));
    defparam \uart_drone.bit_Count_0_LC_11_6_6 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_11_6_6 .LUT_INIT=16'b0000111101000000;
    LogicCell40 \uart_drone.bit_Count_0_LC_11_6_6  (
            .in0(N__35608),
            .in1(N__33918),
            .in2(N__33881),
            .in3(N__35409),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59079),
            .ce(),
            .sr(N__57500));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_11_6_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_11_6_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_11_6_7  (
            .in0(N__33860),
            .in1(N__35607),
            .in2(_gnd_net_),
            .in3(N__33798),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_11_7_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_11_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__33722),
            .in2(N__33705),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_11_7_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__33680),
            .in2(_gnd_net_),
            .in3(N__33663),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_11_7_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__33659),
            .in2(_gnd_net_),
            .in3(N__33648),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__59082),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_11_7_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_11_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__33645),
            .in2(_gnd_net_),
            .in3(N__33633),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__59082),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_11_7_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_11_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__34068),
            .in2(_gnd_net_),
            .in3(N__34056),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__59082),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_11_7_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_11_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__34052),
            .in2(_gnd_net_),
            .in3(N__34041),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__59082),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_11_7_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_11_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__34038),
            .in2(_gnd_net_),
            .in3(N__34026),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__59082),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_11_7_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_11_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__34023),
            .in2(_gnd_net_),
            .in3(N__34011),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__59082),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_11_8_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_11_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__34007),
            .in2(_gnd_net_),
            .in3(N__33993),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_11_8_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_11_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__34286),
            .in2(_gnd_net_),
            .in3(N__33990),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_11_8_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_11_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__34301),
            .in2(_gnd_net_),
            .in3(N__33987),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_11_8_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_11_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__33983),
            .in2(_gnd_net_),
            .in3(N__33972),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_11_8_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_11_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__34206),
            .in2(_gnd_net_),
            .in3(N__34137),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_11_8_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_11_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__34313),
            .in2(_gnd_net_),
            .in3(N__34134),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_11_8_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_11_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__34230),
            .in2(_gnd_net_),
            .in3(N__34131),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_11_8_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_11_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__34128),
            .in2(_gnd_net_),
            .in3(N__34116),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__59085),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_11_9_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_11_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__34274),
            .in2(_gnd_net_),
            .in3(N__34113),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__59090),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_11_9_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_11_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__34110),
            .in2(_gnd_net_),
            .in3(N__34098),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__59090),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_11_9_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_11_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__34239),
            .in2(_gnd_net_),
            .in3(N__34095),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__59090),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_11_9_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_11_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__34088),
            .in2(_gnd_net_),
            .in3(N__34074),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__59090),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_11_9_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_11_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__34217),
            .in2(_gnd_net_),
            .in3(N__34071),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59090),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_9_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_9_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_11_9_5  (
            .in0(N__35485),
            .in1(N__35559),
            .in2(_gnd_net_),
            .in3(N__35419),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNISRMR1_10_LC_11_9_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNISRMR1_10_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNISRMR1_10_LC_11_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNISRMR1_10_LC_11_9_6  (
            .in0(N__34314),
            .in1(N__34302),
            .in2(N__34290),
            .in3(N__34275),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_11_9_7 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_11_9_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_11_9_7  (
            .in0(N__34238),
            .in1(N__34229),
            .in2(N__34218),
            .in3(N__34205),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_0_LC_11_10_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_11_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__34173),
            .in2(N__34188),
            .in3(N__34187),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_1_LC_11_10_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_11_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__34167),
            .in2(_gnd_net_),
            .in3(N__34161),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_2_LC_11_10_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_11_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__34158),
            .in2(_gnd_net_),
            .in3(N__34152),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_3_LC_11_10_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_11_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__34149),
            .in2(_gnd_net_),
            .in3(N__34143),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_4_LC_11_10_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_11_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__34493),
            .in2(_gnd_net_),
            .in3(N__34140),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_5_LC_11_10_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_11_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__34541),
            .in2(_gnd_net_),
            .in3(N__34347),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_6_LC_11_10_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_11_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__34508),
            .in2(_gnd_net_),
            .in3(N__34344),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_7_LC_11_10_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_11_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__34526),
            .in2(_gnd_net_),
            .in3(N__34341),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__59096),
            .ce(),
            .sr(N__40875));
    defparam \dron_frame_decoder_1.WDT_8_LC_11_11_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_11_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__34407),
            .in2(_gnd_net_),
            .in3(N__34338),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_9_LC_11_11_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_11_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__34479),
            .in2(_gnd_net_),
            .in3(N__34335),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_10_LC_11_11_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_11_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__34442),
            .in2(_gnd_net_),
            .in3(N__34332),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_11_LC_11_11_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_11_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__34422),
            .in2(_gnd_net_),
            .in3(N__34329),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_12_LC_11_11_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_11_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__34394),
            .in2(_gnd_net_),
            .in3(N__34326),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_13_LC_11_11_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_11_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__34455),
            .in2(_gnd_net_),
            .in3(N__34323),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_14_LC_11_11_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_11_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__34581),
            .in2(_gnd_net_),
            .in3(N__34566),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_15_LC_11_11_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_11_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__34559),
            .in2(_gnd_net_),
            .in3(N__34563),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59104),
            .ce(),
            .sr(N__40871));
    defparam \dron_frame_decoder_1.WDT_RNIIVJ1_4_LC_11_12_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIIVJ1_4_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIIVJ1_4_LC_11_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIIVJ1_4_LC_11_12_0  (
            .in0(N__34542),
            .in1(N__34527),
            .in2(N__34512),
            .in3(N__34494),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT_RNIIVJ1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_9_LC_11_12_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_9_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_9_LC_11_12_1 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIATMH2_9_LC_11_12_1  (
            .in0(N__34478),
            .in1(N__34428),
            .in2(N__34467),
            .in3(N__34377),
            .lcout(\dron_frame_decoder_1.WDT10lt14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_11_12_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_11_12_2 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_11_12_2  (
            .in0(N__34454),
            .in1(N__34393),
            .in2(N__34443),
            .in3(N__34421),
            .lcout(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI2LQQ_8_LC_11_12_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI2LQQ_8_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI2LQQ_8_LC_11_12_3 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI2LQQ_8_LC_11_12_3  (
            .in0(N__34420),
            .in1(N__34406),
            .in2(N__34395),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.WDT10lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_11_12_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_11_12_7 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \dron_frame_decoder_1.state_RNITC181_2_LC_11_12_7  (
            .in0(N__36153),
            .in1(N__40974),
            .in2(N__34370),
            .in3(N__57841),
            .lcout(\dron_frame_decoder_1.N_481_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_5_LC_11_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_11_13_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_11_13_1  (
            .in0(N__34596),
            .in1(N__34632),
            .in2(N__45314),
            .in3(N__43216),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59120),
            .ce(),
            .sr(N__57528));
    defparam \dron_frame_decoder_1.state_2_LC_11_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_11_13_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_11_13_3  (
            .in0(N__36152),
            .in1(N__40983),
            .in2(N__34371),
            .in3(N__34691),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59120),
            .ce(),
            .sr(N__57528));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_11_14_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_11_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__36248),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_11_14_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__41435),
            .in2(N__42295),
            .in3(N__34644),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_11_14_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_11_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__37613),
            .in2(_gnd_net_),
            .in3(N__34641),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_11_14_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_11_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__36086),
            .in2(N__42296),
            .in3(N__34638),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_11_14_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_11_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__36020),
            .in2(_gnd_net_),
            .in3(N__34635),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_11_14_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_11_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__34631),
            .in2(_gnd_net_),
            .in3(N__34590),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_11_14_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_11_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__36125),
            .in2(N__42297),
            .in3(N__34587),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_11_14_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__36219),
            .in2(_gnd_net_),
            .in3(N__34584),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_11_15_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__35978),
            .in2(_gnd_net_),
            .in3(N__34785),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_11_15_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__36065),
            .in2(_gnd_net_),
            .in3(N__34782),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_11_15_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_11_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__34728),
            .in2(_gnd_net_),
            .in3(N__34779),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_11_15_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_11_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__40046),
            .in2(_gnd_net_),
            .in3(N__34776),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_11_15_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_11_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__35939),
            .in2(_gnd_net_),
            .in3(N__34773),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_11_15_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_11_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__42258),
            .in2(N__34764),
            .in3(N__34770),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_11_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_11_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34767),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59147),
            .ce(N__46762),
            .sr(N__57541));
    defparam \ppm_encoder_1.throttle_13_LC_11_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_11_16_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_11_16_0 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_11_16_0  (
            .in0(N__34760),
            .in1(N__34734),
            .in2(N__45387),
            .in3(N__37813),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59159),
            .ce(),
            .sr(N__57551));
    defparam \ppm_encoder_1.aileron_9_LC_11_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_11_16_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_11_16_4  (
            .in0(N__42849),
            .in1(N__34875),
            .in2(N__45386),
            .in3(N__39974),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59159),
            .ce(),
            .sr(N__57551));
    defparam \ppm_encoder_1.throttle_10_LC_11_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_11_16_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_11_16_5  (
            .in0(N__34727),
            .in1(N__34815),
            .in2(N__40552),
            .in3(N__45321),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59159),
            .ce(),
            .sr(N__57551));
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__43293),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__41547),
            .in2(N__42364),
            .in3(N__34809),
            .lcout(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_0 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_17_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__41124),
            .in2(_gnd_net_),
            .in3(N__34806),
            .lcout(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_1 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_17_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__43952),
            .in2(N__42365),
            .in3(N__34803),
            .lcout(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_2 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_17_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__43247),
            .in2(_gnd_net_),
            .in3(N__34800),
            .lcout(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_3 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_17_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__43275),
            .in2(_gnd_net_),
            .in3(N__34797),
            .lcout(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_4 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_17_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__42336),
            .in2(N__42974),
            .in3(N__34794),
            .lcout(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_5 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_17_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42929),
            .in3(N__34791),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_18_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__42884),
            .in2(_gnd_net_),
            .in3(N__34788),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_18_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__42848),
            .in2(_gnd_net_),
            .in3(N__34866),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_18_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__43044),
            .in2(_gnd_net_),
            .in3(N__34863),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_18_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__43011),
            .in2(_gnd_net_),
            .in3(N__34860),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_18_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__45597),
            .in2(_gnd_net_),
            .in3(N__34857),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_18_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__48066),
            .in2(N__42366),
            .in3(N__34854),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34851),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59190),
            .ce(N__46782),
            .sr(N__57571));
    defparam \pid_alt.error_axb_2_LC_11_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_11_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34836),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_11_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_2_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50383),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59200),
            .ce(N__34953),
            .sr(N__57576));
    defparam \pid_alt.error_axb_3_LC_11_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_11_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34959),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_11_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_11_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_3_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52683),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59200),
            .ce(N__34953),
            .sr(N__57576));
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_11_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_11_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34923),
            .lcout(\pid_alt.error_d_reg_prev_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_1_LC_11_19_5 .C_ON=1'b0;
    defparam \pid_front.error_axb_1_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_1_LC_11_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_1_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36255),
            .lcout(\pid_front.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIUJRT3_12_LC_11_20_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIUJRT3_12_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIUJRT3_12_LC_11_20_0 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIUJRT3_12_LC_11_20_0  (
            .in0(N__36957),
            .in1(N__37008),
            .in2(N__37146),
            .in3(N__35330),
            .lcout(\pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12 ),
            .ltout(\pid_front.pid_prereg_esr_RNIUJRT3Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI3F0N8_10_LC_11_20_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI3F0N8_10_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI3F0N8_10_LC_11_20_1 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI3F0N8_10_LC_11_20_1  (
            .in0(N__35297),
            .in1(N__35233),
            .in2(N__34884),
            .in3(_gnd_net_),
            .lcout(\pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10 ),
            .ltout(\pid_front.pid_prereg_esr_RNI3F0N8Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_1_LC_11_20_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_1_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_1_LC_11_20_2 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_front.source_pid_1_esr_1_LC_11_20_2  (
            .in0(N__50442),
            .in1(N__36725),
            .in2(N__34881),
            .in3(N__35065),
            .lcout(front_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59215),
            .ce(N__35209),
            .sr(N__35187));
    defparam \pid_front.source_pid_1_esr_2_LC_11_20_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_2_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_2_LC_11_20_3 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pid_front.source_pid_1_esr_2_LC_11_20_3  (
            .in0(N__35066),
            .in1(N__36726),
            .in2(N__36335),
            .in3(N__35053),
            .lcout(front_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59215),
            .ce(N__35209),
            .sr(N__35187));
    defparam \pid_front.pid_prereg_esr_RNIDT6R8_5_LC_11_20_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIDT6R8_5_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIDT6R8_5_LC_11_20_4 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIDT6R8_5_LC_11_20_4  (
            .in0(N__35234),
            .in1(N__35298),
            .in2(N__36686),
            .in3(N__35269),
            .lcout(\pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5 ),
            .ltout(\pid_front.pid_prereg_esr_RNIDT6R8Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_0_LC_11_20_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_0_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_0_LC_11_20_5 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \pid_front.source_pid_1_esr_0_LC_11_20_5  (
            .in0(N__36724),
            .in1(N__49431),
            .in2(N__34878),
            .in3(N__35052),
            .lcout(front_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59215),
            .ce(N__35209),
            .sr(N__35187));
    defparam \pid_front.source_pid_1_esr_4_LC_11_20_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_4_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_4_LC_11_20_6 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \pid_front.source_pid_1_esr_4_LC_11_20_6  (
            .in0(N__35055),
            .in1(N__36723),
            .in2(N__36687),
            .in3(N__35270),
            .lcout(front_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59215),
            .ce(N__35209),
            .sr(N__35187));
    defparam \pid_front.source_pid_1_esr_3_LC_11_20_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_3_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_3_LC_11_20_7 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pid_front.source_pid_1_esr_3_LC_11_20_7  (
            .in0(N__35067),
            .in1(N__36727),
            .in2(N__36776),
            .in3(N__35054),
            .lcout(front_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59215),
            .ce(N__35209),
            .sr(N__35187));
    defparam \pid_front.error_d_reg_esr_RNI7KE8_7_LC_11_21_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNI7KE8_7_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNI7KE8_7_LC_11_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_esr_RNI7KE8_7_LC_11_21_0  (
            .in0(N__35040),
            .in1(N__35119),
            .in2(_gnd_net_),
            .in3(N__59395),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_60_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI94TV_6_LC_11_21_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI94TV_6_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI94TV_6_LC_11_21_1 .LUT_INIT=16'b0100101101001011;
    LogicCell40 \pid_front.error_p_reg_esr_RNI94TV_6_LC_11_21_1  (
            .in0(N__35009),
            .in1(N__34979),
            .in2(N__35016),
            .in3(N__36606),
            .lcout(\pid_front.error_p_reg_esr_RNI94TVZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_6_LC_11_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_11_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_6_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52217),
            .lcout(\pid_front.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59232),
            .ce(N__49366),
            .sr(N__57596));
    defparam \pid_front.error_p_reg_esr_RNIG0G7_6_LC_11_21_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIG0G7_6_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIG0G7_6_LC_11_21_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIG0G7_6_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__35007),
            .in2(_gnd_net_),
            .in3(N__34977),
            .lcout(),
            .ltout(\pid_front.N_1447_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIIFUF_6_LC_11_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIIFUF_6_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIIFUF_6_LC_11_21_4 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \pid_front.error_d_reg_esr_RNIIFUF_6_LC_11_21_4  (
            .in0(N__52218),
            .in1(N__38049),
            .in2(N__35013),
            .in3(N__38304),
            .lcout(\pid_front.error_d_reg_esr_RNIIFUFZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNI4HE8_6_LC_11_21_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNI4HE8_6_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNI4HE8_6_LC_11_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_esr_RNI4HE8_6_LC_11_21_5  (
            .in0(N__52216),
            .in1(N__35008),
            .in2(_gnd_net_),
            .in3(N__34978),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_50_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH8R01_5_LC_11_21_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH8R01_5_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH8R01_5_LC_11_21_6 .LUT_INIT=16'b0011110000001111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH8R01_5_LC_11_21_6  (
            .in0(N__38013),
            .in1(N__38048),
            .in2(N__34962),
            .in3(N__38303),
            .lcout(\pid_front.error_p_reg_esr_RNIH8R01Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_7_LC_11_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_11_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_11_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_7_LC_11_21_7  (
            .in0(N__59396),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59232),
            .ce(N__49366),
            .sr(N__57596));
    defparam \pid_front.pid_prereg_esr_RNII3QG_6_LC_11_22_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNII3QG_6_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNII3QG_6_LC_11_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNII3QG_6_LC_11_22_0  (
            .in0(N__36524),
            .in1(N__36625),
            .in2(N__36580),
            .in3(N__36451),
            .lcout(\pid_front.m26_e_5 ),
            .ltout(\pid_front.m26_e_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIVDO51_10_LC_11_22_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIVDO51_10_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIVDO51_10_LC_11_22_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIVDO51_10_LC_11_22_1  (
            .in0(N__37055),
            .in1(_gnd_net_),
            .in2(N__35106),
            .in3(N__36371),
            .lcout(\pid_front.pid_prereg_esr_RNIVDO51Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIHEUK_12_LC_11_22_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIHEUK_12_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIHEUK_12_LC_11_22_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIHEUK_12_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__37002),
            .in2(_gnd_net_),
            .in3(N__36942),
            .lcout(),
            .ltout(\pid_front.m26_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIGSMQ1_10_LC_11_22_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIGSMQ1_10_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIGSMQ1_10_LC_11_22_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIGSMQ1_10_LC_11_22_3  (
            .in0(N__37053),
            .in1(N__36369),
            .in2(N__35103),
            .in3(N__35100),
            .lcout(\pid_front.pid_prereg_esr_RNIGSMQ1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIEUJ31_10_LC_11_22_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIEUJ31_10_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIEUJ31_10_LC_11_22_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIEUJ31_10_LC_11_22_4  (
            .in0(N__36370),
            .in1(N__37054),
            .in2(N__36731),
            .in3(N__37003),
            .lcout(\pid_front.m18_s_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNII3QG_0_6_LC_11_22_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNII3QG_0_6_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNII3QG_0_6_LC_11_22_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNII3QG_0_6_LC_11_22_5  (
            .in0(N__36514),
            .in1(N__36626),
            .in2(N__36581),
            .in3(N__36452),
            .lcout(\pid_front.m18_s_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_12_LC_11_22_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_12_LC_11_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_12_LC_11_22_6 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \pid_front.source_pid_1_esr_12_LC_11_22_6  (
            .in0(N__36949),
            .in1(N__37004),
            .in2(N__37139),
            .in3(N__35325),
            .lcout(front_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59250),
            .ce(N__35220),
            .sr(N__35188));
    defparam \pid_front.source_pid_1_esr_13_LC_11_22_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_13_LC_11_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_13_LC_11_22_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_13_LC_11_22_7  (
            .in0(N__35326),
            .in1(N__37124),
            .in2(_gnd_net_),
            .in3(N__36948),
            .lcout(front_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59250),
            .ce(N__35220),
            .sr(N__35188));
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_11_23_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_11_23_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIMHT91_16_LC_11_23_0  (
            .in0(N__36831),
            .in1(N__36801),
            .in2(N__37278),
            .in3(N__37245),
            .lcout(\pid_front.m9_e_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIEREV_14_LC_11_23_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIEREV_14_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIEREV_14_LC_11_23_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIEREV_14_LC_11_23_1  (
            .in0(N__36864),
            .in1(N__36900),
            .in2(_gnd_net_),
            .in3(N__37158),
            .lcout(),
            .ltout(\pid_front.m9_e_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIJRCU2_20_LC_11_23_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIJRCU2_20_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIJRCU2_20_LC_11_23_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIJRCU2_20_LC_11_23_2  (
            .in0(N__37179),
            .in1(N__37212),
            .in2(N__35340),
            .in3(N__35337),
            .lcout(\pid_front.pid_prereg_esr_RNIJRCU2Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_5_LC_11_23_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_5_LC_11_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_5_LC_11_23_3 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \pid_front.source_pid_1_esr_5_LC_11_23_3  (
            .in0(N__35296),
            .in1(N__35280),
            .in2(N__36685),
            .in3(N__35241),
            .lcout(front_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59265),
            .ce(N__35219),
            .sr(N__35193));
    defparam \pid_front.state_RNIVIRQ_0_LC_11_23_4 .C_ON=1'b0;
    defparam \pid_front.state_RNIVIRQ_0_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVIRQ_0_LC_11_23_4 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \pid_front.state_RNIVIRQ_0_LC_11_23_4  (
            .in0(N__50625),
            .in1(N__47709),
            .in2(N__50507),
            .in3(N__57835),
            .lcout(),
            .ltout(\pid_front.state_RNIVIRQZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNISV141_0_LC_11_23_5 .C_ON=1'b0;
    defparam \pid_front.state_RNISV141_0_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNISV141_0_LC_11_23_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_front.state_RNISV141_0_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35160),
            .in3(N__58320),
            .lcout(\pid_front.N_543_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNI9NAB3_10_LC_11_24_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNI9NAB3_10_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNI9NAB3_10_LC_11_24_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_d_reg_esr_RNI9NAB3_10_LC_11_24_0  (
            .in0(N__54314),
            .in1(N__35646),
            .in2(N__37082),
            .in3(N__35634),
            .lcout(\pid_front.error_d_reg_esr_RNI9NAB3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI653N_0_10_LC_11_24_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI653N_0_10_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI653N_0_10_LC_11_24_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_p_reg_esr_RNI653N_0_10_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__35153),
            .in2(_gnd_net_),
            .in3(N__35684),
            .lcout(\pid_front.N_1463_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI653N_10_LC_11_24_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI653N_10_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI653N_10_LC_11_24_4 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_front.error_p_reg_esr_RNI653N_10_LC_11_24_4  (
            .in0(N__35685),
            .in1(_gnd_net_),
            .in2(N__35157),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNI653NZ0Z_10 ),
            .ltout(\pid_front.error_p_reg_esr_RNI653NZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIESET1_0_10_LC_11_24_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIESET1_0_10_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIESET1_0_10_LC_11_24_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIESET1_0_10_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__35674),
            .in2(N__35133),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNIESET1_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_10_LC_11_24_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_11_24_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_10_LC_11_24_6  (
            .in0(N__54315),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59278),
            .ce(N__49362),
            .sr(N__57616));
    defparam \pid_front.error_p_reg_esr_RNIESET1_10_LC_11_24_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIESET1_10_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIESET1_10_LC_11_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIESET1_10_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__35675),
            .in2(_gnd_net_),
            .in3(N__35657),
            .lcout(\pid_front.error_p_reg_esr_RNIESET1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNISPQT1_10_LC_11_25_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNISPQT1_10_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNISPQT1_10_LC_11_25_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_esr_RNISPQT1_10_LC_11_25_7  (
            .in0(N__54308),
            .in1(N__35645),
            .in2(N__36420),
            .in3(N__35633),
            .lcout(\pid_front.error_d_reg_esr_RNISPQT1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_12_6_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_12_6_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_12_6_2  (
            .in0(N__35537),
            .in1(N__35464),
            .in2(_gnd_net_),
            .in3(N__35389),
            .lcout(\uart_drone.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIL5IF_0_LC_12_9_0 .C_ON=1'b0;
    defparam \pid_side.state_RNIL5IF_0_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIL5IF_0_LC_12_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNIL5IF_0_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__47621),
            .in2(_gnd_net_),
            .in3(N__57834),
            .lcout(\pid_side.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_12_9_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_12_9_1 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_12_9_1  (
            .in0(N__35564),
            .in1(N__35497),
            .in2(N__35426),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_12_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_12_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56479),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_12_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_12_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56284),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_12_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_12_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56124),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_12_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_12_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55353),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_12_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_12_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53379),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_12_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_12_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55903),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_12_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_12_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55733),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_12_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_12_11_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_12_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55567),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59097),
            .ce(N__35760),
            .sr(N__57525));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_12_12_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_12_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__41160),
            .in2(N__41206),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_12_12_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__35748),
            .in2(N__35742),
            .in3(N__35730),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_12_12_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__35727),
            .in2(N__35721),
            .in3(N__35709),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_12_12_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__35706),
            .in2(N__35700),
            .in3(N__35688),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_12_12_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__35901),
            .in2(N__35895),
            .in3(N__35880),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_12_12_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_12_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__35877),
            .in2(N__35871),
            .in3(N__35859),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_12_12_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_12_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__35856),
            .in2(N__35847),
            .in3(N__35838),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_12_12_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_12_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__35835),
            .in2(_gnd_net_),
            .in3(N__35820),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_12_13_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_12_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__35766),
            .in2(N__42298),
            .in3(N__35817),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_12_13_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_12_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35814),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_1849_i_l_ofx_LC_12_13_2 .C_ON=1'b0;
    defparam \scaler_4.N_1849_i_l_ofx_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_1849_i_l_ofx_LC_12_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_1849_i_l_ofx_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__35811),
            .in2(_gnd_net_),
            .in3(N__35783),
            .lcout(\scaler_4.N_1849_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_12_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_12_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__45203),
            .in2(_gnd_net_),
            .in3(N__57845),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_12_13_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_12_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI4N6K_2_LC_12_13_6  (
            .in0(N__40975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36148),
            .lcout(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_6_LC_12_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_12_14_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_12_14_2 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_12_14_2  (
            .in0(N__36132),
            .in1(N__36126),
            .in2(N__40171),
            .in3(N__45354),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59121),
            .ce(),
            .sr(N__57542));
    defparam \ppm_encoder_1.throttle_3_LC_12_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_12_14_3 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_12_14_3  (
            .in0(N__36096),
            .in1(N__36090),
            .in2(N__45398),
            .in3(N__44216),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59121),
            .ce(),
            .sr(N__57542));
    defparam \ppm_encoder_1.throttle_9_LC_12_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_12_15_1 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_12_15_1  (
            .in0(N__36066),
            .in1(N__45344),
            .in2(N__40251),
            .in3(N__36036),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59133),
            .ce(),
            .sr(N__57552));
    defparam \ppm_encoder_1.aileron_4_LC_12_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_4_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_4_LC_12_15_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_4_LC_12_15_4  (
            .in0(N__36030),
            .in1(N__43248),
            .in2(N__45396),
            .in3(N__46951),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59133),
            .ce(),
            .sr(N__57552));
    defparam \ppm_encoder_1.throttle_4_LC_12_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_12_15_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_12_15_5  (
            .in0(N__41872),
            .in1(N__45343),
            .in2(N__36021),
            .in3(N__35985),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59133),
            .ce(),
            .sr(N__57552));
    defparam \ppm_encoder_1.throttle_8_LC_12_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_12_15_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_12_15_6  (
            .in0(N__35979),
            .in1(N__35949),
            .in2(N__45397),
            .in3(N__40469),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59133),
            .ce(),
            .sr(N__57552));
    defparam \ppm_encoder_1.throttle_12_LC_12_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_12_15_7 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_12_15_7  (
            .in0(N__35943),
            .in1(N__45342),
            .in2(N__39952),
            .in3(N__35916),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59133),
            .ce(),
            .sr(N__57552));
    defparam \ppm_encoder_1.aileron_2_LC_12_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_2_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_2_LC_12_16_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_2_LC_12_16_0  (
            .in0(N__35910),
            .in1(N__41123),
            .in2(N__43792),
            .in3(N__45340),
            .lcout(\ppm_encoder_1.aileronZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59148),
            .ce(),
            .sr(N__57561));
    defparam \ppm_encoder_1.throttle_0_LC_12_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_12_16_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_12_16_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_12_16_1  (
            .in0(N__45333),
            .in1(N__36249),
            .in2(_gnd_net_),
            .in3(N__43660),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59148),
            .ce(),
            .sr(N__57561));
    defparam \ppm_encoder_1.throttle_7_LC_12_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_12_16_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_12_16_3  (
            .in0(N__36228),
            .in1(N__36214),
            .in2(N__45395),
            .in3(N__40342),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59148),
            .ce(),
            .sr(N__57561));
    defparam \ppm_encoder_1.elevator_10_LC_12_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_12_16_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_12_16_5  (
            .in0(N__37917),
            .in1(N__37884),
            .in2(N__45394),
            .in3(N__40520),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59148),
            .ce(),
            .sr(N__57561));
    defparam \ppm_encoder_1.elevator_2_LC_12_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_2_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_2_LC_12_16_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_2_LC_12_16_6  (
            .in0(N__37791),
            .in1(N__37773),
            .in2(N__47032),
            .in3(N__45341),
            .lcout(\ppm_encoder_1.elevatorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59148),
            .ce(),
            .sr(N__57561));
    defparam \ppm_encoder_1.elevator_8_LC_12_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_12_17_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_12_17_0  (
            .in0(N__37995),
            .in1(N__37968),
            .in2(N__45388),
            .in3(N__40455),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59160),
            .ce(),
            .sr(N__57572));
    defparam \ppm_encoder_1.aileron_10_LC_12_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_12_17_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_12_17_1  (
            .in0(N__43043),
            .in1(N__36186),
            .in2(N__45399),
            .in3(N__40496),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59160),
            .ce(),
            .sr(N__57572));
    defparam \ppm_encoder_1.aileron_13_LC_12_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_12_17_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_12_17_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_12_17_6  (
            .in0(N__48062),
            .in1(N__36180),
            .in2(N__38175),
            .in3(N__45358),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59160),
            .ce(),
            .sr(N__57572));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_12_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_12_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_12_18_1  (
            .in0(N__47163),
            .in1(N__37821),
            .in2(_gnd_net_),
            .in3(N__38124),
            .lcout(\ppm_encoder_1.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_12_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_12_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNI14DT_2_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__36170),
            .in2(_gnd_net_),
            .in3(N__57865),
            .lcout(\dron_frame_decoder_1.N_489_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICVO11_2_LC_12_19_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICVO11_2_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICVO11_2_LC_12_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNICVO11_2_LC_12_19_0  (
            .in0(N__36291),
            .in1(N__38246),
            .in2(N__36282),
            .in3(N__38230),
            .lcout(\pid_front.error_p_reg_esr_RNICVO11Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_19_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_19_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_19_1  (
            .in0(N__36311),
            .in1(N__36263),
            .in2(_gnd_net_),
            .in3(N__50866),
            .lcout(\pid_front.un1_pid_prereg_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_19_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_19_2 .LUT_INIT=16'b0110100101101001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_19_2  (
            .in0(N__50867),
            .in1(N__36312),
            .in2(N__36267),
            .in3(_gnd_net_),
            .lcout(\pid_front.un1_pid_prereg_2 ),
            .ltout(\pid_front.un1_pid_prereg_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJCSG_2_LC_12_19_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJCSG_2_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJCSG_2_LC_12_19_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJCSG_2_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36294),
            .in3(N__36290),
            .lcout(\pid_front.error_p_reg_esr_RNIJCSGZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_19_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_19_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_19_4  (
            .in0(N__38103),
            .in1(N__38082),
            .in2(_gnd_net_),
            .in3(N__49301),
            .lcout(\pid_front.un1_pid_prereg_0 ),
            .ltout(\pid_front.un1_pid_prereg_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH7Q01_1_LC_12_19_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH7Q01_1_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH7Q01_1_LC_12_19_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH7Q01_1_LC_12_19_5  (
            .in0(N__38568),
            .in1(N__36278),
            .in2(N__36270),
            .in3(N__38551),
            .lcout(\pid_front.error_p_reg_esr_RNIH7Q01Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_19_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_19_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_3_LC_12_19_6  (
            .in0(N__50868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59191),
            .ce(N__49372),
            .sr(N__57583));
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_19_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_2_LC_12_19_7  (
            .in0(N__49302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59191),
            .ce(N__49372),
            .sr(N__57583));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_12_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_12_20_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_12_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52291),
            .lcout(drone_H_disp_front_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50779),
            .lcout(drone_H_disp_front_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50398),
            .lcout(drone_H_disp_front_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52693),
            .lcout(drone_H_disp_front_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_20_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52598),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_12_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_12_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52477),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_12_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_12_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53211),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_12_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_12_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52391),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59201),
            .ce(N__36354),
            .sr(N__57597));
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_21_0 .C_ON=1'b1;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_0_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__49460),
            .in2(N__56939),
            .in3(N__56935),
            .lcout(\pid_front.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\pid_front.un1_pid_prereg_cry_0 ),
            .clk(N__59216),
            .ce(N__49369),
            .sr(N__57603));
    defparam \pid_front.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_12_21_1 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_12_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__50519),
            .in2(_gnd_net_),
            .in3(N__36339),
            .lcout(\pid_front.un1_pid_prereg_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_0 ),
            .carryout(\pid_front.un1_pid_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_2_LC_12_21_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_2_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_2_LC_12_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_2_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__38208),
            .in2(N__38589),
            .in3(N__36315),
            .lcout(\pid_front.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_1 ),
            .carryout(\pid_front.un1_pid_prereg_cry_0_0 ),
            .clk(N__59216),
            .ce(N__49369),
            .sr(N__57603));
    defparam \pid_front.pid_prereg_esr_3_LC_12_21_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_3_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_3_LC_12_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_3_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__38535),
            .in2(N__36792),
            .in3(N__36756),
            .lcout(\pid_front.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_0_0 ),
            .carryout(\pid_front.un1_pid_prereg_cry_1_0 ),
            .clk(N__59216),
            .ce(N__49369),
            .sr(N__57603));
    defparam \pid_front.pid_prereg_esr_4_LC_12_21_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_4_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_4_LC_12_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_4_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__36753),
            .in2(N__36744),
            .in3(N__36690),
            .lcout(\pid_front.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_1_0 ),
            .carryout(\pid_front.un1_pid_prereg_cry_2 ),
            .clk(N__59216),
            .ce(N__49369),
            .sr(N__57603));
    defparam \pid_front.pid_prereg_esr_5_LC_12_21_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_5_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_5_LC_12_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_5_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__38217),
            .in2(N__38070),
            .in3(N__36645),
            .lcout(\pid_front.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_2 ),
            .carryout(\pid_front.un1_pid_prereg_cry_3 ),
            .clk(N__59216),
            .ce(N__49369),
            .sr(N__57603));
    defparam \pid_front.pid_prereg_esr_6_LC_12_21_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_6_LC_12_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_6_LC_12_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_6_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__38006),
            .in2(N__36642),
            .in3(N__36609),
            .lcout(\pid_front.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_3 ),
            .carryout(\pid_front.un1_pid_prereg_cry_4 ),
            .clk(N__59216),
            .ce(N__49369),
            .sr(N__57603));
    defparam \pid_front.pid_prereg_esr_7_LC_12_21_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_7_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_7_LC_12_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_7_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__36605),
            .in2(N__36594),
            .in3(N__36555),
            .lcout(\pid_front.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_4 ),
            .carryout(\pid_front.un1_pid_prereg_cry_5 ),
            .clk(N__59216),
            .ce(N__49369),
            .sr(N__57603));
    defparam \pid_front.pid_prereg_esr_8_LC_12_22_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_8_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_8_LC_12_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_8_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__36552),
            .in2(N__36540),
            .in3(N__36495),
            .lcout(\pid_front.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\pid_front.un1_pid_prereg_cry_6 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_9_LC_12_22_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_9_LC_12_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_9_LC_12_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_9_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__36492),
            .in2(N__36474),
            .in3(N__36435),
            .lcout(\pid_front.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_6 ),
            .carryout(\pid_front.un1_pid_prereg_cry_7 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_10_LC_12_22_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_10_LC_12_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_10_LC_12_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_10_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__36432),
            .in2(N__36419),
            .in3(N__37095),
            .lcout(\pid_front.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_7 ),
            .carryout(\pid_front.un1_pid_prereg_cry_8 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_11_LC_12_22_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_11_LC_12_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_11_LC_12_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_11_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__37092),
            .in2(N__37083),
            .in3(N__37038),
            .lcout(\pid_front.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_8 ),
            .carryout(\pid_front.un1_pid_prereg_cry_9 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_12_LC_12_22_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_12_LC_12_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_12_LC_12_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_12_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__37035),
            .in2(N__37023),
            .in3(N__36987),
            .lcout(\pid_front.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_9 ),
            .carryout(\pid_front.un1_pid_prereg_cry_10 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_13_LC_12_22_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_13_LC_12_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_13_LC_12_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_13_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__36984),
            .in2(N__36969),
            .in3(N__36924),
            .lcout(\pid_front.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_10 ),
            .carryout(\pid_front.un1_pid_prereg_cry_11 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_14_LC_12_22_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_14_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_14_LC_12_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_14_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(N__36921),
            .in2(N__36912),
            .in3(N__36894),
            .lcout(\pid_front.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_11 ),
            .carryout(\pid_front.un1_pid_prereg_cry_12 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_15_LC_12_22_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_15_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_15_LC_12_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_15_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(N__36891),
            .in2(N__36879),
            .in3(N__36858),
            .lcout(\pid_front.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_12 ),
            .carryout(\pid_front.un1_pid_prereg_cry_13 ),
            .clk(N__59233),
            .ce(N__49367),
            .sr(N__57610));
    defparam \pid_front.pid_prereg_esr_16_LC_12_23_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_16_LC_12_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_16_LC_12_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_16_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__36855),
            .in2(N__36846),
            .in3(N__36825),
            .lcout(\pid_front.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(bfn_12_23_0_),
            .carryout(\pid_front.un1_pid_prereg_cry_14 ),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \pid_front.pid_prereg_esr_17_LC_12_23_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_17_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_17_LC_12_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_17_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__36822),
            .in2(N__36813),
            .in3(N__36795),
            .lcout(\pid_front.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_14 ),
            .carryout(\pid_front.un1_pid_prereg_cry_15 ),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \pid_front.pid_prereg_esr_18_LC_12_23_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_18_LC_12_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_18_LC_12_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_18_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__37299),
            .in2(N__37290),
            .in3(N__37269),
            .lcout(\pid_front.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_15 ),
            .carryout(\pid_front.un1_pid_prereg_cry_16 ),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \pid_front.pid_prereg_esr_19_LC_12_23_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_19_LC_12_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_19_LC_12_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_19_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__37266),
            .in2(N__37257),
            .in3(N__37239),
            .lcout(\pid_front.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_16 ),
            .carryout(\pid_front.un1_pid_prereg_cry_17 ),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \pid_front.pid_prereg_esr_20_LC_12_23_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_20_LC_12_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_20_LC_12_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_20_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__37236),
            .in2(N__37227),
            .in3(N__37206),
            .lcout(\pid_front.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_17 ),
            .carryout(\pid_front.un1_pid_prereg_cry_18 ),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \pid_front.pid_prereg_esr_21_LC_12_23_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_21_LC_12_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_21_LC_12_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_21_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__37203),
            .in2(N__37194),
            .in3(N__37173),
            .lcout(\pid_front.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_18 ),
            .carryout(\pid_front.un1_pid_prereg_cry_19 ),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \pid_front.pid_prereg_esr_22_LC_12_23_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_22_LC_12_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_22_LC_12_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_22_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__37170),
            .in2(N__42516),
            .in3(N__37152),
            .lcout(\pid_front.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_19 ),
            .carryout(\pid_front.un1_pid_prereg_cry_20 ),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \pid_front.pid_prereg_esr_23_LC_12_23_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_23_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_23_LC_12_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.pid_prereg_esr_23_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__37320),
            .in2(_gnd_net_),
            .in3(N__37149),
            .lcout(\pid_front.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59251),
            .ce(N__49365),
            .sr(N__57617));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_24_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_24_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56506),
            .lcout(front_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_24_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56311),
            .lcout(front_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_24_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_24_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56142),
            .lcout(front_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_24_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_24_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_12_24_3  (
            .in0(N__55356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(front_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_24_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53409),
            .lcout(front_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_24_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55932),
            .lcout(front_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_24_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_24_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55755),
            .lcout(front_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_24_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_24_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_12_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55584),
            .lcout(front_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59266),
            .ce(N__37338),
            .sr(N__57624));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_25_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39417),
            .lcout(drone_H_disp_front_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNO_0_23_LC_12_25_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNO_0_23_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNO_0_23_LC_12_25_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_front.pid_prereg_esr_RNO_0_23_LC_12_25_1  (
            .in0(N__42539),
            .in1(N__42609),
            .in2(N__42552),
            .in3(N__42610),
            .lcout(\pid_front.un1_pid_prereg_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_8_l_ofx_LC_12_25_2 .C_ON=1'b0;
    defparam \pid_front.error_axb_8_l_ofx_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_8_l_ofx_LC_12_25_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_front.error_axb_8_l_ofx_LC_12_25_2  (
            .in0(N__39411),
            .in1(_gnd_net_),
            .in2(N__37311),
            .in3(N__39398),
            .lcout(\pid_front.error_axb_8_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_7_LC_12_25_3 .C_ON=1'b0;
    defparam \pid_front.error_axb_7_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_7_LC_12_25_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_axb_7_LC_12_25_3  (
            .in0(_gnd_net_),
            .in1(N__37307),
            .in2(_gnd_net_),
            .in3(N__39410),
            .lcout(\pid_front.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_25_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39397),
            .lcout(drone_H_disp_front_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_12_25_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_12_25_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_12_25_6  (
            .in0(N__59501),
            .in1(_gnd_net_),
            .in2(N__43059),
            .in3(N__37362),
            .lcout(\pid_front.un1_pid_prereg_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_12_25_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_12_25_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8QE61_20_LC_12_25_7  (
            .in0(N__37361),
            .in1(N__43055),
            .in2(_gnd_net_),
            .in3(N__59500),
            .lcout(\pid_front.un1_pid_prereg_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIFCSD1_0_LC_13_8_0 .C_ON=1'b0;
    defparam \pid_alt.state_RNIFCSD1_0_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIFCSD1_0_LC_13_8_0 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_alt.state_RNIFCSD1_0_LC_13_8_0  (
            .in0(N__47684),
            .in1(N__39717),
            .in2(N__39595),
            .in3(N__57828),
            .lcout(\pid_alt.state_RNIFCSD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_LC_13_9_0 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_esr_LC_13_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_data_valid_esr_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39718),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59080),
            .ce(N__39840),
            .sr(N__57519));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__37595),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__37427),
            .in2(_gnd_net_),
            .in3(N__37347),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_10_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__39800),
            .in2(_gnd_net_),
            .in3(N__37344),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_10_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__39830),
            .in2(_gnd_net_),
            .in3(N__37341),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_10_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__39782),
            .in2(_gnd_net_),
            .in3(N__37410),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_10_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39552),
            .in3(N__37407),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_10_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__39528),
            .in2(_gnd_net_),
            .in3(N__37404),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_10_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__39761),
            .in2(N__42315),
            .in3(N__37401),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_13_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_13_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__37476),
            .in2(_gnd_net_),
            .in3(N__37398),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59088),
            .ce(N__46776),
            .sr(N__57529));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_13_12_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_13_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__41235),
            .in2(N__41139),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_13_12_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__37388),
            .in2(N__41245),
            .in3(N__37395),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__59094),
            .ce(N__37466),
            .sr(N__57535));
    defparam \scaler_4.source_data_1_esr_7_LC_13_12_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__37373),
            .in2(N__37392),
            .in3(N__37380),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__59094),
            .ce(N__37466),
            .sr(N__57535));
    defparam \scaler_4.source_data_1_esr_8_LC_13_12_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__37559),
            .in2(N__37377),
            .in3(N__37365),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__59094),
            .ce(N__37466),
            .sr(N__57535));
    defparam \scaler_4.source_data_1_esr_9_LC_13_12_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__37544),
            .in2(N__37563),
            .in3(N__37551),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__59094),
            .ce(N__37466),
            .sr(N__57535));
    defparam \scaler_4.source_data_1_esr_10_LC_13_12_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_13_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__37529),
            .in2(N__37548),
            .in3(N__37536),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__59094),
            .ce(N__37466),
            .sr(N__57535));
    defparam \scaler_4.source_data_1_esr_11_LC_13_12_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_13_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__37514),
            .in2(N__37533),
            .in3(N__37521),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__59094),
            .ce(N__37466),
            .sr(N__57535));
    defparam \scaler_4.source_data_1_esr_12_LC_13_12_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_13_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__37502),
            .in2(N__37518),
            .in3(N__37506),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__59094),
            .ce(N__37466),
            .sr(N__57535));
    defparam \scaler_4.source_data_1_esr_13_LC_13_13_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_13_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__37503),
            .in2(N__37491),
            .in3(N__37482),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__59102),
            .ce(N__37467),
            .sr(N__57543));
    defparam \scaler_4.source_data_1_esr_14_LC_13_13_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_13_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37479),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59102),
            .ce(N__37467),
            .sr(N__57543));
    defparam \ppm_encoder_1.rudder_7_LC_13_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_13_14_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_13_14_0  (
            .in0(N__37437),
            .in1(N__37428),
            .in2(N__45370),
            .in3(N__40576),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59111),
            .ce(),
            .sr(N__57553));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_13_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_13_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__43629),
            .in2(_gnd_net_),
            .in3(N__43538),
            .lcout(),
            .ltout(\ppm_encoder_1.N_134_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_14_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_14_2 .LUT_INIT=16'b1100110011110100;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_13_14_2  (
            .in0(N__43590),
            .in1(N__37634),
            .in2(N__37644),
            .in3(N__42654),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59111),
            .ce(),
            .sr(N__57553));
    defparam \ppm_encoder_1.throttle_2_LC_13_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_13_14_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_13_14_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_13_14_6  (
            .in0(N__37623),
            .in1(N__37614),
            .in2(N__45371),
            .in3(N__46993),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59111),
            .ce(),
            .sr(N__57553));
    defparam \ppm_encoder_1.elevator_4_LC_13_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_4_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_4_LC_13_15_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_4_LC_13_15_0  (
            .in0(N__37737),
            .in1(N__37761),
            .in2(N__45297),
            .in3(N__41852),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \ppm_encoder_1.elevator_5_LC_13_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_5_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_5_LC_13_15_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_5_LC_13_15_1  (
            .in0(N__37728),
            .in1(N__37698),
            .in2(N__43199),
            .in3(N__45200),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \ppm_encoder_1.elevator_9_LC_13_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_13_15_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_13_15_2  (
            .in0(N__37929),
            .in1(N__37959),
            .in2(N__45298),
            .in3(N__40227),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \ppm_encoder_1.rudder_6_LC_13_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_13_15_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_13_15_3 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_13_15_3  (
            .in0(N__37596),
            .in1(N__45190),
            .in2(_gnd_net_),
            .in3(N__40610),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \ppm_encoder_1.elevator_11_LC_13_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_13_15_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_13_15_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_13_15_4  (
            .in0(N__37875),
            .in1(N__37842),
            .in2(N__45296),
            .in3(N__40099),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \ppm_encoder_1.aileron_5_LC_13_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_5_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_5_LC_13_15_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_5_LC_13_15_5  (
            .in0(N__43274),
            .in1(N__37578),
            .in2(N__45295),
            .in3(N__51269),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \pid_alt.state_1_LC_13_15_6 .C_ON=1'b0;
    defparam \pid_alt.state_1_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_1_LC_13_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.state_1_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39599),
            .lcout(\pid_alt.N_72_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \ppm_encoder_1.elevator_6_LC_13_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_13_15_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_13_15_7 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_13_15_7  (
            .in0(N__45186),
            .in1(N__37689),
            .in2(N__40149),
            .in3(N__37656),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59118),
            .ce(),
            .sr(N__57562));
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_16_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__45428),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_16_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__41480),
            .in2(N__42316),
            .in3(N__37794),
            .lcout(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_0 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_16_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__37790),
            .in2(_gnd_net_),
            .in3(N__37767),
            .lcout(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_1 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_16_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__43886),
            .in2(N__42317),
            .in3(N__37764),
            .lcout(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_2 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_16_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(N__37760),
            .in2(_gnd_net_),
            .in3(N__37731),
            .lcout(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_3 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_16_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(N__37727),
            .in2(_gnd_net_),
            .in3(N__37692),
            .lcout(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_4 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_16_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__42278),
            .in2(N__37688),
            .in3(N__37650),
            .lcout(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_5 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_16_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(N__40292),
            .in2(_gnd_net_),
            .in3(N__37647),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__37994),
            .in2(_gnd_net_),
            .in3(N__37962),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__37955),
            .in2(_gnd_net_),
            .in3(N__37920),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_17_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__37916),
            .in2(_gnd_net_),
            .in3(N__37878),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_17_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__37874),
            .in2(_gnd_net_),
            .in3(N__37833),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_17_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__39890),
            .in2(_gnd_net_),
            .in3(N__37830),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_17_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__38153),
            .in2(N__42352),
            .in3(N__37827),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37824),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59145),
            .ce(N__46777),
            .sr(N__57577));
    defparam \ppm_encoder_1.throttle_RNIM4PT2_13_LC_13_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIM4PT2_13_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIM4PT2_13_LC_13_18_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIM4PT2_13_LC_13_18_0  (
            .in0(N__44372),
            .in1(N__37820),
            .in2(N__41361),
            .in3(N__44069),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIMC2D6_13_LC_13_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIMC2D6_13_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIMC2D6_13_LC_13_18_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIMC2D6_13_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__44400),
            .in2(N__37797),
            .in3(N__38187),
            .lcout(\ppm_encoder_1.elevator_RNIMC2D6Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_13_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_13_18_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNI68LH2_13_LC_13_18_2  (
            .in0(N__38122),
            .in1(N__38170),
            .in2(N__44202),
            .in3(N__45553),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_18_4  (
            .in0(N__51431),
            .in1(N__38181),
            .in2(_gnd_net_),
            .in3(N__38171),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_13_LC_13_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_13_18_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_13_18_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_13_18_6  (
            .in0(N__38123),
            .in1(N__38157),
            .in2(N__45401),
            .in3(N__38130),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59157),
            .ce(),
            .sr(N__57584));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38109),
            .lcout(drone_H_disp_front_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_13_19_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_13_19_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_13_19_7  (
            .in0(N__38102),
            .in1(N__38081),
            .in2(_gnd_net_),
            .in3(N__49295),
            .lcout(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIOBP11_5_LC_13_20_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIOBP11_5_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIOBP11_5_LC_13_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_esr_RNIOBP11_5_LC_13_20_0  (
            .in0(N__38232),
            .in1(N__38061),
            .in2(N__38250),
            .in3(N__38055),
            .lcout(\pid_front.error_d_reg_esr_RNIOBP11Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNI1EE8_5_LC_13_20_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNI1EE8_5_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNI1EE8_5_LC_13_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_esr_RNI1EE8_5_LC_13_20_1  (
            .in0(N__38046),
            .in1(N__38293),
            .in2(_gnd_net_),
            .in3(N__53080),
            .lcout(\pid_front.un1_pid_prereg_40_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_13_20_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_13_20_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_4_LC_13_20_2  (
            .in0(N__38279),
            .in1(N__38258),
            .in2(_gnd_net_),
            .in3(N__59425),
            .lcout(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ),
            .ltout(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIVOSG_5_LC_13_20_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIVOSG_5_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIVOSG_5_LC_13_20_3 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \pid_front.error_d_reg_esr_RNIVOSG_5_LC_13_20_3  (
            .in0(N__38047),
            .in1(N__38294),
            .in2(N__38016),
            .in3(N__53081),
            .lcout(\pid_front.error_d_reg_esr_RNIVOSGZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_5_LC_13_20_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_13_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_13_20_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_5_LC_13_20_4  (
            .in0(N__53082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59188),
            .ce(N__49373),
            .sr(N__57604));
    defparam \pid_front.error_d_reg_prev_esr_4_LC_13_20_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_13_20_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_4_LC_13_20_5  (
            .in0(N__59427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59188),
            .ce(N__49373),
            .sr(N__57604));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_13_20_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_13_20_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_13_20_6  (
            .in0(N__38280),
            .in1(N__38259),
            .in2(_gnd_net_),
            .in3(N__59426),
            .lcout(\pid_front.un1_pid_prereg_17 ),
            .ltout(\pid_front.un1_pid_prereg_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIPISG_3_LC_13_20_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIPISG_3_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIPISG_3_LC_13_20_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIPISG_3_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38235),
            .in3(N__38231),
            .lcout(\pid_front.error_p_reg_esr_RNIPISGZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6MF7_0_1_LC_13_21_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6MF7_0_1_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6MF7_0_1_LC_13_21_0 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6MF7_0_1_LC_13_21_0  (
            .in0(N__46919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38201),
            .lcout(\pid_front.N_1427_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI4KF7_0_LC_13_21_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI4KF7_0_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI4KF7_0_LC_13_21_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \pid_front.error_p_reg_esr_RNI4KF7_0_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__38396),
            .in2(_gnd_net_),
            .in3(N__38348),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNI4KF7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNINGRV_1_LC_13_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNINGRV_1_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNINGRV_1_LC_13_21_2 .LUT_INIT=16'b1100000011111100;
    LogicCell40 \pid_front.error_d_reg_esr_RNINGRV_1_LC_13_21_2  (
            .in0(N__38588),
            .in1(N__56894),
            .in2(N__38211),
            .in3(N__38325),
            .lcout(\pid_front.error_d_reg_esr_RNINGRVZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_13_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_13_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40721),
            .lcout(drone_H_disp_front_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6MF7_1_LC_13_21_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6MF7_1_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6MF7_1_LC_13_21_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6MF7_1_LC_13_21_4  (
            .in0(N__46920),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38202),
            .lcout(\pid_front.error_p_reg_esr_RNI6MF7Z0Z_1 ),
            .ltout(\pid_front.error_p_reg_esr_RNI6MF7Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUQTF_0_1_LC_13_21_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUQTF_0_1_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUQTF_0_1_LC_13_21_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUQTF_0_1_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38592),
            .in3(N__38552),
            .lcout(\pid_front.un1_pid_prereg ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_3_LC_13_21_6 .C_ON=1'b0;
    defparam \pid_front.error_axb_3_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_3_LC_13_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_3_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38574),
            .lcout(\pid_front.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUQTF_1_LC_13_21_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUQTF_1_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUQTF_1_LC_13_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUQTF_1_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__38564),
            .in2(_gnd_net_),
            .in3(N__38553),
            .lcout(\pid_front.error_p_reg_esr_RNIUQTFZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_13_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_13_22_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_13_22_1  (
            .in0(N__38528),
            .in1(N__38490),
            .in2(_gnd_net_),
            .in3(N__38457),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_22_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38415),
            .lcout(drone_H_disp_front_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_22_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38406),
            .lcout(drone_H_disp_front_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_RNIPLTF_1_LC_13_22_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_RNIPLTF_1_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_esr_RNIPLTF_1_LC_13_22_4 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \pid_front.error_d_reg_esr_RNIPLTF_1_LC_13_22_4  (
            .in0(N__38397),
            .in1(N__38347),
            .in2(N__56893),
            .in3(N__38324),
            .lcout(\pid_front.un1_pid_prereg_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_22_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38313),
            .lcout(drone_H_disp_front_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_2_LC_13_22_6 .C_ON=1'b0;
    defparam \pid_front.error_axb_2_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_2_LC_13_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_2_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38925),
            .lcout(\pid_front.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_22_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39360),
            .lcout(drone_H_disp_front_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_inv_LC_13_23_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_inv_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_inv_LC_13_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_cry_0_c_inv_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__38871),
            .in2(_gnd_net_),
            .in3(N__38902),
            .lcout(\pid_front.error_axb_0 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\pid_front.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_13_23_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_13_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_0_c_RNIC7KB_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__38865),
            .in2(_gnd_net_),
            .in3(N__38811),
            .lcout(\pid_front.error_1 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0 ),
            .carryout(\pid_front.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_13_23_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_13_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_1_c_RNIEALB_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__38808),
            .in2(_gnd_net_),
            .in3(N__38763),
            .lcout(\pid_front.error_2 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1 ),
            .carryout(\pid_front.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_13_23_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_13_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_2_c_RNIGDMB_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__38760),
            .in2(_gnd_net_),
            .in3(N__38712),
            .lcout(\pid_front.error_3 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2 ),
            .carryout(\pid_front.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_13_23_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_13_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_c_RNIABAG_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__38709),
            .in2(N__38703),
            .in3(N__38652),
            .lcout(\pid_front.error_4 ),
            .ltout(),
            .carryin(\pid_front.error_cry_3 ),
            .carryout(\pid_front.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_23_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__38649),
            .in2(N__38643),
            .in3(N__38595),
            .lcout(\pid_front.error_5 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0_0 ),
            .carryout(\pid_front.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_23_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__39342),
            .in2(N__39336),
            .in3(N__39294),
            .lcout(\pid_front.error_6 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1_0 ),
            .carryout(\pid_front.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_13_23_7 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_13_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIU61K_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__39291),
            .in2(N__39279),
            .in3(N__39231),
            .lcout(\pid_front.error_7 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2_0 ),
            .carryout(\pid_front.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_24_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__39228),
            .in2(N__39219),
            .in3(N__39171),
            .lcout(\pid_front.error_8 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\pid_front.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_13_24_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_13_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_4_c_RNILNBG_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__50799),
            .in2(N__39168),
            .in3(N__39120),
            .lcout(\pid_front.error_9 ),
            .ltout(),
            .carryin(\pid_front.error_cry_4 ),
            .carryout(\pid_front.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_13_24_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_13_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_5_c_RNIVNFF_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__39117),
            .in2(N__39111),
            .in3(N__39060),
            .lcout(\pid_front.error_10 ),
            .ltout(),
            .carryin(\pid_front.error_cry_5 ),
            .carryout(\pid_front.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_13_24_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_13_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_6_c_RNI3VJG_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__39057),
            .in2(_gnd_net_),
            .in3(N__39012),
            .lcout(\pid_front.error_11 ),
            .ltout(),
            .carryin(\pid_front.error_cry_6 ),
            .carryout(\pid_front.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_13_24_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_13_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_7_c_RNIAPPM_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__39009),
            .in2(N__39402),
            .in3(N__38970),
            .lcout(\pid_front.error_12 ),
            .ltout(),
            .carryin(\pid_front.error_cry_7 ),
            .carryout(\pid_front.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_13_24_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_13_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_8_c_RNIAC2E_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__38967),
            .in2(N__40731),
            .in3(N__38928),
            .lcout(\pid_front.error_13 ),
            .ltout(),
            .carryin(\pid_front.error_cry_8 ),
            .carryout(\pid_front.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_13_24_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_13_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_9_c_RNIDG3E_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__39507),
            .in2(N__39384),
            .in3(N__39459),
            .lcout(\pid_front.error_14 ),
            .ltout(),
            .carryin(\pid_front.error_cry_9 ),
            .carryout(\pid_front.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_13_24_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_13_24_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_cry_10_c_RNINTDI_LC_13_24_7  (
            .in0(N__39369),
            .in1(N__39383),
            .in2(_gnd_net_),
            .in3(N__39456),
            .lcout(\pid_front.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_13_25_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_13_25_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_13_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50403),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59263),
            .ce(N__50697),
            .sr(N__57636));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_25_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_25_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52708),
            .lcout(drone_H_disp_front_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59263),
            .ce(N__50697),
            .sr(N__57636));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_25_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_25_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52597),
            .lcout(drone_H_disp_front_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59263),
            .ce(N__50697),
            .sr(N__57636));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_13_25_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_13_25_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_13_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_13_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53228),
            .lcout(drone_H_disp_front_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59263),
            .ce(N__50697),
            .sr(N__57636));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_25_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_25_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52395),
            .lcout(drone_H_disp_front_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59263),
            .ce(N__50697),
            .sr(N__57636));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_25_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_25_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52300),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59263),
            .ce(N__50697),
            .sr(N__57636));
    defparam \pid_alt.state_RNIH1EN_0_LC_13_29_4 .C_ON=1'b0;
    defparam \pid_alt.state_RNIH1EN_0_LC_13_29_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIH1EN_0_LC_13_29_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIH1EN_0_LC_13_29_4  (
            .in0(_gnd_net_),
            .in1(N__39600),
            .in2(_gnd_net_),
            .in3(N__57836),
            .lcout(\pid_alt.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_RNO_LC_14_9_7 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_14_9_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_alt.source_data_valid_esr_RNO_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__39588),
            .in2(_gnd_net_),
            .in3(N__57870),
            .lcout(\pid_alt.state_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_9_LC_14_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_14_10_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_14_10_1  (
            .in0(N__39831),
            .in1(N__39813),
            .in2(N__45202),
            .in3(N__40204),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59091),
            .ce(),
            .sr(N__57530));
    defparam \ppm_encoder_1.rudder_8_LC_14_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_14_10_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_14_10_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_14_10_4  (
            .in0(N__39807),
            .in1(N__39801),
            .in2(N__46231),
            .in3(N__45132),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59091),
            .ce(),
            .sr(N__57530));
    defparam \ppm_encoder_1.rudder_10_LC_14_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_14_10_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_14_10_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_14_10_5  (
            .in0(N__39783),
            .in1(N__39768),
            .in2(N__45201),
            .in3(N__46291),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59091),
            .ce(),
            .sr(N__57530));
    defparam \ppm_encoder_1.rudder_13_LC_14_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_14_11_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_14_11_1 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_14_11_1  (
            .in0(N__39762),
            .in1(N__39744),
            .in2(N__45374),
            .in3(N__44365),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59098),
            .ce(),
            .sr(N__57536));
    defparam \pid_alt.state_0_LC_14_11_2 .C_ON=1'b0;
    defparam \pid_alt.state_0_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_0_LC_14_11_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_alt.state_0_LC_14_11_2  (
            .in0(N__39584),
            .in1(N__47705),
            .in2(_gnd_net_),
            .in3(N__39676),
            .lcout(\pid_alt.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59098),
            .ce(),
            .sr(N__57536));
    defparam \ppm_encoder_1.rudder_11_LC_14_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_14_11_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_14_11_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_14_11_3  (
            .in0(N__39551),
            .in1(N__39534),
            .in2(N__45372),
            .in3(N__40850),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59098),
            .ce(),
            .sr(N__57536));
    defparam \ppm_encoder_1.rudder_12_LC_14_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_14_11_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_14_11_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_14_11_5  (
            .in0(N__39527),
            .in1(N__39513),
            .in2(N__45373),
            .in3(N__46712),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59098),
            .ce(),
            .sr(N__57536));
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_12_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_12_0  (
            .in0(N__39859),
            .in1(N__39907),
            .in2(N__45558),
            .in3(N__44189),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_12_2  (
            .in0(N__39953),
            .in1(N__46708),
            .in2(N__41353),
            .in3(N__44053),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_12_3  (
            .in0(N__47178),
            .in1(N__39954),
            .in2(_gnd_net_),
            .in3(N__39860),
            .lcout(),
            .ltout(\ppm_encoder_1.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_12_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__51409),
            .in2(N__39930),
            .in3(N__39908),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_12_LC_14_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_14_12_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_14_12_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_14_12_5  (
            .in0(N__39909),
            .in1(N__45294),
            .in2(N__39927),
            .in3(N__45590),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59105),
            .ce(),
            .sr(N__57544));
    defparam \ppm_encoder_1.elevator_12_LC_14_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_14_12_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_14_12_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_14_12_6  (
            .in0(N__39861),
            .in1(N__39897),
            .in2(N__45375),
            .in3(N__39873),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59105),
            .ce(),
            .sr(N__57544));
    defparam \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_13_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_13_0  (
            .in0(N__40000),
            .in1(N__40851),
            .in2(N__44070),
            .in3(N__41357),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_13_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__47490),
            .in2(N__39849),
            .in3(N__39846),
            .lcout(\ppm_encoder_1.elevator_RNIC22D6Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_13_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_13_2  (
            .in0(N__40100),
            .in1(N__40063),
            .in2(N__44201),
            .in3(N__45513),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_13_3  (
            .in0(N__47164),
            .in1(N__40001),
            .in2(_gnd_net_),
            .in3(N__40101),
            .lcout(),
            .ltout(\ppm_encoder_1.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_13_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__51426),
            .in2(N__40083),
            .in3(N__40064),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_14_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_14_13_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_14_13_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_14_13_5  (
            .in0(N__40065),
            .in1(N__45389),
            .in2(N__43010),
            .in3(N__40080),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59112),
            .ce(),
            .sr(N__57554));
    defparam \ppm_encoder_1.throttle_11_LC_14_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_14_13_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_14_13_7  (
            .in0(N__40053),
            .in1(N__40017),
            .in2(N__40005),
            .in3(N__45390),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59112),
            .ce(),
            .sr(N__57554));
    defparam \ppm_encoder_1.throttle_RNI04QV2_9_LC_14_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI04QV2_9_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI04QV2_9_LC_14_14_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNI04QV2_9_LC_14_14_0  (
            .in0(N__40249),
            .in1(N__40205),
            .in2(N__41352),
            .in3(N__44054),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIV9PO6_9_LC_14_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIV9PO6_9_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIV9PO6_9_LC_14_14_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIV9PO6_9_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__46161),
            .in2(N__39987),
            .in3(N__39960),
            .lcout(\ppm_encoder_1.throttle_RNIV9PO6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_14_2  (
            .in0(N__51410),
            .in1(N__40212),
            .in2(_gnd_net_),
            .in3(N__39981),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_14_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_14_14_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__44660),
            .in2(N__39984),
            .in3(N__40188),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59122),
            .ce(N__44613),
            .sr(N__57563));
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_14_4 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_14_4  (
            .in0(N__40225),
            .in1(N__39980),
            .in2(N__45532),
            .in3(N__44166),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_14_5  (
            .in0(N__47171),
            .in1(N__40250),
            .in2(_gnd_net_),
            .in3(N__40226),
            .lcout(\ppm_encoder_1.N_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_14_6 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_14_6  (
            .in0(N__46389),
            .in1(N__46566),
            .in2(N__46140),
            .in3(N__40206),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_14_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_14_7  (
            .in0(N__46565),
            .in1(N__46388),
            .in2(_gnd_net_),
            .in3(N__46070),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIQTPV2_6_LC_14_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQTPV2_6_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQTPV2_6_LC_14_15_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIQTPV2_6_LC_14_15_0  (
            .in0(N__40172),
            .in1(N__40606),
            .in2(N__44073),
            .in3(N__41327),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIGQOO6_6_LC_14_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIGQOO6_6_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIGQOO6_6_LC_14_15_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIGQOO6_6_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__45834),
            .in2(N__40182),
            .in3(N__40179),
            .lcout(\ppm_encoder_1.throttle_RNIGQOO6Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_14_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_14_15_2 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.elevator_RNIAH7O2_6_LC_14_15_2  (
            .in0(N__40111),
            .in1(N__45483),
            .in2(N__40148),
            .in3(N__44125),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_14_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_14_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_14_15_3  (
            .in0(N__47165),
            .in1(N__40173),
            .in2(_gnd_net_),
            .in3(N__40144),
            .lcout(),
            .ltout(\ppm_encoder_1.N_292_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_15_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_15_4  (
            .in0(N__40112),
            .in1(_gnd_net_),
            .in2(N__40128),
            .in3(N__51456),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_14_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_14_15_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_14_15_5 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_14_15_5  (
            .in0(N__40125),
            .in1(N__40113),
            .in2(N__42975),
            .in3(N__45363),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59134),
            .ce(),
            .sr(N__57573));
    defparam \ppm_encoder_1.throttle_RNISVPV2_7_LC_14_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNISVPV2_7_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNISVPV2_7_LC_14_16_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_RNISVPV2_7_LC_14_16_0  (
            .in0(N__40343),
            .in1(N__40577),
            .in2(N__44071),
            .in3(N__41332),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNILVOO6_7_LC_14_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNILVOO6_7_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNILVOO6_7_LC_14_16_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.throttle_RNILVOO6_7_LC_14_16_1  (
            .in0(N__45924),
            .in1(_gnd_net_),
            .in2(N__40353),
            .in3(N__40350),
            .lcout(\ppm_encoder_1.throttle_RNILVOO6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_14_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_14_16_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNICJ7O2_7_LC_14_16_2  (
            .in0(N__40264),
            .in1(N__40309),
            .in2(N__44200),
            .in3(N__45516),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_16_3  (
            .in0(N__47169),
            .in1(N__40344),
            .in2(_gnd_net_),
            .in3(N__40265),
            .lcout(),
            .ltout(\ppm_encoder_1.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_16_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__51436),
            .in2(N__40326),
            .in3(N__40310),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_7_LC_14_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_14_16_5 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_14_16_5  (
            .in0(N__40311),
            .in1(N__40323),
            .in2(N__42930),
            .in3(N__45362),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59149),
            .ce(),
            .sr(N__57578));
    defparam \ppm_encoder_1.elevator_7_LC_14_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_14_16_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_14_16_6  (
            .in0(N__40266),
            .in1(N__40299),
            .in2(N__45400),
            .in3(N__40293),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59149),
            .ce(),
            .sr(N__57578));
    defparam \ppm_encoder_1.throttle_RNIU1QV2_8_LC_14_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIU1QV2_8_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIU1QV2_8_LC_14_17_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIU1QV2_8_LC_14_17_0  (
            .in0(N__40475),
            .in1(N__46232),
            .in2(N__44072),
            .in3(N__41348),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_14_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_14_17_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_14_17_1  (
            .in0(N__46257),
            .in1(_gnd_net_),
            .in2(N__40254),
            .in3(N__40482),
            .lcout(\ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_17_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_17_2  (
            .in0(N__40453),
            .in1(N__40417),
            .in2(N__44190),
            .in3(N__45546),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_17_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_17_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_17_3  (
            .in0(N__47177),
            .in1(N__40476),
            .in2(_gnd_net_),
            .in3(N__40454),
            .lcout(),
            .ltout(\ppm_encoder_1.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_17_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_17_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_17_4  (
            .in0(N__51415),
            .in1(_gnd_net_),
            .in2(N__40434),
            .in3(N__40418),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_8_LC_14_17_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_14_17_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_14_17_5  (
            .in0(N__40419),
            .in1(N__42885),
            .in2(N__45402),
            .in3(N__40431),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59161),
            .ce(),
            .sr(N__57585));
    defparam \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_14_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_14_18_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_14_18_0  (
            .in0(N__44059),
            .in1(N__40385),
            .in2(N__41356),
            .in3(N__44816),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_14_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_14_18_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_14_18_1  (
            .in0(N__44325),
            .in1(_gnd_net_),
            .in2(N__40407),
            .in3(N__40404),
            .lcout(\ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_14_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_14_18_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_14_18_2  (
            .in0(N__40397),
            .in1(N__40364),
            .in2(N__45561),
            .in3(N__44194),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_14_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_14_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_14_18_3  (
            .in0(N__47150),
            .in1(N__40398),
            .in2(_gnd_net_),
            .in3(N__40386),
            .lcout(),
            .ltout(\ppm_encoder_1.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_18_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_18_4  (
            .in0(N__51452),
            .in1(_gnd_net_),
            .in2(N__40368),
            .in3(N__40365),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_18_5 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_18_5  (
            .in0(N__45759),
            .in1(N__46570),
            .in2(N__46444),
            .in3(N__40611),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIGUOT2_10_LC_14_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIGUOT2_10_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIGUOT2_10_LC_14_18_6 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \ppm_encoder_1.throttle_RNIGUOT2_10_LC_14_18_6  (
            .in0(N__44058),
            .in1(N__40553),
            .in2(N__41355),
            .in3(N__46302),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48854),
            .lcout(\ppm_encoder_1.N_2150_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_14_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_14_19_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNI02LH2_10_LC_14_19_1  (
            .in0(N__40526),
            .in1(N__40502),
            .in2(N__45560),
            .in3(N__44195),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI7T1D6_10_LC_14_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI7T1D6_10_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI7T1D6_10_LC_14_19_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI7T1D6_10_LC_14_19_2  (
            .in0(N__46608),
            .in1(_gnd_net_),
            .in2(N__40590),
            .in3(N__40587),
            .lcout(\ppm_encoder_1.elevator_RNI7T1D6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_19_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_19_3 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_19_3  (
            .in0(N__45900),
            .in1(N__46569),
            .in2(N__46445),
            .in3(N__40581),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_19_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_19_4  (
            .in0(N__40557),
            .in1(N__47128),
            .in2(_gnd_net_),
            .in3(N__40527),
            .lcout(),
            .ltout(\ppm_encoder_1.N_296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_14_19_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_14_19_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__51451),
            .in2(N__40506),
            .in3(N__40503),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_14_19_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_14_19_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_14_19_7  (
            .in0(N__46977),
            .in1(N__51450),
            .in2(_gnd_net_),
            .in3(N__43794),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_14_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_14_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52467),
            .lcout(drone_H_disp_front_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59202),
            .ce(N__50692),
            .sr(N__57611));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_21_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_21_0  (
            .in0(N__40689),
            .in1(N__42770),
            .in2(N__40662),
            .in3(N__42810),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_21_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_21_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_14_21_1  (
            .in0(N__44704),
            .in1(N__40710),
            .in2(_gnd_net_),
            .in3(N__40698),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59217),
            .ce(N__44612),
            .sr(N__57618));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_21_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_14_21_2  (
            .in0(N__40683),
            .in1(N__40674),
            .in2(_gnd_net_),
            .in3(N__44705),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59217),
            .ce(N__44612),
            .sr(N__57618));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_14_21_3  (
            .in0(N__44703),
            .in1(N__40653),
            .in2(_gnd_net_),
            .in3(N__44346),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59217),
            .ce(N__44612),
            .sr(N__57618));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_21_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_21_4  (
            .in0(N__42720),
            .in1(N__40644),
            .in2(N__41925),
            .in3(N__41769),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_14_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_14_21_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_14_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_14_21_5  (
            .in0(N__44706),
            .in1(N__40638),
            .in2(_gnd_net_),
            .in3(N__46188),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59217),
            .ce(N__44612),
            .sr(N__57618));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_21_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_21_6  (
            .in0(N__40626),
            .in1(N__44519),
            .in2(N__42696),
            .in3(N__40620),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_14_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_14_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_14_22_0  (
            .in0(N__42076),
            .in1(N__42025),
            .in2(N__42057),
            .in3(N__43586),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_14_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_14_22_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_14_22_3  (
            .in0(N__40800),
            .in1(_gnd_net_),
            .in2(N__44727),
            .in3(N__44301),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59234),
            .ce(N__44592),
            .sr(N__57625));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_14_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_14_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_14_22_5  (
            .in0(N__44720),
            .in1(N__50214),
            .in2(_gnd_net_),
            .in3(N__40791),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59234),
            .ce(N__44592),
            .sr(N__57625));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_14_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_14_22_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_14_22_6  (
            .in0(N__42075),
            .in1(N__40779),
            .in2(N__40773),
            .in3(N__44455),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_14_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_14_22_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_14_22_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_14_22_7  (
            .in0(N__44721),
            .in1(_gnd_net_),
            .in2(N__41562),
            .in3(N__43824),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59234),
            .ce(N__44592),
            .sr(N__57625));
    defparam \ppm_encoder_1.counter_0_LC_14_23_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_14_23_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_14_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__44459),
            .in2(N__40764),
            .in3(N__40763),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_1_LC_14_23_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_14_23_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_14_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__42078),
            .in2(_gnd_net_),
            .in3(N__40743),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_2_LC_14_23_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_14_23_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_14_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__42026),
            .in2(_gnd_net_),
            .in3(N__40740),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_3_LC_14_23_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_14_23_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_14_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__42056),
            .in2(_gnd_net_),
            .in3(N__40737),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_4_LC_14_23_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_14_23_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_14_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(N__42746),
            .in2(_gnd_net_),
            .in3(N__40734),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_5_LC_14_23_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_14_23_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_14_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_14_23_5  (
            .in0(_gnd_net_),
            .in1(N__42789),
            .in2(_gnd_net_),
            .in3(N__40830),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_6_LC_14_23_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_14_23_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_14_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__42809),
            .in2(_gnd_net_),
            .in3(N__40827),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_7_LC_14_23_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_14_23_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_14_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__42769),
            .in2(_gnd_net_),
            .in3(N__40824),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__59252),
            .ce(),
            .sr(N__41046));
    defparam \ppm_encoder_1.counter_8_LC_14_24_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_14_24_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_14_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(N__42692),
            .in2(_gnd_net_),
            .in3(N__40821),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_9_LC_14_24_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_14_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_14_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(N__44518),
            .in2(_gnd_net_),
            .in3(N__40818),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_10_LC_14_24_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_14_24_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_14_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(N__44551),
            .in2(_gnd_net_),
            .in3(N__40815),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_11_LC_14_24_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_14_24_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_14_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__44491),
            .in2(_gnd_net_),
            .in3(N__40812),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_12_LC_14_24_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_14_24_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_14_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(N__42719),
            .in2(_gnd_net_),
            .in3(N__40809),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_13_LC_14_24_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_14_24_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_14_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__41921),
            .in2(_gnd_net_),
            .in3(N__40806),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_14_LC_14_24_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_14_24_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_14_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__41945),
            .in2(_gnd_net_),
            .in3(N__40803),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_15_LC_14_24_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_14_24_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_14_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(N__43103),
            .in2(_gnd_net_),
            .in3(N__41058),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__59267),
            .ce(),
            .sr(N__41045));
    defparam \ppm_encoder_1.counter_16_LC_14_25_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_14_25_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_14_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__43143),
            .in2(_gnd_net_),
            .in3(N__41055),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__59279),
            .ce(),
            .sr(N__41044));
    defparam \ppm_encoder_1.counter_17_LC_14_25_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_14_25_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_14_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(N__43124),
            .in2(_gnd_net_),
            .in3(N__41052),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__59279),
            .ce(),
            .sr(N__41044));
    defparam \ppm_encoder_1.counter_18_LC_14_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_14_25_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_14_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__43158),
            .in2(_gnd_net_),
            .in3(N__41049),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59279),
            .ce(),
            .sr(N__41044));
    defparam \ppm_encoder_1.aileron_0_LC_15_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_0_LC_15_10_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_0_LC_15_10_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.aileron_0_LC_15_10_4  (
            .in0(N__45405),
            .in1(N__43289),
            .in2(_gnd_net_),
            .in3(N__50233),
            .lcout(\ppm_encoder_1.aileronZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59099),
            .ce(),
            .sr(N__57537));
    defparam \scaler_4.source_data_1_4_LC_15_11_4 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_15_11_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_15_11_4 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_15_11_4  (
            .in0(N__41021),
            .in1(N__41217),
            .in2(N__46817),
            .in3(N__41173),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59106),
            .ce(),
            .sr(N__57545));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_12_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__40982),
            .in2(_gnd_net_),
            .in3(N__57842),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_12_1 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_12_1  (
            .in0(N__57843),
            .in1(N__41072),
            .in2(N__46353),
            .in3(N__48743),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59113),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_12_3  (
            .in0(N__46332),
            .in1(N__48330),
            .in2(_gnd_net_),
            .in3(N__40849),
            .lcout(),
            .ltout(\ppm_encoder_1.N_313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_12_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__46501),
            .in2(N__41088),
            .in3(N__46664),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_12_5 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_12_5  (
            .in0(N__47172),
            .in1(N__43482),
            .in2(_gnd_net_),
            .in3(N__43351),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_15_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_15_12_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_15_12_7  (
            .in0(N__47173),
            .in1(N__43483),
            .in2(_gnd_net_),
            .in3(N__43350),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_13_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_13_0 .LUT_INIT=16'b1101110111001110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_13_0  (
            .in0(N__48740),
            .in1(N__57887),
            .in2(N__49082),
            .in3(N__43485),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59123),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_13_1 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_13_1  (
            .in0(N__57886),
            .in1(N__43409),
            .in2(N__43170),
            .in3(N__48742),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59123),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_13_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__43316),
            .in2(_gnd_net_),
            .in3(N__43699),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_13_3 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_13_3  (
            .in0(N__57885),
            .in1(N__43388),
            .in2(N__41073),
            .in3(N__48741),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59123),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIH72D6_12_LC_15_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIH72D6_12_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIH72D6_12_LC_15_13_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIH72D6_12_LC_15_13_4  (
            .in0(N__46641),
            .in1(N__41085),
            .in2(_gnd_net_),
            .in3(N__41079),
            .lcout(\ppm_encoder_1.elevator_RNIH72D6Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_13_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_13_5  (
            .in0(N__46352),
            .in1(N__47162),
            .in2(N__51448),
            .in3(N__49061),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_13_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_13_6  (
            .in0(N__48739),
            .in1(N__57888),
            .in2(N__41262),
            .in3(N__41103),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59123),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_15_13_7 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_15_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_15_13_7  (
            .in0(N__41259),
            .in1(N__41213),
            .in2(_gnd_net_),
            .in3(N__41175),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_1_LC_15_14_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_1_LC_15_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_1_LC_15_14_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \pid_side.source_pid_1_esr_1_LC_15_14_0  (
            .in0(N__47745),
            .in1(N__44854),
            .in2(N__49695),
            .in3(N__45625),
            .lcout(side_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59135),
            .ce(N__48036),
            .sr(N__47994));
    defparam \pid_side.source_pid_1_esr_2_LC_15_14_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_2_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_2_LC_15_14_1 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \pid_side.source_pid_1_esr_2_LC_15_14_1  (
            .in0(N__45626),
            .in1(N__49681),
            .in2(N__44859),
            .in3(N__49755),
            .lcout(side_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59135),
            .ce(N__48036),
            .sr(N__47994));
    defparam \pid_side.source_pid_1_esr_3_LC_15_14_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_3_LC_15_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_3_LC_15_14_2 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \pid_side.source_pid_1_esr_3_LC_15_14_2  (
            .in0(N__49728),
            .in1(N__44858),
            .in2(N__49696),
            .in3(N__45627),
            .lcout(side_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59135),
            .ce(N__48036),
            .sr(N__47994));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_15_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_15_14_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_15_14_3  (
            .in0(N__43481),
            .in1(N__43692),
            .in2(N__43445),
            .in3(N__43517),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_14_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_14_5  (
            .in0(N__43480),
            .in1(N__43436),
            .in2(N__48735),
            .in3(N__43691),
            .lcout(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_14_6 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43410),
            .in3(N__41102),
            .lcout(\ppm_encoder_1.N_221 ),
            .ltout(\ppm_encoder_1.N_221_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_14_7  (
            .in0(N__48635),
            .in1(N__43479),
            .in2(N__41091),
            .in3(N__43435),
            .lcout(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_15_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_15_0  (
            .in0(N__41848),
            .in1(N__46952),
            .in2(N__45514),
            .in3(N__44123),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_15_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_15_15_1 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_15_15_1  (
            .in0(N__41873),
            .in1(N__46800),
            .in2(N__41354),
            .in3(N__44048),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFISN6_4_LC_15_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFISN6_4_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFISN6_4_LC_15_15_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIFISN6_4_LC_15_15_2  (
            .in0(N__44424),
            .in1(_gnd_net_),
            .in2(N__41385),
            .in3(N__41382),
            .lcout(\ppm_encoder_1.elevator_RNIFISN6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_15_4 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_15_4  (
            .in0(N__43189),
            .in1(N__51265),
            .in2(N__45515),
            .in3(N__44124),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_15_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_15_15_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_15_15_5  (
            .in0(N__43357),
            .in1(N__43389),
            .in2(N__43317),
            .in3(N__48642),
            .lcout(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_15_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_15_15_6 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_15_15_6  (
            .in0(N__44049),
            .in1(N__43223),
            .in2(N__41376),
            .in3(N__45971),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIKNSN6_5_LC_15_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIKNSN6_5_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIKNSN6_5_LC_15_15_7 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIKNSN6_5_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__46004),
            .in2(N__41373),
            .in3(N__41370),
            .lcout(\ppm_encoder_1.elevator_RNIKNSN6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_15_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_15_16_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.elevator_RNI077O2_1_LC_15_16_0  (
            .in0(N__41461),
            .in1(N__41509),
            .in2(N__45545),
            .in3(N__44170),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIUINC6_1_LC_15_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIUINC6_1_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIUINC6_1_LC_15_16_1 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIUINC6_1_LC_15_16_1  (
            .in0(N__43845),
            .in1(N__41268),
            .in2(N__41364),
            .in3(N__41328),
            .lcout(\ppm_encoder_1.throttle_RNIUINC6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIEES71_1_LC_15_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIEES71_1_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIEES71_1_LC_15_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIEES71_1_LC_15_16_2  (
            .in0(N__41410),
            .in1(N__43703),
            .in2(N__43809),
            .in3(N__48696),
            .lcout(\ppm_encoder_1.throttle_m_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_16_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_16_3  (
            .in0(N__47170),
            .in1(N__41462),
            .in2(_gnd_net_),
            .in3(N__41411),
            .lcout(),
            .ltout(\ppm_encoder_1.N_287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_16_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__51411),
            .in2(N__41565),
            .in3(N__41510),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_1_LC_15_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_1_LC_15_16_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_1_LC_15_16_5 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \ppm_encoder_1.aileron_1_LC_15_16_5  (
            .in0(N__45376),
            .in1(N__41546),
            .in2(N__41526),
            .in3(N__41511),
            .lcout(\ppm_encoder_1.aileronZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59162),
            .ce(),
            .sr(N__57586));
    defparam \ppm_encoder_1.elevator_1_LC_15_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_1_LC_15_16_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_1_LC_15_16_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \ppm_encoder_1.elevator_1_LC_15_16_6  (
            .in0(N__41463),
            .in1(N__41496),
            .in2(N__41487),
            .in3(N__45380),
            .lcout(\ppm_encoder_1.elevatorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59162),
            .ce(),
            .sr(N__57586));
    defparam \ppm_encoder_1.throttle_1_LC_15_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_15_16_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_15_16_7  (
            .in0(N__41451),
            .in1(N__41439),
            .in2(N__45403),
            .in3(N__41412),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59162),
            .ce(),
            .sr(N__57586));
    defparam \ppm_encoder_1.elevator_RNINSH16_0_LC_15_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.elevator_RNINSH16_0_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNINSH16_0_LC_15_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNINSH16_0_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__43638),
            .in2(N__46044),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__43841),
            .in2(N__41400),
            .in3(N__41391),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_17_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__44276),
            .in2(N__43758),
            .in3(N__41388),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_17_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__44237),
            .in2(N__43968),
            .in3(N__41685),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_17_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__44417),
            .in2(N__41682),
            .in3(N__41670),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_17_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__46005),
            .in2(N__41667),
            .in3(N__41655),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_17_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__45833),
            .in2(N__41652),
            .in3(N__41640),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_17_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__45923),
            .in2(N__41637),
            .in3(N__41628),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_18_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__46253),
            .in2(N__41625),
            .in3(N__41616),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_18_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__46160),
            .in2(N__41613),
            .in3(N__41598),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_18_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__46604),
            .in2(N__41595),
            .in3(N__41586),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_18_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__47483),
            .in2(N__41583),
            .in3(N__41568),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_18_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__46637),
            .in2(N__41757),
            .in3(N__41742),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_18_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__44393),
            .in2(N__41739),
            .in3(N__41727),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_18_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__44321),
            .in2(N__41724),
            .in3(N__41715),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_18_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__45795),
            .in2(N__45816),
            .in3(N__41712),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__43071),
            .in2(_gnd_net_),
            .in3(N__41709),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__44259),
            .in2(_gnd_net_),
            .in3(N__41706),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__41700),
            .in2(_gnd_net_),
            .in3(N__41703),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_15_19_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_15_19_3 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_18_LC_15_19_3  (
            .in0(N__48851),
            .in1(N__47883),
            .in2(N__49105),
            .in3(N__49074),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_15_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_15_19_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__41694),
            .in2(_gnd_net_),
            .in3(N__43618),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_19_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_19_5  (
            .in0(N__47127),
            .in1(N__41877),
            .in2(_gnd_net_),
            .in3(N__41853),
            .lcout(\ppm_encoder_1.N_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_19_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_19_6 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_19_6  (
            .in0(N__47109),
            .in1(N__57896),
            .in2(N__51449),
            .in3(N__48852),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59203),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_15_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_15_20_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_15_20_1  (
            .in0(N__46092),
            .in1(N__44684),
            .in2(_gnd_net_),
            .in3(N__46932),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59218),
            .ce(N__44602),
            .sr(N__57619));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_15_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_15_20_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_15_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_15_20_2  (
            .in0(N__44685),
            .in1(N__51246),
            .in2(_gnd_net_),
            .in3(N__45951),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59218),
            .ce(N__44602),
            .sr(N__57619));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_15_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_15_20_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_15_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_15_20_3  (
            .in0(N__41829),
            .in1(N__47511),
            .in2(_gnd_net_),
            .in3(N__44681),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59218),
            .ce(N__44602),
            .sr(N__57619));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_20_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_20_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_20_4  (
            .in0(N__44492),
            .in1(N__41823),
            .in2(N__41793),
            .in3(N__44552),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_15_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_15_20_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_15_20_5  (
            .in0(N__41817),
            .in1(N__44682),
            .in2(_gnd_net_),
            .in3(N__41805),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59218),
            .ce(N__44602),
            .sr(N__57619));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_15_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_15_20_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_15_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_15_20_6  (
            .in0(N__44683),
            .in1(N__41784),
            .in2(_gnd_net_),
            .in3(N__46653),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59218),
            .ce(N__44602),
            .sr(N__57619));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_15_21_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_15_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__41763),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_15_21_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_15_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__42003),
            .in2(N__42449),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_15_21_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_15_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__41979),
            .in2(N__42439),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_15_21_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_15_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__41901),
            .in2(N__42446),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_15_21_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_15_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__41895),
            .in2(N__42440),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_15_21_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_15_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__41889),
            .in2(N__42447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_15_21_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_15_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__41883),
            .in2(N__42441),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_15_21_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_15_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__42084),
            .in2(N__42448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_15_22_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_15_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__42504),
            .in2(N__42450),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_15_22_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_15_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__42468),
            .in2(N__42442),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42087),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_15_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_15_22_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_15_22_3  (
            .in0(N__44733),
            .in1(N__43104),
            .in2(N__46869),
            .in3(N__41946),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_22_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_22_4  (
            .in0(N__43536),
            .in1(N__42052),
            .in2(N__42027),
            .in3(N__42077),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_22_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_22_5  (
            .in0(N__42051),
            .in1(N__42033),
            .in2(N__44622),
            .in3(N__42021),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_22_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_22_7  (
            .in0(N__42787),
            .in1(N__41997),
            .in2(N__42747),
            .in3(N__41988),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_23_0  (
            .in0(N__41973),
            .in1(N__44438),
            .in2(N__43083),
            .in3(N__42672),
            .lcout(\ppm_encoder_1.N_232 ),
            .ltout(\ppm_encoder_1.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_23_1 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_23_1  (
            .in0(N__44988),
            .in1(N__43608),
            .in2(N__41967),
            .in3(N__43537),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_23_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__41944),
            .in2(_gnd_net_),
            .in3(N__41920),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_15_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_15_23_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_15_23_3  (
            .in0(N__42808),
            .in1(N__42788),
            .in2(N__42771),
            .in3(N__42745),
            .lcout(),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_15_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_15_23_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.counter_RNIAEV01_8_LC_15_23_4  (
            .in0(N__42726),
            .in1(N__42718),
            .in2(N__42699),
            .in3(N__42691),
            .lcout(\ppm_encoder_1.N_139_17 ),
            .ltout(\ppm_encoder_1.N_139_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_15_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_15_23_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_15_23_5  (
            .in0(N__44439),
            .in1(N__42666),
            .in2(N__42657),
            .in3(N__43082),
            .lcout(\ppm_encoder_1.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIGKTC2_20_LC_15_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGKTC2_20_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGKTC2_20_LC_15_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGKTC2_20_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__42627),
            .in2(_gnd_net_),
            .in3(N__42561),
            .lcout(\pid_front.error_p_reg_esr_RNIGKTC2Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_15_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_15_24_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_15_24_0  (
            .in0(N__42491),
            .in1(N__43120),
            .in2(N__45011),
            .in3(N__43141),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_16_LC_15_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_16_LC_15_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_16_LC_15_24_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ppm_encoder_1.pulses2count_16_LC_15_24_1  (
            .in0(N__46907),
            .in1(N__44772),
            .in2(N__42495),
            .in3(N__48870),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59280),
            .ce(),
            .sr(N__57640));
    defparam \ppm_encoder_1.pulses2count_18_LC_15_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_18_LC_15_24_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_18_LC_15_24_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_18_LC_15_24_4  (
            .in0(N__48869),
            .in1(N__46908),
            .in2(N__42480),
            .in3(N__49113),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59280),
            .ce(),
            .sr(N__57640));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_24_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__42476),
            .in2(_gnd_net_),
            .in3(N__43156),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_15_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_15_24_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNI637H_18_LC_15_24_6  (
            .in0(N__43157),
            .in1(N__43142),
            .in2(N__43128),
            .in3(N__43102),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_15_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_15_24_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_15_24_7  (
            .in0(N__49083),
            .in1(N__44771),
            .in2(_gnd_net_),
            .in3(N__48868),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_20_LC_15_25_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_15_25_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_15_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_20_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59502),
            .lcout(\pid_front.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59289),
            .ce(N__49368),
            .sr(N__57644));
    defparam \pid_side.source_pid_1_10_LC_16_10_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_10_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_10_LC_16_10_2 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_side.source_pid_1_10_LC_16_10_2  (
            .in0(N__47578),
            .in1(N__45695),
            .in2(N__43033),
            .in3(N__49967),
            .lcout(side_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59107),
            .ce(),
            .sr(N__47986));
    defparam \pid_side.source_pid_1_11_LC_16_10_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_11_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_11_LC_16_10_3 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_side.source_pid_1_11_LC_16_10_3  (
            .in0(N__45696),
            .in1(N__47579),
            .in2(N__43006),
            .in3(N__49928),
            .lcout(side_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59107),
            .ce(),
            .sr(N__47986));
    defparam \pid_side.source_pid_1_6_LC_16_10_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_6_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_6_LC_16_10_4 .LUT_INIT=16'b1101100011111010;
    LogicCell40 \pid_side.source_pid_1_6_LC_16_10_4  (
            .in0(N__47580),
            .in1(N__49568),
            .in2(N__42961),
            .in3(N__45697),
            .lcout(side_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59107),
            .ce(),
            .sr(N__47986));
    defparam \pid_side.source_pid_1_7_LC_16_10_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_7_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_7_LC_16_10_5 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \pid_side.source_pid_1_7_LC_16_10_5  (
            .in0(N__45698),
            .in1(N__49542),
            .in2(N__42916),
            .in3(N__47581),
            .lcout(side_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59107),
            .ce(),
            .sr(N__47986));
    defparam \pid_side.source_pid_1_8_LC_16_10_6 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_8_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_8_LC_16_10_6 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_side.source_pid_1_8_LC_16_10_6  (
            .in0(N__47582),
            .in1(N__45699),
            .in2(N__42871),
            .in3(N__49509),
            .lcout(side_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59107),
            .ce(),
            .sr(N__47986));
    defparam \pid_side.source_pid_1_9_LC_16_10_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_9_LC_16_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_9_LC_16_10_7 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_side.source_pid_1_9_LC_16_10_7  (
            .in0(N__45700),
            .in1(N__47583),
            .in2(N__42835),
            .in3(N__49488),
            .lcout(side_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59107),
            .ce(),
            .sr(N__47986));
    defparam \pid_side.state_RNID6CB8_1_LC_16_11_2 .C_ON=1'b0;
    defparam \pid_side.state_RNID6CB8_1_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNID6CB8_1_LC_16_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNID6CB8_1_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__47577),
            .in2(_gnd_net_),
            .in3(N__47982),
            .lcout(\pid_side.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_0_LC_16_11_6 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_0_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_0_LC_16_11_6 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \pid_side.source_pid_1_esr_0_LC_16_11_6  (
            .in0(N__47769),
            .in1(N__44843),
            .in2(N__49697),
            .in3(N__45613),
            .lcout(side_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59114),
            .ce(N__48020),
            .sr(N__47983));
    defparam \pid_side.source_pid_1_esr_5_LC_16_11_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_5_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_5_LC_16_11_7 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \pid_side.source_pid_1_esr_5_LC_16_11_7  (
            .in0(N__45643),
            .in1(N__45701),
            .in2(N__49619),
            .in3(N__45663),
            .lcout(side_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59114),
            .ce(N__48020),
            .sr(N__47983));
    defparam \pid_side.source_pid_1_esr_4_LC_16_12_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_4_LC_16_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_4_LC_16_12_0 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \pid_side.source_pid_1_esr_4_LC_16_12_0  (
            .in0(N__49698),
            .in1(N__45702),
            .in2(N__49620),
            .in3(N__45614),
            .lcout(side_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59124),
            .ce(N__48021),
            .sr(N__47987));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_13_0  (
            .in0(N__43437),
            .in1(N__45870),
            .in2(_gnd_net_),
            .in3(N__43668),
            .lcout(\ppm_encoder_1.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_13_1  (
            .in0(N__47151),
            .in1(N__43227),
            .in2(_gnd_net_),
            .in3(N__43200),
            .lcout(\ppm_encoder_1.N_291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_16_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_16_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__48274),
            .in2(_gnd_net_),
            .in3(N__48736),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_13_4 .LUT_INIT=16'b0100000010101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_13_4  (
            .in0(N__43355),
            .in1(N__47152),
            .in2(N__51432),
            .in3(N__46360),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_13_5 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_13_5  (
            .in0(N__57889),
            .in1(N__43356),
            .in2(N__43161),
            .in3(N__48738),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59136),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_16_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_16_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_16_13_6  (
            .in0(N__43438),
            .in1(N__43387),
            .in2(N__43359),
            .in3(N__43484),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_16_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_16_13_7 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__48275),
            .in2(N__43449),
            .in3(N__48737),
            .lcout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_14_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_14_0 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_14_0  (
            .in0(N__57890),
            .in1(N__51382),
            .in2(N__43446),
            .in3(N__48645),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59150),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_14_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__43722),
            .in2(_gnd_net_),
            .in3(N__43743),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_16_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_16_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__43382),
            .in2(_gnd_net_),
            .in3(N__43408),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_16_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_16_14_3 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_16_14_3  (
            .in0(N__43383),
            .in1(N__43358),
            .in2(N__43320),
            .in3(N__43312),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_16_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_16_14_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43296),
            .in3(N__48643),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_5 .LUT_INIT=16'b1111111101010010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_5  (
            .in0(N__48644),
            .in1(N__48994),
            .in2(N__43728),
            .in3(N__57894),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59150),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_6 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_6  (
            .in0(N__43745),
            .in1(N__51381),
            .in2(N__57902),
            .in3(N__48646),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59150),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_14_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__43744),
            .in2(_gnd_net_),
            .in3(N__43723),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_15_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_15_0  (
            .in0(N__47000),
            .in1(N__43793),
            .in2(N__44159),
            .in3(N__44020),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_15_1 .LUT_INIT=16'b1000111110001111;
    LogicCell40 \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_15_1  (
            .in0(N__45504),
            .in1(N__47039),
            .in2(N__43761),
            .in3(N__44280),
            .lcout(\ppm_encoder_1.elevator_RNIPVQ05Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_16_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_16_15_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_16_15_2  (
            .in0(N__43746),
            .in1(N__43724),
            .in2(N__43704),
            .in3(N__48636),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIGCMK2_0_LC_16_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIGCMK2_0_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIGCMK2_0_LC_16_15_3 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIGCMK2_0_LC_16_15_3  (
            .in0(N__43667),
            .in1(N__50240),
            .in2(N__43644),
            .in3(N__44126),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0 ),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_15_4 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_15_4  (
            .in0(N__45879),
            .in1(N__46040),
            .in2(N__43641),
            .in3(N__45503),
            .lcout(\ppm_encoder_1.elevator_RNIHNQ05Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_16_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_16_15_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__43510),
            .in2(_gnd_net_),
            .in3(N__43573),
            .lcout(\ppm_encoder_1.PPM_STATE_53_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_16_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_16_15_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_16_15_6 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_16_15_6  (
            .in0(N__43511),
            .in1(_gnd_net_),
            .in2(N__43560),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59163),
            .ce(),
            .sr(N__57587));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_16_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_16_15_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_16_15_7 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_16_15_7  (
            .in0(N__43628),
            .in1(N__43574),
            .in2(N__43539),
            .in3(N__43556),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59163),
            .ce(),
            .sr(N__57587));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_16_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_16_0  (
            .in0(N__43865),
            .in1(N__47161),
            .in2(_gnd_net_),
            .in3(N__44226),
            .lcout(\ppm_encoder_1.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIMIMK2_3_LC_16_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIMIMK2_3_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIMIMK2_3_LC_16_16_1 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIMIMK2_3_LC_16_16_1  (
            .in0(N__44225),
            .in1(N__43915),
            .in2(N__44199),
            .in3(N__44021),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIT3R05_3_LC_16_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIT3R05_3_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIT3R05_3_LC_16_16_2 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \ppm_encoder_1.elevator_RNIT3R05_3_LC_16_16_2  (
            .in0(N__43864),
            .in1(N__44241),
            .in2(N__43971),
            .in3(N__45559),
            .lcout(\ppm_encoder_1.elevator_RNIT3R05Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_16_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_16_3  (
            .in0(N__51404),
            .in1(N__43959),
            .in2(_gnd_net_),
            .in3(N__43916),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_3_LC_16_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_3_LC_16_16_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_3_LC_16_16_4 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \ppm_encoder_1.aileron_3_LC_16_16_4  (
            .in0(N__45381),
            .in1(N__43917),
            .in2(N__43953),
            .in3(N__43929),
            .lcout(\ppm_encoder_1.aileronZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59176),
            .ce(),
            .sr(N__57598));
    defparam \ppm_encoder_1.elevator_3_LC_16_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_3_LC_16_16_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_3_LC_16_16_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.elevator_3_LC_16_16_6  (
            .in0(N__43866),
            .in1(N__43902),
            .in2(N__45404),
            .in3(N__43890),
            .lcout(\ppm_encoder_1.elevatorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59176),
            .ce(),
            .sr(N__57598));
    defparam \ppm_encoder_1.init_pulses_1_LC_16_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_16_17_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_16_17_0 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_16_17_0  (
            .in0(N__47277),
            .in1(N__47467),
            .in2(N__43854),
            .in3(N__48189),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59192),
            .ce(),
            .sr(N__57605));
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_17_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_17_2  (
            .in0(N__47815),
            .in1(N__49025),
            .in2(_gnd_net_),
            .in3(N__48789),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_17_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_17_3 .LUT_INIT=16'b1111110001010101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_17_3  (
            .in0(N__46684),
            .in1(N__46447),
            .in2(N__47822),
            .in3(N__46553),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_17_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_17_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_17_4  (
            .in0(N__46448),
            .in1(N__45779),
            .in2(N__46572),
            .in3(N__46685),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_2_LC_16_17_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_16_17_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_16_17_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_16_17_5  (
            .in0(N__47466),
            .in1(N__48153),
            .in2(N__47318),
            .in3(N__44286),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59192),
            .ce(),
            .sr(N__57605));
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_16_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_16_17_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI87N01_2_LC_16_17_6  (
            .in0(N__45778),
            .in1(N__49026),
            .in2(_gnd_net_),
            .in3(N__48790),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_17_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_17_7 .LUT_INIT=16'b1110111000001111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_17_7  (
            .in0(N__48236),
            .in1(N__46449),
            .in2(N__46689),
            .in3(N__46554),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_17_LC_16_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_16_18_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_16_18_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_16_18_0  (
            .in0(N__47422),
            .in1(N__49128),
            .in2(N__47319),
            .in3(N__44265),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59204),
            .ce(),
            .sr(N__57612));
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_16_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_16_18_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_16_18_1  (
            .in0(N__48794),
            .in1(N__45025),
            .in2(_gnd_net_),
            .in3(N__49078),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_16_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_16_18_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_16_18_2  (
            .in0(N__49077),
            .in1(_gnd_net_),
            .in2(N__45032),
            .in3(N__48793),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_3_LC_16_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_16_18_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_16_18_3  (
            .in0(N__47327),
            .in1(N__48132),
            .in2(N__44253),
            .in3(N__47424),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59204),
            .ce(),
            .sr(N__57612));
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_16_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_16_18_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI98N01_3_LC_16_18_4  (
            .in0(N__49075),
            .in1(N__48232),
            .in2(_gnd_net_),
            .in3(N__48791),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_4_LC_16_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_16_18_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_16_18_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_16_18_6  (
            .in0(N__47423),
            .in1(N__48111),
            .in2(N__47320),
            .in3(N__44430),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59204),
            .ce(),
            .sr(N__57612));
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_16_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_16_18_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_16_18_7  (
            .in0(N__48792),
            .in1(N__46108),
            .in2(_gnd_net_),
            .in3(N__49076),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_16_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_16_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__48291),
            .in2(_gnd_net_),
            .in3(N__48832),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_16_19_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_16_19_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_16_19_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_16_19_3  (
            .in0(N__47417),
            .in1(N__49233),
            .in2(N__47348),
            .in3(N__44406),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59219),
            .ce(),
            .sr(N__57620));
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_19_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_19_4  (
            .in0(N__49073),
            .in1(N__47836),
            .in2(_gnd_net_),
            .in3(N__48833),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_18_LC_16_19_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_16_19_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_16_19_6  (
            .in0(N__47418),
            .in1(N__48519),
            .in2(N__47349),
            .in3(N__44382),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59219),
            .ce(),
            .sr(N__57620));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_19_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_19_7 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_19_7  (
            .in0(N__47837),
            .in1(N__46573),
            .in2(N__46453),
            .in3(N__44376),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_14_LC_16_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_16_20_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_16_20_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_16_20_0  (
            .in0(N__47419),
            .in1(N__49206),
            .in2(N__47350),
            .in3(N__44334),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59235),
            .ce(),
            .sr(N__57626));
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_16_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_16_20_1 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_16_20_1  (
            .in0(N__44830),
            .in1(_gnd_net_),
            .in2(N__48867),
            .in3(N__49069),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_20_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_20_2  (
            .in0(N__49067),
            .in1(N__48834),
            .in2(_gnd_net_),
            .in3(N__44831),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_20_3 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_20_3  (
            .in0(N__44832),
            .in1(N__46574),
            .in2(N__46454),
            .in3(N__44820),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_16_20_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_16_20_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_16_20_4  (
            .in0(N__47420),
            .in1(N__49182),
            .in2(N__47351),
            .in3(N__44787),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59235),
            .ce(),
            .sr(N__57626));
    defparam \ppm_encoder_1.init_pulses_16_LC_16_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_16_20_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_16_20_6  (
            .in0(N__47421),
            .in1(N__49155),
            .in2(N__47352),
            .in3(N__44778),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59235),
            .ce(),
            .sr(N__57626));
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_16_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_16_20_7 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_16_20_7  (
            .in0(N__44765),
            .in1(_gnd_net_),
            .in2(N__48866),
            .in3(N__49068),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_16_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_16_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_16_21_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_16_21_2  (
            .in0(N__44751),
            .in1(N__44725),
            .in2(_gnd_net_),
            .in3(N__44739),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59253),
            .ce(N__44580),
            .sr(N__57632));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_16_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_16_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_16_21_4  (
            .in0(N__44726),
            .in1(N__44640),
            .in2(_gnd_net_),
            .in3(N__44631),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59253),
            .ce(N__44580),
            .sr(N__57632));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_16_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_16_22_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__57844),
            .in2(_gnd_net_),
            .in3(N__48853),
            .lcout(\ppm_encoder_1.N_2150_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_16_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_16_22_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.counter_RNIK1KG_0_LC_16_22_2  (
            .in0(N__44553),
            .in1(N__44523),
            .in2(N__44496),
            .in3(N__44463),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_14_LC_16_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_16_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_16_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_14_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59458),
            .lcout(\pid_front.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59281),
            .ce(N__49374),
            .sr(N__57641));
    defparam \ppm_encoder_1.pulses2count_17_LC_16_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_17_LC_16_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_17_LC_16_24_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ppm_encoder_1.pulses2count_17_LC_16_24_1  (
            .in0(N__45033),
            .in1(N__46900),
            .in2(N__45012),
            .in3(N__48871),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59290),
            .ce(),
            .sr(N__57645));
    defparam \pid_side.pid_prereg_esr_RNIOPAK1_2_LC_17_9_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIOPAK1_2_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIOPAK1_2_LC_17_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIOPAK1_2_LC_17_9_5  (
            .in0(N__49748),
            .in1(N__47731),
            .in2(N__49724),
            .in3(N__47761),
            .lcout(\pid_side.m32_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIKRVH2_5_LC_17_10_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIKRVH2_5_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIKRVH2_5_LC_17_10_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIKRVH2_5_LC_17_10_0  (
            .in0(N__44994),
            .in1(N__47552),
            .in2(N__49618),
            .in3(N__44980),
            .lcout(\pid_side.un1_reset_0_i_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI2NBO1_6_LC_17_10_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI2NBO1_6_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI2NBO1_6_LC_17_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI2NBO1_6_LC_17_10_2  (
            .in0(N__49564),
            .in1(N__49486),
            .in2(N__49541),
            .in3(N__49507),
            .lcout(\pid_side.m26_e_5 ),
            .ltout(\pid_side.m26_e_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI7JSP1_10_LC_17_10_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI7JSP1_10_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI7JSP1_10_LC_17_10_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI7JSP1_10_LC_17_10_3  (
            .in0(N__49927),
            .in1(_gnd_net_),
            .in2(N__44865),
            .in3(N__49966),
            .lcout(\pid_side.pid_prereg_esr_RNI7JSP1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI2NBO1_0_6_LC_17_10_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI2NBO1_0_6_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI2NBO1_0_6_LC_17_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI2NBO1_0_6_LC_17_10_4  (
            .in0(N__49487),
            .in1(N__49537),
            .in2(N__49569),
            .in3(N__49508),
            .lcout(\pid_side.m18_s_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIQEI8_13_LC_17_11_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIQEI8_13_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIQEI8_13_LC_17_11_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \pid_side.pid_prereg_esr_RNIQEI8_13_LC_17_11_0  (
            .in0(N__50014),
            .in1(N__49854),
            .in2(_gnd_net_),
            .in3(N__48084),
            .lcout(\pid_side.N_11_0 ),
            .ltout(\pid_side.N_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNILRSP2_5_LC_17_11_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNILRSP2_5_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNILRSP2_5_LC_17_11_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNILRSP2_5_LC_17_11_1  (
            .in0(N__49611),
            .in1(N__45645),
            .in2(N__44862),
            .in3(N__45694),
            .lcout(\pid_side.pid_prereg_esr_RNILRSP2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIGJDR1_10_LC_17_11_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIGJDR1_10_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIGJDR1_10_LC_17_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIGJDR1_10_LC_17_11_2  (
            .in0(N__49929),
            .in1(N__49968),
            .in2(N__45735),
            .in3(N__47517),
            .lcout(),
            .ltout(\pid_side.pid_prereg_esr_RNIGJDR1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIQBAH2_23_LC_17_11_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIQBAH2_23_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIQBAH2_23_LC_17_11_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIQBAH2_23_LC_17_11_3  (
            .in0(N__48085),
            .in1(N__49664),
            .in2(N__45726),
            .in3(N__50015),
            .lcout(),
            .ltout(\pid_side.pid_prereg_esr_RNIQBAH2Z0Z_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIKNK25_10_LC_17_11_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIKNK25_10_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIKNK25_10_LC_17_11_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIKNK25_10_LC_17_11_4  (
            .in0(N__47592),
            .in1(N__45723),
            .in2(N__45717),
            .in3(N__45661),
            .lcout(),
            .ltout(\pid_side.i19_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIKC058_23_LC_17_11_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIKC058_23_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIKC058_23_LC_17_11_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIKC058_23_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__45714),
            .in2(N__45705),
            .in3(N__47523),
            .lcout(\pid_side.un1_reset_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIEUA9_12_LC_17_11_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIEUA9_12_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIEUA9_12_LC_17_11_6 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \pid_side.pid_prereg_esr_RNIEUA9_12_LC_17_11_6  (
            .in0(N__50016),
            .in1(N__49855),
            .in2(N__49893),
            .in3(N__48086),
            .lcout(\pid_side.pid_prereg_esr_RNIEUA9Z0Z_12 ),
            .ltout(\pid_side.pid_prereg_esr_RNIEUA9Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIF0QB2_10_LC_17_11_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIF0QB2_10_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIF0QB2_10_LC_17_11_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIF0QB2_10_LC_17_11_7  (
            .in0(N__45662),
            .in1(_gnd_net_),
            .in2(N__45648),
            .in3(N__45644),
            .lcout(\pid_side.N_82_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_12_LC_17_12_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_12_LC_17_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_12_LC_17_12_4 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \pid_side.source_pid_1_esr_12_LC_17_12_4  (
            .in0(N__49857),
            .in1(N__48087),
            .in2(N__50028),
            .in3(N__49892),
            .lcout(side_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59137),
            .ce(N__48025),
            .sr(N__47984));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_13_0 .LUT_INIT=16'b0110110001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_13_0  (
            .in0(N__45570),
            .in1(N__46036),
            .in2(N__45878),
            .in3(N__45557),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_0_LC_17_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_0_LC_17_13_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_0_LC_17_13_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \ppm_encoder_1.elevator_0_LC_17_13_1  (
            .in0(N__45429),
            .in1(N__45385),
            .in2(_gnd_net_),
            .in3(N__45874),
            .lcout(\ppm_encoder_1.elevatorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59151),
            .ce(),
            .sr(N__57579));
    defparam \ppm_encoder_1.init_pulses_6_LC_17_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_17_13_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_17_13_5  (
            .in0(N__47468),
            .in1(N__48465),
            .in2(N__47315),
            .in3(N__45849),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59151),
            .ce(),
            .sr(N__57579));
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_17_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_17_13_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICBN01_6_LC_17_13_6  (
            .in0(N__45751),
            .in1(N__48990),
            .in2(_gnd_net_),
            .in3(N__48797),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_13_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_13_7  (
            .in0(N__48798),
            .in1(_gnd_net_),
            .in2(N__49043),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_17_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_17_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__48931),
            .in2(_gnd_net_),
            .in3(N__48637),
            .lcout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ),
            .ltout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_17_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_17_14_1 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNILVE13_0_LC_17_14_1  (
            .in0(N__48640),
            .in1(N__46063),
            .in2(N__45798),
            .in3(N__48286),
            .lcout(\ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_17_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_17_14_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_17_14_2  (
            .in0(N__47871),
            .in1(N__48935),
            .in2(N__48864),
            .in3(N__47912),
            .lcout(\ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_14_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_14_3  (
            .in0(N__48641),
            .in1(N__45783),
            .in2(N__48296),
            .in3(N__47869),
            .lcout(\ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_14_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_14_4  (
            .in0(N__47870),
            .in1(N__48290),
            .in2(N__48865),
            .in3(N__45752),
            .lcout(\ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_14_5 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_14_5  (
            .in0(N__48639),
            .in1(N__48285),
            .in2(N__46071),
            .in3(N__47872),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_17_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_17_14_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_17_14_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_17_14_6  (
            .in0(N__47241),
            .in1(N__46080),
            .in2(N__46074),
            .in3(N__47469),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59164),
            .ce(),
            .sr(N__57588));
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_17_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_17_14_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI65N01_0_LC_17_14_7  (
            .in0(N__48638),
            .in1(_gnd_net_),
            .in2(N__48995),
            .in3(N__46062),
            .lcout(\ppm_encoder_1.un1_init_pulses_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_5_LC_17_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_17_15_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_17_15_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_17_15_0  (
            .in0(N__47456),
            .in1(N__48495),
            .in2(N__47316),
            .in3(N__46017),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59177),
            .ce(),
            .sr(N__57599));
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_15_1  (
            .in0(N__48986),
            .in1(N__45983),
            .in2(_gnd_net_),
            .in3(N__48702),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_17_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_17_15_2 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_17_15_2  (
            .in0(N__45982),
            .in1(_gnd_net_),
            .in2(N__48795),
            .in3(N__48987),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_15_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_15_3  (
            .in0(N__46575),
            .in1(N__45984),
            .in2(N__46446),
            .in3(N__45972),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_7_LC_17_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_17_15_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_17_15_4  (
            .in0(N__47457),
            .in1(N__48441),
            .in2(N__47317),
            .in3(N__45936),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59177),
            .ce(),
            .sr(N__57599));
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_15_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_15_5  (
            .in0(N__48989),
            .in1(N__48709),
            .in2(_gnd_net_),
            .in3(N__45892),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_17_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_17_15_6 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_17_15_6  (
            .in0(N__45893),
            .in1(_gnd_net_),
            .in2(N__48796),
            .in3(N__48988),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_8_LC_17_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_17_16_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_17_16_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_17_16_0  (
            .in0(N__47461),
            .in1(N__48423),
            .in2(N__47346),
            .in3(N__46269),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59193),
            .ce(),
            .sr(N__57606));
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_17_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_17_16_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_17_16_1  (
            .in0(N__46198),
            .in1(N__49021),
            .in2(_gnd_net_),
            .in3(N__48700),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_17_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_17_16_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_17_16_2  (
            .in0(N__48698),
            .in1(_gnd_net_),
            .in2(N__49065),
            .in3(N__46199),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3  (
            .in0(N__46236),
            .in1(N__46436),
            .in2(N__46203),
            .in3(N__46564),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_9_LC_17_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_17_16_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_17_16_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_17_16_4  (
            .in0(N__47462),
            .in1(N__48408),
            .in2(N__47347),
            .in3(N__46173),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59193),
            .ce(),
            .sr(N__57606));
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_17_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_17_16_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_17_16_5  (
            .in0(N__46127),
            .in1(N__49022),
            .in2(_gnd_net_),
            .in3(N__48701),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_17_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_17_16_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_17_16_6  (
            .in0(N__48699),
            .in1(_gnd_net_),
            .in2(N__49066),
            .in3(N__46126),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_16_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_16_7  (
            .in0(N__46113),
            .in1(N__49014),
            .in2(_gnd_net_),
            .in3(N__48697),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_17_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_17_0  (
            .in0(N__46567),
            .in1(N__46112),
            .in2(N__46437),
            .in3(N__46796),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_4_LC_17_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_17_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46824),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59205),
            .ce(N__46781),
            .sr(N__57613));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_17_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_17_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_17_17_2  (
            .in0(N__46407),
            .in1(N__47190),
            .in2(_gnd_net_),
            .in3(N__46716),
            .lcout(),
            .ltout(\ppm_encoder_1.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_17_17_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_17_17_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__46568),
            .in2(N__46692),
            .in3(N__46676),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_17_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_17_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_17_4  (
            .in0(N__49023),
            .in1(N__48815),
            .in2(_gnd_net_),
            .in3(N__47189),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_17_17_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_17_17_5 .LUT_INIT=16'b0110101001101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_17_17_5  (
            .in0(N__47188),
            .in1(N__49024),
            .in2(N__48863),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_17_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_17_18_0 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_17_18_0  (
            .in0(N__47343),
            .in1(N__47464),
            .in2(N__48390),
            .in3(N__46617),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59220),
            .ce(),
            .sr(N__57621));
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_17_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_17_18_1 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINSJT_10_LC_17_18_1  (
            .in0(N__46585),
            .in1(_gnd_net_),
            .in2(N__48861),
            .in3(N__49080),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_17_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_17_18_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_17_18_2  (
            .in0(N__49079),
            .in1(N__48808),
            .in2(_gnd_net_),
            .in3(N__46586),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_18_3 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_18_3  (
            .in0(N__46587),
            .in1(N__46571),
            .in2(N__46455),
            .in3(N__46301),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_11_LC_17_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_17_18_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_17_18_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_17_18_4  (
            .in0(N__47344),
            .in1(N__47465),
            .in2(N__48366),
            .in3(N__47499),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59220),
            .ce(),
            .sr(N__57621));
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_17_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_17_18_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_17_18_5  (
            .in0(N__48313),
            .in1(_gnd_net_),
            .in2(N__48862),
            .in3(N__49081),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_12_LC_17_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_17_18_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_17_18_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_17_18_7  (
            .in0(N__47463),
            .in1(N__47345),
            .in2(N__48345),
            .in3(N__47199),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59220),
            .ce(),
            .sr(N__57621));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_19_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_19_0  (
            .in0(N__47126),
            .in1(N__47040),
            .in2(_gnd_net_),
            .in3(N__47004),
            .lcout(\ppm_encoder_1.N_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_17_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_17_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_17_19_2  (
            .in0(N__51427),
            .in1(N__46968),
            .in2(_gnd_net_),
            .in3(N__46959),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_1_LC_17_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_17_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_17_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_1_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56895),
            .lcout(\pid_front.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59268),
            .ce(N__49376),
            .sr(N__57637));
    defparam \ppm_encoder_1.pulses2count_15_LC_17_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_15_LC_17_22_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_15_LC_17_22_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_15_LC_17_22_1  (
            .in0(N__47905),
            .in1(N__46865),
            .in2(N__46906),
            .in3(N__48873),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59282),
            .ce(),
            .sr(N__57642));
    defparam \pid_front.error_d_reg_prev_esr_11_LC_17_23_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_17_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_17_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_11_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56822),
            .lcout(\pid_front.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59291),
            .ce(N__49375),
            .sr(N__57646));
    defparam \pid_alt.state_RNICP2N1_0_LC_18_6_0 .C_ON=1'b0;
    defparam \pid_alt.state_RNICP2N1_0_LC_18_6_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNICP2N1_0_LC_18_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNICP2N1_0_LC_18_6_0  (
            .in0(_gnd_net_),
            .in1(N__47796),
            .in2(_gnd_net_),
            .in3(N__58319),
            .lcout(\pid_alt.N_664_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_0_LC_18_9_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_0_LC_18_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_0_LC_18_9_1 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_side.pid_prereg_0_LC_18_9_1  (
            .in0(N__47618),
            .in1(N__50940),
            .in2(N__53511),
            .in3(N__47762),
            .lcout(\pid_side.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59115),
            .ce(),
            .sr(N__57555));
    defparam \pid_side.pid_prereg_1_LC_18_9_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_1_LC_18_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_1_LC_18_9_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pid_side.pid_prereg_1_LC_18_9_2  (
            .in0(N__49266),
            .in1(N__50832),
            .in2(N__47741),
            .in3(N__47619),
            .lcout(\pid_side.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59115),
            .ce(),
            .sr(N__57555));
    defparam \pid_side.state_0_LC_18_9_4 .C_ON=1'b0;
    defparam \pid_side.state_0_LC_18_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_0_LC_18_9_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_side.state_0_LC_18_9_4  (
            .in0(N__47711),
            .in1(N__47617),
            .in2(_gnd_net_),
            .in3(N__47554),
            .lcout(\pid_side.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59115),
            .ce(),
            .sr(N__57555));
    defparam \pid_side.state_RNINK4U_0_LC_18_9_5 .C_ON=1'b0;
    defparam \pid_side.state_RNINK4U_0_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNINK4U_0_LC_18_9_5 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \pid_side.state_RNINK4U_0_LC_18_9_5  (
            .in0(N__47553),
            .in1(N__47710),
            .in2(N__47622),
            .in3(N__57830),
            .lcout(\pid_side.state_RNINK4UZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_1_LC_18_9_7 .C_ON=1'b0;
    defparam \pid_side.state_1_LC_18_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_1_LC_18_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.state_1_LC_18_9_7  (
            .in0(N__47620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59115),
            .ce(),
            .sr(N__57555));
    defparam \pid_side.pid_prereg_esr_RNIU5CG_10_LC_18_10_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIU5CG_10_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIU5CG_10_LC_18_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIU5CG_10_LC_18_10_0  (
            .in0(N__49926),
            .in1(N__49965),
            .in2(N__49694),
            .in3(N__49882),
            .lcout(\pid_side.m18_s_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNICPBG_23_LC_18_10_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNICPBG_23_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNICPBG_23_LC_18_10_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \pid_side.pid_prereg_esr_RNICPBG_23_LC_18_10_3  (
            .in0(N__57829),
            .in1(N__47551),
            .in2(_gnd_net_),
            .in3(N__50024),
            .lcout(\pid_side.un1_reset_0_i_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI90H1_12_LC_18_10_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI90H1_12_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI90H1_12_LC_18_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI90H1_12_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__49881),
            .in2(_gnd_net_),
            .in3(N__49842),
            .lcout(\pid_side.m26_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI2MA2_14_LC_18_10_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI2MA2_14_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI2MA2_14_LC_18_10_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI2MA2_14_LC_18_10_7  (
            .in0(N__49821),
            .in1(N__50046),
            .in2(_gnd_net_),
            .in3(N__49806),
            .lcout(\pid_side.m9_e_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_11_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_11_0  (
            .in0(N__50085),
            .in1(N__49794),
            .in2(N__49770),
            .in3(N__49782),
            .lcout(),
            .ltout(\pid_side.m9_e_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIFB07_20_LC_18_11_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIFB07_20_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIFB07_20_LC_18_11_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIFB07_20_LC_18_11_1  (
            .in0(N__48096),
            .in1(N__50070),
            .in2(N__48090),
            .in3(N__50058),
            .lcout(\pid_side.pid_prereg_esr_RNIFB07Z0Z_20 ),
            .ltout(\pid_side.pid_prereg_esr_RNIFB07Z0Z_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_13_LC_18_11_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_13_LC_18_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_13_LC_18_11_2 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \pid_side.source_pid_1_esr_13_LC_18_11_2  (
            .in0(N__50020),
            .in1(_gnd_net_),
            .in2(N__48069),
            .in3(N__49856),
            .lcout(side_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59138),
            .ce(N__48035),
            .sr(N__47985));
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_18_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_18_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIC08S_3_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__47945),
            .in2(_gnd_net_),
            .in3(N__57858),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_14_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_14_0  (
            .in0(N__47913),
            .in1(N__48999),
            .in2(_gnd_net_),
            .in3(N__48823),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_18_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_18_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_18_14_1  (
            .in0(N__48825),
            .in1(N__47873),
            .in2(N__48297),
            .in3(N__47847),
            .lcout(\ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_18_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_18_14_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_18_14_2  (
            .in0(N__47823),
            .in1(N__48996),
            .in2(_gnd_net_),
            .in3(N__48819),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_18_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_18_14_3 .LUT_INIT=16'b1101110011011110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_18_14_3  (
            .in0(N__48824),
            .in1(N__57895),
            .in2(N__51400),
            .in3(N__49013),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59178),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_14_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_14_4  (
            .in0(N__48326),
            .in1(N__48998),
            .in2(_gnd_net_),
            .in3(N__48821),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_18_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_18_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_18_14_5  (
            .in0(N__48822),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48292),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_18_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_18_14_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_18_14_6  (
            .in0(N__48240),
            .in1(N__48997),
            .in2(_gnd_net_),
            .in3(N__48820),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_18_15_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_18_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__48216),
            .in2(N__48204),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_15_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__48195),
            .in2(_gnd_net_),
            .in3(N__48177),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_15_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__48174),
            .in2(N__48168),
            .in3(N__48141),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_15_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__48138),
            .in2(_gnd_net_),
            .in3(N__48120),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_15_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__48117),
            .in2(_gnd_net_),
            .in3(N__48099),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_15_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__48501),
            .in2(_gnd_net_),
            .in3(N__48489),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_15_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__48486),
            .in2(N__48480),
            .in3(N__48453),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_15_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48450),
            .in3(N__48435),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_16_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__48432),
            .in2(_gnd_net_),
            .in3(N__48417),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_16_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__48414),
            .in2(_gnd_net_),
            .in3(N__48402),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_16_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__48399),
            .in2(_gnd_net_),
            .in3(N__48378),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_16_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__48375),
            .in2(_gnd_net_),
            .in3(N__48354),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_16_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__48351),
            .in2(_gnd_net_),
            .in3(N__48333),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_16_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__49254),
            .in2(N__49245),
            .in3(N__49221),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_16_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__49218),
            .in2(_gnd_net_),
            .in3(N__49194),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_16_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__49191),
            .in2(_gnd_net_),
            .in3(N__49170),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__49167),
            .in2(_gnd_net_),
            .in3(N__49143),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__49140),
            .in2(_gnd_net_),
            .in3(N__49116),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_17_2 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_17_2  (
            .in0(N__49112),
            .in1(N__49060),
            .in2(N__48872),
            .in3(N__48522),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_18_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_18_17_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__48507),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_18_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_18_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_18_18_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__52484),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59236),
            .ce(N__50297),
            .sr(N__57627));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_18_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_18_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_18_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53224),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59236),
            .ce(N__50297),
            .sr(N__57627));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_18_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_18_18_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_18_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52374),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59236),
            .ce(N__50297),
            .sr(N__57627));
    defparam \pid_front.pid_prereg_0_LC_18_20_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_0_LC_18_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_0_LC_18_20_4 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_front.pid_prereg_0_LC_18_20_4  (
            .in0(N__50508),
            .in1(N__49461),
            .in2(N__56940),
            .in3(N__49423),
            .lcout(\pid_front.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59269),
            .ce(),
            .sr(N__57638));
    defparam \pid_front.error_d_reg_prev_esr_18_LC_18_22_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_18_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_18_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_18_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59573),
            .lcout(\pid_front.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59292),
            .ce(N__49377),
            .sr(N__57647));
    defparam \pid_front.error_d_reg_esr_2_LC_18_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_2_LC_18_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_2_LC_18_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_2_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49311),
            .lcout(\pid_front.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59302),
            .ce(N__58455),
            .sr(N__58179));
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6.C_ON=1'b0;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57827),
            .lcout(GB_BUFFER_reset_system_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_1_LC_20_8_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_20_8_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_20_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_1_LC_20_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53436),
            .lcout(\pid_side.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59125),
            .ce(N__57948),
            .sr(N__57564));
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_9_0 .C_ON=1'b1;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_0_LC_20_9_0  (
            .in0(_gnd_net_),
            .in1(N__50936),
            .in2(N__53510),
            .in3(N__53509),
            .lcout(\pid_side.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(bfn_20_9_0_),
            .carryout(\pid_side.un1_pid_prereg_cry_0 ),
            .clk(N__59140),
            .ce(N__57950),
            .sr(N__57574));
    defparam \pid_side.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_20_9_1 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_20_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_0_THRU_LUT4_0_LC_20_9_1  (
            .in0(_gnd_net_),
            .in1(N__50828),
            .in2(_gnd_net_),
            .in3(N__49257),
            .lcout(\pid_side.un1_pid_prereg_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_0 ),
            .carryout(\pid_side.un1_pid_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_2_LC_20_9_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_2_LC_20_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_2_LC_20_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_2_LC_20_9_2  (
            .in0(_gnd_net_),
            .in1(N__50814),
            .in2(N__50967),
            .in3(N__49731),
            .lcout(\pid_side.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_1 ),
            .carryout(\pid_side.un1_pid_prereg_cry_0_0 ),
            .clk(N__59140),
            .ce(N__57950),
            .sr(N__57574));
    defparam \pid_side.pid_prereg_esr_3_LC_20_9_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_3_LC_20_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_3_LC_20_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_3_LC_20_9_3  (
            .in0(_gnd_net_),
            .in1(N__50925),
            .in2(N__53043),
            .in3(N__49701),
            .lcout(\pid_side.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_0_0 ),
            .carryout(\pid_side.un1_pid_prereg_cry_1_0 ),
            .clk(N__59140),
            .ce(N__57950),
            .sr(N__57574));
    defparam \pid_side.pid_prereg_esr_4_LC_20_9_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_4_LC_20_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_4_LC_20_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_4_LC_20_9_4  (
            .in0(_gnd_net_),
            .in1(N__53655),
            .in2(N__52803),
            .in3(N__49623),
            .lcout(\pid_side.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_1_0 ),
            .carryout(\pid_side.un1_pid_prereg_cry_2 ),
            .clk(N__59140),
            .ce(N__57950),
            .sr(N__57574));
    defparam \pid_side.pid_prereg_esr_5_LC_20_9_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_5_LC_20_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_5_LC_20_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_5_LC_20_9_5  (
            .in0(_gnd_net_),
            .in1(N__52833),
            .in2(N__52857),
            .in3(N__49572),
            .lcout(\pid_side.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_2 ),
            .carryout(\pid_side.un1_pid_prereg_cry_3 ),
            .clk(N__59140),
            .ce(N__57950),
            .sr(N__57574));
    defparam \pid_side.pid_prereg_esr_6_LC_20_9_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_6_LC_20_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_6_LC_20_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_6_LC_20_9_6  (
            .in0(_gnd_net_),
            .in1(N__52877),
            .in2(N__50847),
            .in3(N__49545),
            .lcout(\pid_side.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_3 ),
            .carryout(\pid_side.un1_pid_prereg_cry_4 ),
            .clk(N__59140),
            .ce(N__57950),
            .sr(N__57574));
    defparam \pid_side.pid_prereg_esr_7_LC_20_9_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_7_LC_20_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_7_LC_20_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_7_LC_20_9_7  (
            .in0(_gnd_net_),
            .in1(N__54633),
            .in2(N__54612),
            .in3(N__49512),
            .lcout(\pid_side.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_4 ),
            .carryout(\pid_side.un1_pid_prereg_cry_5 ),
            .clk(N__59140),
            .ce(N__57950),
            .sr(N__57574));
    defparam \pid_side.pid_prereg_esr_8_LC_20_10_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_8_LC_20_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_8_LC_20_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_8_LC_20_10_0  (
            .in0(_gnd_net_),
            .in1(N__54942),
            .in2(N__54591),
            .in3(N__49491),
            .lcout(\pid_side.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(bfn_20_10_0_),
            .carryout(\pid_side.un1_pid_prereg_cry_6 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_9_LC_20_10_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_9_LC_20_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_9_LC_20_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_9_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__53703),
            .in2(N__53727),
            .in3(N__49464),
            .lcout(\pid_side.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_6 ),
            .carryout(\pid_side.un1_pid_prereg_cry_7 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_10_LC_20_10_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_10_LC_20_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_10_LC_20_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_10_LC_20_10_2  (
            .in0(_gnd_net_),
            .in1(N__51078),
            .in2(N__53757),
            .in3(N__49932),
            .lcout(\pid_side.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_7 ),
            .carryout(\pid_side.un1_pid_prereg_cry_8 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_11_LC_20_10_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_11_LC_20_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_11_LC_20_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_11_LC_20_10_3  (
            .in0(_gnd_net_),
            .in1(N__51063),
            .in2(N__51183),
            .in3(N__49896),
            .lcout(\pid_side.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_8 ),
            .carryout(\pid_side.un1_pid_prereg_cry_9 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_12_LC_20_10_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_12_LC_20_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_12_LC_20_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_12_LC_20_10_4  (
            .in0(_gnd_net_),
            .in1(N__51195),
            .in2(N__51135),
            .in3(N__49860),
            .lcout(\pid_side.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_9 ),
            .carryout(\pid_side.un1_pid_prereg_cry_10 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_13_LC_20_10_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_13_LC_20_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_13_LC_20_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_13_LC_20_10_5  (
            .in0(_gnd_net_),
            .in1(N__51102),
            .in2(N__51122),
            .in3(N__49824),
            .lcout(\pid_side.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_10 ),
            .carryout(\pid_side.un1_pid_prereg_cry_11 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_14_LC_20_10_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_14_LC_20_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_14_LC_20_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_14_LC_20_10_6  (
            .in0(_gnd_net_),
            .in1(N__51093),
            .in2(N__51003),
            .in3(N__49809),
            .lcout(\pid_side.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_11 ),
            .carryout(\pid_side.un1_pid_prereg_cry_12 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_15_LC_20_10_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_15_LC_20_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_15_LC_20_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_15_LC_20_10_7  (
            .in0(_gnd_net_),
            .in1(N__51057),
            .in2(N__50916),
            .in3(N__49797),
            .lcout(\pid_side.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_12 ),
            .carryout(\pid_side.un1_pid_prereg_cry_13 ),
            .clk(N__59153),
            .ce(N__57951),
            .sr(N__57581));
    defparam \pid_side.pid_prereg_esr_16_LC_20_11_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_16_LC_20_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_16_LC_20_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_16_LC_20_11_0  (
            .in0(_gnd_net_),
            .in1(N__51084),
            .in2(N__50181),
            .in3(N__49785),
            .lcout(\pid_side.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(bfn_20_11_0_),
            .carryout(\pid_side.un1_pid_prereg_cry_14 ),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.pid_prereg_esr_17_LC_20_11_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_17_LC_20_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_17_LC_20_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_17_LC_20_11_1  (
            .in0(_gnd_net_),
            .in1(N__49974),
            .in2(N__50106),
            .in3(N__49773),
            .lcout(\pid_side.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_14 ),
            .carryout(\pid_side.un1_pid_prereg_cry_15 ),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.pid_prereg_esr_18_LC_20_11_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_18_LC_20_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_18_LC_20_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_18_LC_20_11_2  (
            .in0(_gnd_net_),
            .in1(N__50157),
            .in2(N__52923),
            .in3(N__49758),
            .lcout(\pid_side.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_15 ),
            .carryout(\pid_side.un1_pid_prereg_cry_16 ),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.pid_prereg_esr_19_LC_20_11_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_19_LC_20_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_19_LC_20_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_19_LC_20_11_3  (
            .in0(_gnd_net_),
            .in1(N__50172),
            .in2(N__53553),
            .in3(N__50073),
            .lcout(\pid_side.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_16 ),
            .carryout(\pid_side.un1_pid_prereg_cry_17 ),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.pid_prereg_esr_20_LC_20_11_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_20_LC_20_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_20_LC_20_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_20_LC_20_11_4  (
            .in0(_gnd_net_),
            .in1(N__49980),
            .in2(N__50166),
            .in3(N__50061),
            .lcout(\pid_side.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_17 ),
            .carryout(\pid_side.un1_pid_prereg_cry_18 ),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.pid_prereg_esr_21_LC_20_11_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_21_LC_20_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_21_LC_20_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_21_LC_20_11_5  (
            .in0(_gnd_net_),
            .in1(N__50094),
            .in2(N__50196),
            .in3(N__50049),
            .lcout(\pid_side.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_18 ),
            .carryout(\pid_side.un1_pid_prereg_cry_19 ),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.pid_prereg_esr_22_LC_20_11_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_22_LC_20_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_22_LC_20_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_22_LC_20_11_6  (
            .in0(_gnd_net_),
            .in1(N__50274),
            .in2(N__51204),
            .in3(N__50034),
            .lcout(\pid_side.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_19 ),
            .carryout(\pid_side.un1_pid_prereg_cry_20 ),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.pid_prereg_esr_23_LC_20_11_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_23_LC_20_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_23_LC_20_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.pid_prereg_esr_23_LC_20_11_7  (
            .in0(_gnd_net_),
            .in1(N__50265),
            .in2(_gnd_net_),
            .in3(N__50031),
            .lcout(\pid_side.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59166),
            .ce(N__57952),
            .sr(N__57590));
    defparam \pid_side.error_d_reg_prev_esr_RNILHF23_18_LC_20_12_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNILHF23_18_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNILHF23_18_LC_20_12_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNILHF23_18_LC_20_12_0  (
            .in0(N__51833),
            .in1(N__51227),
            .in2(N__53991),
            .in3(N__52956),
            .lcout(\pid_side.error_d_reg_prev_esr_RNILHF23Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIJV5H1_15_LC_20_12_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIJV5H1_15_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIJV5H1_15_LC_20_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIJV5H1_15_LC_20_12_3  (
            .in0(N__50134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50117),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIJV5H1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_12_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_12_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_12_4  (
            .in0(N__54378),
            .in1(N__52989),
            .in2(_gnd_net_),
            .in3(N__54813),
            .lcout(\pid_side.un1_pid_prereg_30 ),
            .ltout(\pid_side.un1_pid_prereg_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0PB23_14_LC_20_12_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0PB23_14_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0PB23_14_LC_20_12_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0PB23_14_LC_20_12_5  (
            .in0(N__50135),
            .in1(N__50994),
            .in2(N__50184),
            .in3(N__52974),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI0PB23Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI4UC23_17_LC_20_12_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI4UC23_17_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI4UC23_17_LC_20_12_6 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI4UC23_17_LC_20_12_6  (
            .in0(N__52896),
            .in1(N__52954),
            .in2(N__51228),
            .in3(N__54102),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI4UC23Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI5I6H1_18_LC_20_12_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5I6H1_18_LC_20_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5I6H1_18_LC_20_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5I6H1_18_LC_20_12_7  (
            .in0(N__52955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51226),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI5I6H1Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIP56H1_16_LC_20_13_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIP56H1_16_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIP56H1_16_LC_20_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIP56H1_16_LC_20_13_2  (
            .in0(N__54121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52934),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIP56H1Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_16_LC_20_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_20_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_20_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_16_LC_20_13_3  (
            .in0(N__56628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59195),
            .ce(N__57956),
            .sr(N__57607));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_20_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_20_13_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_20_13_4  (
            .in0(N__54179),
            .in1(N__50144),
            .in2(_gnd_net_),
            .in3(N__56626),
            .lcout(\pid_side.un1_pid_prereg_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_20_13_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_20_13_5 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_20_13_5  (
            .in0(N__56627),
            .in1(_gnd_net_),
            .in2(N__50148),
            .in3(N__54180),
            .lcout(\pid_side.un1_pid_prereg_36 ),
            .ltout(\pid_side.un1_pid_prereg_36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIC5C23_15_LC_20_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIC5C23_15_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIC5C23_15_LC_20_13_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIC5C23_15_LC_20_13_6  (
            .in0(N__54122),
            .in1(N__50136),
            .in2(N__50121),
            .in3(N__50118),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIC5C23Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI89K23_19_LC_20_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI89K23_19_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI89K23_19_LC_20_14_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI89K23_19_LC_20_14_1  (
            .in0(N__54029),
            .in1(N__53983),
            .in2(N__51834),
            .in3(N__53980),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI89K23Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIGJM23_20_LC_20_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIGJM23_20_LC_20_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIGJM23_20_LC_20_14_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIGJM23_20_LC_20_14_2  (
            .in0(N__54028),
            .in1(N__53979),
            .in2(N__54035),
            .in3(N__53978),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIGJM23Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNO_0_23_LC_20_14_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNO_0_23_LC_20_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNO_0_23_LC_20_14_5 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_side.pid_prereg_esr_RNO_0_23_LC_20_14_5  (
            .in0(N__54030),
            .in1(N__53981),
            .in2(N__54036),
            .in3(N__53982),
            .lcout(\pid_side.un1_pid_prereg_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_20_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_20_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_20_14_6  (
            .in0(N__51365),
            .in1(N__50256),
            .in2(_gnd_net_),
            .in3(N__50244),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIGV8H1_19_LC_20_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIGV8H1_19_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIGV8H1_19_LC_20_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIGV8H1_19_LC_20_15_3  (
            .in0(_gnd_net_),
            .in1(N__53974),
            .in2(_gnd_net_),
            .in3(N__51826),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIGV8H1Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_20_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_20_16_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_20_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_20_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56285),
            .lcout(side_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59238),
            .ce(N__51810),
            .sr(N__57628));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_20_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_20_16_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_20_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_20_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56132),
            .lcout(side_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59238),
            .ce(N__51810),
            .sr(N__57628));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_20_16_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_20_16_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_20_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_20_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56507),
            .lcout(side_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59238),
            .ce(N__51810),
            .sr(N__57628));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_20_16_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_20_16_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_20_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_20_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53397),
            .lcout(side_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59238),
            .ce(N__51810),
            .sr(N__57628));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_20_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_20_16_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_20_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_20_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55926),
            .lcout(side_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59238),
            .ce(N__51810),
            .sr(N__57628));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_20_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_20_16_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_20_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_20_16_6  (
            .in0(N__55749),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(side_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59238),
            .ce(N__51810),
            .sr(N__57628));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_20_16_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_20_16_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_20_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_20_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55574),
            .lcout(side_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59238),
            .ce(N__51810),
            .sr(N__57628));
    defparam \pid_side.error_axb_1_LC_20_17_0 .C_ON=1'b0;
    defparam \pid_side.error_axb_1_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_1_LC_20_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_1_LC_20_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50409),
            .lcout(\pid_side.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_20_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_20_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_20_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50780),
            .lcout(drone_H_disp_side_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59254),
            .ce(N__50298),
            .sr(N__57633));
    defparam \pid_side.error_axb_2_LC_20_17_2 .C_ON=1'b0;
    defparam \pid_side.error_axb_2_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_2_LC_20_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_2_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50310),
            .lcout(\pid_side.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_20_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_20_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_20_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50402),
            .lcout(drone_H_disp_side_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59254),
            .ce(N__50298),
            .sr(N__57633));
    defparam \pid_side.error_axb_3_LC_20_17_4 .C_ON=1'b0;
    defparam \pid_side.error_axb_3_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_3_LC_20_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_3_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50304),
            .lcout(\pid_side.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_20_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_20_17_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_20_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_20_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52709),
            .lcout(drone_H_disp_side_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59254),
            .ce(N__50298),
            .sr(N__57633));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_20_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_20_17_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_20_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_20_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52307),
            .lcout(drone_H_disp_side_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59254),
            .ce(N__50298),
            .sr(N__57633));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_20_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_20_17_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_20_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_20_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52605),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59254),
            .ce(N__50298),
            .sr(N__57633));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_20_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_20_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_20_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50703),
            .lcout(drone_H_disp_front_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_20_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_20_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_20_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50781),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59271),
            .ce(N__50696),
            .sr(N__57639));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_20_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_20_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_20_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52406),
            .lcout(drone_H_disp_side_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_20_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_20_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_20_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50649),
            .lcout(drone_H_disp_side_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_20_18_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_20_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_20_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50643),
            .lcout(drone_H_disp_side_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_20_18_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_20_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_20_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50634),
            .lcout(drone_H_disp_side_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_20_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_20_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52236),
            .lcout(drone_H_disp_side_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_1_LC_20_19_2 .C_ON=1'b0;
    defparam \pid_front.state_1_LC_20_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_1_LC_20_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.state_1_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50505),
            .lcout(\pid_front.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59284),
            .ce(),
            .sr(N__57643));
    defparam \pid_front.pid_prereg_1_LC_20_19_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_1_LC_20_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_1_LC_20_19_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pid_front.pid_prereg_1_LC_20_19_4  (
            .in0(N__50544),
            .in1(N__50529),
            .in2(N__50434),
            .in3(N__50506),
            .lcout(\pid_front.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59284),
            .ce(),
            .sr(N__57643));
    defparam \pid_side.error_axb_8_l_ofx_LC_20_19_5 .C_ON=1'b0;
    defparam \pid_side.error_axb_8_l_ofx_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_8_l_ofx_LC_20_19_5 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_side.error_axb_8_l_ofx_LC_20_19_5  (
            .in0(N__52614),
            .in1(_gnd_net_),
            .in2(N__50892),
            .in3(N__52502),
            .lcout(\pid_side.error_axb_8_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_7_LC_20_19_6 .C_ON=1'b0;
    defparam \pid_side.error_axb_7_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_7_LC_20_19_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_axb_7_LC_20_19_6  (
            .in0(_gnd_net_),
            .in1(N__50888),
            .in2(_gnd_net_),
            .in3(N__52613),
            .lcout(\pid_side.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_20_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_20_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_20_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52501),
            .lcout(drone_H_disp_side_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_3_LC_20_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_3_LC_20_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_3_LC_20_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_3_LC_20_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50877),
            .lcout(\pid_front.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59315),
            .ce(N__58494),
            .sr(N__58180));
    defparam \pid_side.error_p_reg_esr_RNI5QI23_5_LC_21_7_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5QI23_5_LC_21_7_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5QI23_5_LC_21_7_0 .LUT_INIT=16'b0011100100111001;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5QI23_5_LC_21_7_0  (
            .in0(N__53784),
            .in1(N__54894),
            .in2(N__53823),
            .in3(N__52878),
            .lcout(\pid_side.error_p_reg_esr_RNI5QI23Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_5_LC_21_7_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_21_7_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_21_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_5_LC_21_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54753),
            .lcout(\pid_side.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59126),
            .ce(N__57949),
            .sr(N__57565));
    defparam \pid_side.error_d_reg_esr_RNI5QKD1_1_LC_21_9_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI5QKD1_1_LC_21_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI5QKD1_1_LC_21_9_0 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \pid_side.error_d_reg_esr_RNI5QKD1_1_LC_21_9_0  (
            .in0(N__53022),
            .in1(N__50952),
            .in2(N__53435),
            .in3(N__50807),
            .lcout(\pid_side.un1_pid_prereg_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISH6J_0_LC_21_9_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISH6J_0_LC_21_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISH6J_0_LC_21_9_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pid_side.error_p_reg_esr_RNISH6J_0_LC_21_9_1  (
            .in0(N__50950),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53020),
            .lcout(),
            .ltout(\pid_side.error_p_reg_esr_RNISH6JZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNIFP9R2_1_LC_21_9_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNIFP9R2_1_LC_21_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNIFP9R2_1_LC_21_9_2 .LUT_INIT=16'b1010000011111010;
    LogicCell40 \pid_side.error_d_reg_esr_RNIFP9R2_1_LC_21_9_2  (
            .in0(N__53431),
            .in1(N__50966),
            .in2(N__50817),
            .in3(N__50808),
            .lcout(\pid_side.error_d_reg_esr_RNIFP9R2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIUJ6J_0_1_LC_21_9_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIUJ6J_0_1_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIUJ6J_0_1_LC_21_9_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIUJ6J_0_1_LC_21_9_3  (
            .in0(_gnd_net_),
            .in1(N__54257),
            .in2(_gnd_net_),
            .in3(N__50978),
            .lcout(\pid_side.N_1546_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIUJ6J_1_LC_21_9_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIUJ6J_1_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIUJ6J_1_LC_21_9_4 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIUJ6J_1_LC_21_9_4  (
            .in0(N__50979),
            .in1(_gnd_net_),
            .in2(N__54261),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1 ),
            .ltout(\pid_side.error_p_reg_esr_RNIUJ6JZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIAVKD1_0_1_LC_21_9_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIAVKD1_0_1_LC_21_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIAVKD1_0_1_LC_21_9_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIAVKD1_0_1_LC_21_9_5  (
            .in0(_gnd_net_),
            .in1(N__53645),
            .in2(N__50970),
            .in3(_gnd_net_),
            .lcout(\pid_side.un1_pid_prereg ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISH6J_0_0_LC_21_9_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISH6J_0_0_LC_21_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISH6J_0_0_LC_21_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_p_reg_esr_RNISH6J_0_0_LC_21_9_6  (
            .in0(N__53021),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50951),
            .lcout(\pid_side.un1_pid_prereg_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIAVKD1_1_LC_21_9_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIAVKD1_1_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIAVKD1_1_LC_21_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIAVKD1_1_LC_21_9_7  (
            .in0(_gnd_net_),
            .in1(N__53646),
            .in2(_gnd_net_),
            .in3(N__53054),
            .lcout(\pid_side.error_p_reg_esr_RNIAVKD1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_21_10_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_21_10_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_21_10_1  (
            .in0(N__54512),
            .in1(N__50900),
            .in2(_gnd_net_),
            .in3(N__55102),
            .lcout(\pid_side.un1_pid_prereg_18 ),
            .ltout(\pid_side.un1_pid_prereg_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_10_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_10_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50919),
            .in3(N__51048),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_10_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_10_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_10_3  (
            .in0(N__54513),
            .in1(N__50901),
            .in2(_gnd_net_),
            .in3(N__55103),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI4NA21_0_12_LC_21_10_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI4NA21_0_12_LC_21_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI4NA21_0_12_LC_21_10_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI4NA21_0_12_LC_21_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50904),
            .in3(N__51523),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI4NA21_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_13_LC_21_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_21_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_21_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_13_LC_21_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55104),
            .lcout(\pid_side.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59167),
            .ce(N__57953),
            .sr(N__57591));
    defparam \pid_side.error_d_reg_prev_esr_RNI4NA21_12_LC_21_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI4NA21_12_LC_21_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI4NA21_12_LC_21_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI4NA21_12_LC_21_10_6  (
            .in0(_gnd_net_),
            .in1(N__51026),
            .in2(_gnd_net_),
            .in3(N__51524),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI4NA21Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_21_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_21_10_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_21_10_7  (
            .in0(N__54431),
            .in1(N__53574),
            .in2(_gnd_net_),
            .in3(N__55169),
            .lcout(\pid_side.un1_pid_prereg_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIDP5H1_14_LC_21_11_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIDP5H1_14_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIDP5H1_14_LC_21_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIDP5H1_14_LC_21_11_0  (
            .in0(_gnd_net_),
            .in1(N__50993),
            .in2(_gnd_net_),
            .in3(N__52970),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIDP5H1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNIKMFP2_10_LC_21_11_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNIKMFP2_10_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNIKMFP2_10_LC_21_11_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_esr_RNIKMFP2_10_LC_21_11_2  (
            .in0(N__55078),
            .in1(N__51072),
            .in2(N__53756),
            .in3(N__52997),
            .lcout(\pid_side.error_d_reg_esr_RNIKMFP2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUQN9_0_10_LC_21_11_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUQN9_0_10_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUQN9_0_10_LC_21_11_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUQN9_0_10_LC_21_11_3  (
            .in0(_gnd_net_),
            .in1(N__54401),
            .in2(_gnd_net_),
            .in3(N__53538),
            .lcout(\pid_side.N_1582_i ),
            .ltout(\pid_side.N_1582_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI104E2_10_LC_21_11_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI104E2_10_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI104E2_10_LC_21_11_4 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_d_reg_esr_RNI104E2_10_LC_21_11_4  (
            .in0(N__55079),
            .in1(N__51179),
            .in2(N__51066),
            .in3(N__52998),
            .lcout(\pid_side.error_d_reg_esr_RNI104E2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKCB23_13_LC_21_11_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKCB23_13_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKCB23_13_LC_21_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKCB23_13_LC_21_11_6  (
            .in0(N__51047),
            .in1(N__50992),
            .in2(N__51015),
            .in3(N__52969),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIKCB23Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBAGJ2_12_LC_21_11_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBAGJ2_12_LC_21_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBAGJ2_12_LC_21_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBAGJ2_12_LC_21_11_7  (
            .in0(N__51525),
            .in1(N__51046),
            .in2(N__51033),
            .in3(N__51011),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIBAGJ2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_21_12_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_21_12_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_21_12_0  (
            .in0(N__54377),
            .in1(N__52985),
            .in2(_gnd_net_),
            .in3(N__54808),
            .lcout(\pid_side.un1_pid_prereg_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIO9BH1_20_LC_21_12_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIO9BH1_20_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIO9BH1_20_LC_21_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIO9BH1_20_LC_21_12_2  (
            .in0(_gnd_net_),
            .in1(N__53990),
            .in2(_gnd_net_),
            .in3(N__54034),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIO9BH1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNILJFJ2_12_LC_21_12_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNILJFJ2_12_LC_21_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNILJFJ2_12_LC_21_12_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNILJFJ2_12_LC_21_12_3  (
            .in0(N__51548),
            .in1(N__51144),
            .in2(N__51165),
            .in3(N__51555),
            .lcout(\pid_side.error_d_reg_prev_esr_RNILJFJ2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUQN9_10_LC_21_12_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUQN9_10_LC_21_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUQN9_10_LC_21_12_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUQN9_10_LC_21_12_4  (
            .in0(N__53537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54405),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIUQN9Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQCA21_0_10_LC_21_12_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQCA21_0_10_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQCA21_0_10_LC_21_12_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQCA21_0_10_LC_21_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51186),
            .in3(N__51158),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQCA21_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_12_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_12_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_12_6  (
            .in0(N__51506),
            .in1(N__51483),
            .in2(_gnd_net_),
            .in3(N__54870),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQCA21_10_LC_21_12_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQCA21_10_LC_21_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQCA21_10_LC_21_12_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQCA21_10_LC_21_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51147),
            .in3(N__51143),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQCA21Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_12_LC_21_13_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_21_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_21_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_12_LC_21_13_0  (
            .in0(N__54711),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59207),
            .ce(N__57958),
            .sr(N__57614));
    defparam \pid_side.error_d_reg_prev_esr_RNI2VN9_0_12_LC_21_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2VN9_0_12_LC_21_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2VN9_0_12_LC_21_13_1 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2VN9_0_12_LC_21_13_1  (
            .in0(N__51537),
            .in1(_gnd_net_),
            .in2(N__54657),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\pid_side.N_1590_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNIVTFJ2_12_LC_21_13_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNIVTFJ2_12_LC_21_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNIVTFJ2_12_LC_21_13_2 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_d_reg_esr_RNIVTFJ2_12_LC_21_13_2  (
            .in0(N__54710),
            .in1(N__51123),
            .in2(N__51105),
            .in3(N__51549),
            .lcout(\pid_side.error_d_reg_esr_RNIVTFJ2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVKIO_12_LC_21_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVKIO_12_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVKIO_12_LC_21_13_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVKIO_12_LC_21_13_3  (
            .in0(N__51536),
            .in1(_gnd_net_),
            .in2(N__54656),
            .in3(N__54709),
            .lcout(\pid_side.un1_pid_prereg_107_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_13_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_13_4  (
            .in0(N__51482),
            .in1(N__51507),
            .in2(_gnd_net_),
            .in3(N__54868),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHIOZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2VN9_12_LC_21_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2VN9_12_LC_21_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2VN9_12_LC_21_13_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2VN9_12_LC_21_13_6  (
            .in0(_gnd_net_),
            .in1(N__54649),
            .in2(_gnd_net_),
            .in3(N__51535),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2VN9Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_13_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_11_LC_21_13_7  (
            .in0(N__54869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59207),
            .ce(N__57958),
            .sr(N__57614));
    defparam \pid_side.error_p_reg_esr_11_LC_21_14_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_11_LC_21_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_11_LC_21_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_11_LC_21_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51495),
            .lcout(\pid_side.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59222),
            .ce(N__56607),
            .sr(N__58188));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_21_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_21_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_21_14_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_21_14_7  (
            .in0(N__51468),
            .in1(N__51405),
            .in2(_gnd_net_),
            .in3(N__51273),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_15_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_15_0  (
            .in0(N__54681),
            .in1(N__51843),
            .in2(_gnd_net_),
            .in3(N__55043),
            .lcout(\pid_side.un1_pid_prereg_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_19_LC_21_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_21_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_21_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_19_LC_21_15_1  (
            .in0(N__55044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59239),
            .ce(N__57962),
            .sr(N__57629));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_15_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_15_2  (
            .in0(N__54680),
            .in1(N__51842),
            .in2(_gnd_net_),
            .in3(N__55042),
            .lcout(\pid_side.un1_pid_prereg_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_21_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_21_16_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_21_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_21_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55372),
            .lcout(side_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59255),
            .ce(N__51809),
            .sr(N__57634));
    defparam \pid_side.error_cry_0_c_inv_LC_21_17_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_inv_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_inv_LC_21_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_cry_0_c_inv_LC_21_17_0  (
            .in0(_gnd_net_),
            .in1(N__51756),
            .in2(_gnd_net_),
            .in3(N__51772),
            .lcout(\pid_side.error_axb_0 ),
            .ltout(),
            .carryin(bfn_21_17_0_),
            .carryout(\pid_side.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_21_17_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_21_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_0_c_RNI43F5_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(N__51750),
            .in2(_gnd_net_),
            .in3(N__51717),
            .lcout(\pid_side.error_1 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0 ),
            .carryout(\pid_side.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_21_17_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_21_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_1_c_RNI66G5_LC_21_17_2  (
            .in0(_gnd_net_),
            .in1(N__51714),
            .in2(_gnd_net_),
            .in3(N__51681),
            .lcout(\pid_side.error_2 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1 ),
            .carryout(\pid_side.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_21_17_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_21_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_2_c_RNI89H5_LC_21_17_3  (
            .in0(_gnd_net_),
            .in1(N__51678),
            .in2(_gnd_net_),
            .in3(N__51648),
            .lcout(\pid_side.error_3 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2 ),
            .carryout(\pid_side.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_21_17_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_21_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_c_RNI1SDJ_LC_21_17_4  (
            .in0(_gnd_net_),
            .in1(N__51645),
            .in2(N__51639),
            .in3(N__51603),
            .lcout(\pid_side.error_4 ),
            .ltout(),
            .carryin(\pid_side.error_cry_3 ),
            .carryout(\pid_side.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_21_17_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_21_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIF3ET_LC_21_17_5  (
            .in0(_gnd_net_),
            .in1(N__51600),
            .in2(N__51591),
            .in3(N__51558),
            .lcout(\pid_side.error_5 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0_0 ),
            .carryout(\pid_side.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_21_17_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_21_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_1_0_c_RNII9K11_LC_21_17_6  (
            .in0(_gnd_net_),
            .in1(N__52191),
            .in2(N__52185),
            .in3(N__52149),
            .lcout(\pid_side.error_6 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1_0 ),
            .carryout(\pid_side.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_21_17_7 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_21_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_2_0_c_RNILFQL_LC_21_17_7  (
            .in0(_gnd_net_),
            .in1(N__52146),
            .in2(N__52140),
            .in3(N__52110),
            .lcout(\pid_side.error_7 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2_0 ),
            .carryout(\pid_side.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_21_18_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_21_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIOL0Q_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__52107),
            .in2(N__52101),
            .in3(N__52065),
            .lcout(\pid_side.error_8 ),
            .ltout(),
            .carryin(bfn_21_18_0_),
            .carryout(\pid_side.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_21_18_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_21_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_4_c_RNIC8FJ_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__52062),
            .in2(N__52044),
            .in3(N__52011),
            .lcout(\pid_side.error_9 ),
            .ltout(),
            .carryin(\pid_side.error_cry_4 ),
            .carryout(\pid_side.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_21_18_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_21_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_5_c_RNIM4IS_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__52008),
            .in2(N__51996),
            .in3(N__51954),
            .lcout(\pid_side.error_10 ),
            .ltout(),
            .carryin(\pid_side.error_cry_5 ),
            .carryout(\pid_side.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_21_18_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_21_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_6_c_RNIQBMT_LC_21_18_3  (
            .in0(_gnd_net_),
            .in1(N__51951),
            .in2(_gnd_net_),
            .in3(N__51918),
            .lcout(\pid_side.error_11 ),
            .ltout(),
            .carryin(\pid_side.error_cry_6 ),
            .carryout(\pid_side.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_21_18_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_21_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_7_c_RNIPRDP1_LC_21_18_4  (
            .in0(_gnd_net_),
            .in1(N__51915),
            .in2(N__52506),
            .in3(N__51882),
            .lcout(\pid_side.error_12 ),
            .ltout(),
            .carryin(\pid_side.error_cry_7 ),
            .carryout(\pid_side.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_21_18_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_21_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_8_c_RNIUUKS_LC_21_18_5  (
            .in0(_gnd_net_),
            .in1(N__51879),
            .in2(N__52410),
            .in3(N__51846),
            .lcout(\pid_side.error_13 ),
            .ltout(),
            .carryin(\pid_side.error_cry_8 ),
            .carryout(\pid_side.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_21_18_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_21_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_9_c_RNI13MS_LC_21_18_6  (
            .in0(_gnd_net_),
            .in1(N__53141),
            .in2(N__52779),
            .in3(N__52746),
            .lcout(\pid_side.error_14 ),
            .ltout(),
            .carryin(\pid_side.error_cry_9 ),
            .carryout(\pid_side.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_21_18_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_21_18_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_cry_10_c_RNIBCT11_LC_21_18_7  (
            .in0(N__53142),
            .in1(N__52317),
            .in2(_gnd_net_),
            .in3(N__52743),
            .lcout(\pid_side.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_21_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_21_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_21_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_21_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52713),
            .lcout(drone_H_disp_side_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59294),
            .ce(N__53129),
            .sr(N__57648));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_21_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_21_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_21_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_21_19_1  (
            .in0(N__52586),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59294),
            .ce(N__53129),
            .sr(N__57648));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_21_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_21_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_21_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_21_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52488),
            .lcout(drone_H_disp_side_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59294),
            .ce(N__53129),
            .sr(N__57648));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_21_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_21_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_21_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_21_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52384),
            .lcout(drone_H_disp_side_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59294),
            .ce(N__53129),
            .sr(N__57648));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_21_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_21_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_21_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_21_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52311),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59294),
            .ce(N__53129),
            .sr(N__57648));
    defparam \pid_front.error_d_reg_esr_6_LC_21_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_6_LC_21_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_6_LC_21_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_6_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52230),
            .lcout(\pid_front.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59319),
            .ce(N__58502),
            .sr(N__58181));
    defparam \pid_side.error_d_reg_esr_RNI76TK1_5_LC_22_9_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI76TK1_5_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI76TK1_5_LC_22_9_0 .LUT_INIT=16'b1011111000101000;
    LogicCell40 \pid_side.error_d_reg_esr_RNI76TK1_5_LC_22_9_0  (
            .in0(N__54752),
            .in1(N__53815),
            .in2(N__53795),
            .in3(N__52845),
            .lcout(\pid_side.error_d_reg_esr_RNI76TK1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNILKEQ_5_LC_22_9_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNILKEQ_5_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNILKEQ_5_LC_22_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_esr_RNILKEQ_5_LC_22_9_1  (
            .in0(N__53814),
            .in1(N__53788),
            .in2(_gnd_net_),
            .in3(N__54751),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_40_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI86Q93_5_LC_22_9_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI86Q93_5_LC_22_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI86Q93_5_LC_22_9_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_esr_RNI86Q93_5_LC_22_9_2  (
            .in0(N__52812),
            .in1(N__53601),
            .in2(N__52860),
            .in3(N__52844),
            .lcout(\pid_side.error_d_reg_esr_RNI86Q93Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_22_9_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_22_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_22_9_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_22_9_3  (
            .in0(N__54278),
            .in1(N__52820),
            .in2(_gnd_net_),
            .in3(N__53458),
            .lcout(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_9_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_9_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_9_4  (
            .in0(N__53459),
            .in1(_gnd_net_),
            .in2(N__52824),
            .in3(N__54279),
            .lcout(\pid_side.un1_pid_prereg_17 ),
            .ltout(\pid_side.un1_pid_prereg_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI10TK1_3_LC_22_9_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI10TK1_3_LC_22_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI10TK1_3_LC_22_9_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI10TK1_3_LC_22_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52836),
            .in3(N__53600),
            .lcout(\pid_side.error_p_reg_esr_RNI10TK1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_4_LC_22_9_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_22_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_22_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_4_LC_22_9_6  (
            .in0(N__53460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59168),
            .ce(N__57954),
            .sr(N__57592));
    defparam \pid_side.error_p_reg_esr_RNISPP93_2_LC_22_9_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISPP93_2_LC_22_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISPP93_2_LC_22_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_p_reg_esr_RNISPP93_2_LC_22_9_7  (
            .in0(N__53672),
            .in1(N__53599),
            .in2(N__53628),
            .in3(N__52811),
            .lcout(\pid_side.error_p_reg_esr_RNISPP93Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_5_LC_22_10_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_5_LC_22_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_5_LC_22_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_p_reg_esr_5_LC_22_10_4  (
            .in0(N__52791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59180),
            .ce(N__56592),
            .sr(N__58196));
    defparam \pid_side.error_p_reg_esr_0_LC_22_10_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_0_LC_22_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_0_LC_22_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_0_LC_22_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53031),
            .lcout(\pid_side.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59180),
            .ce(N__56592),
            .sr(N__58196));
    defparam \pid_side.state_RNIK1B71_0_LC_22_11_1 .C_ON=1'b0;
    defparam \pid_side.state_RNIK1B71_0_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIK1B71_0_LC_22_11_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNIK1B71_0_LC_22_11_1  (
            .in0(_gnd_net_),
            .in1(N__53010),
            .in2(_gnd_net_),
            .in3(N__58321),
            .lcout(\pid_side.N_599_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIE47J_9_LC_22_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIE47J_9_LC_22_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIE47J_9_LC_22_11_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \pid_side.error_p_reg_esr_RNIE47J_9_LC_22_11_2  (
            .in0(_gnd_net_),
            .in1(N__54348),
            .in2(_gnd_net_),
            .in3(N__54139),
            .lcout(\pid_side.error_p_reg_esr_RNIE47JZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_15_LC_22_12_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_22_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_22_12_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_15_LC_22_12_3  (
            .in0(_gnd_net_),
            .in1(N__54812),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59208),
            .ce(N__57959),
            .sr(N__57615));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_12_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_12_7 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_12_7  (
            .in0(N__53573),
            .in1(N__54432),
            .in2(_gnd_net_),
            .in3(N__55168),
            .lcout(\pid_side.un1_pid_prereg_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_13_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_22_13_1  (
            .in0(N__54218),
            .in1(N__52904),
            .in2(_gnd_net_),
            .in3(N__54982),
            .lcout(\pid_side.un1_pid_prereg_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_18_LC_22_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_22_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_22_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_18_LC_22_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54984),
            .lcout(\pid_side.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59223),
            .ce(N__57960),
            .sr(N__57622));
    defparam \pid_side.error_d_reg_prev_esr_RNIOHC23_16_LC_22_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOHC23_16_LC_22_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOHC23_16_LC_22_13_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOHC23_16_LC_22_13_4  (
            .in0(N__52938),
            .in1(N__52889),
            .in2(N__54123),
            .in3(N__54094),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOHC23Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_22_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_22_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_22_13_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_22_13_6  (
            .in0(N__54983),
            .in1(_gnd_net_),
            .in2(N__52908),
            .in3(N__54219),
            .lcout(\pid_side.un1_pid_prereg_47 ),
            .ltout(\pid_side.un1_pid_prereg_47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVB6H1_17_LC_22_13_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVB6H1_17_LC_22_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVB6H1_17_LC_22_13_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVB6H1_17_LC_22_13_7  (
            .in0(N__54095),
            .in1(_gnd_net_),
            .in2(N__53556),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIVB6H1Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_10_LC_22_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_22_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_22_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_10_LC_22_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55080),
            .lcout(\pid_side.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59240),
            .ce(N__57963),
            .sr(N__57630));
    defparam \pid_side.error_d_reg_esr_0_LC_22_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_0_LC_22_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_0_LC_22_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_0_LC_22_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53520),
            .lcout(\pid_side.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59256),
            .ce(N__56593),
            .sr(N__58189));
    defparam \pid_side.error_d_reg_esr_4_LC_22_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_4_LC_22_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_4_LC_22_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_4_LC_22_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53472),
            .lcout(\pid_side.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59256),
            .ce(N__56593),
            .sr(N__58189));
    defparam \pid_side.error_d_reg_esr_1_LC_22_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_1_LC_22_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_1_LC_22_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_1_LC_22_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53445),
            .lcout(\pid_side.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59256),
            .ce(N__56593),
            .sr(N__58189));
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_22_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_22_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_22_17_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_4_LC_22_17_6  (
            .in0(_gnd_net_),
            .in1(N__53396),
            .in2(_gnd_net_),
            .in3(N__58322),
            .lcout(xy_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59285),
            .ce(N__55205),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_22_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_22_18_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_22_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_22_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53229),
            .lcout(drone_H_disp_side_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59295),
            .ce(N__53133),
            .sr(N__57649));
    defparam \pid_front.error_d_reg_esr_5_LC_22_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_5_LC_22_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_5_LC_22_23_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_5_LC_22_23_0  (
            .in0(N__53094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59322),
            .ce(N__58495),
            .sr(N__58182));
    defparam \pid_side.error_p_reg_esr_RNI5PH23_1_LC_23_9_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5PH23_1_LC_23_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5PH23_1_LC_23_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5PH23_1_LC_23_9_0  (
            .in0(N__53058),
            .in1(N__53623),
            .in2(N__53673),
            .in3(N__53644),
            .lcout(\pid_side.error_p_reg_esr_RNI5PH23Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_23_9_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_23_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_23_9_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_23_9_1  (
            .in0(N__54240),
            .in1(N__53610),
            .in2(_gnd_net_),
            .in3(N__55133),
            .lcout(\pid_side.un1_pid_prereg_2 ),
            .ltout(\pid_side.un1_pid_prereg_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIRPSK1_2_LC_23_9_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIRPSK1_2_LC_23_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIRPSK1_2_LC_23_9_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIRPSK1_2_LC_23_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53658),
            .in3(N__53624),
            .lcout(\pid_side.error_p_reg_esr_RNIRPSK1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_23_9_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_23_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_23_9_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_23_9_4  (
            .in0(N__54197),
            .in1(N__53582),
            .in2(_gnd_net_),
            .in3(N__54535),
            .lcout(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_23_9_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_23_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_23_9_5 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_2_LC_23_9_5  (
            .in0(N__54536),
            .in1(_gnd_net_),
            .in2(N__53586),
            .in3(N__54198),
            .lcout(\pid_side.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_3_LC_23_9_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_23_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_23_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_3_LC_23_9_6  (
            .in0(N__55134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59181),
            .ce(N__57955),
            .sr(N__57600));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_23_9_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_23_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_23_9_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_23_9_7  (
            .in0(N__54239),
            .in1(N__53609),
            .in2(_gnd_net_),
            .in3(N__55132),
            .lcout(\pid_side.un1_pid_prereg_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_2_LC_23_10_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_23_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_23_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_2_LC_23_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54537),
            .lcout(\pid_side.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59196),
            .ce(N__57957),
            .sr(N__57608));
    defparam \pid_side.error_d_reg_prev_esr_14_LC_23_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_23_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_23_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_14_LC_23_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55170),
            .lcout(\pid_side.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59196),
            .ce(N__57957),
            .sr(N__57608));
    defparam \pid_side.error_p_reg_esr_RNI8U6J_6_LC_23_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI8U6J_6_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI8U6J_6_LC_23_11_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_p_reg_esr_RNI8U6J_6_LC_23_11_2  (
            .in0(_gnd_net_),
            .in1(N__54930),
            .in2(_gnd_net_),
            .in3(N__54912),
            .lcout(),
            .ltout(\pid_side.N_1566_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNIUJLD1_6_LC_23_11_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNIUJLD1_6_LC_23_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNIUJLD1_6_LC_23_11_3 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \pid_side.error_d_reg_esr_RNIUJLD1_6_LC_23_11_3  (
            .in0(N__53819),
            .in1(N__53796),
            .in2(N__53763),
            .in3(N__55014),
            .lcout(\pid_side.error_d_reg_esr_RNIUJLD1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIE47J_0_9_LC_23_11_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIE47J_0_9_LC_23_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIE47J_0_9_LC_23_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIE47J_0_9_LC_23_11_6  (
            .in0(_gnd_net_),
            .in1(N__54347),
            .in2(_gnd_net_),
            .in3(N__54141),
            .lcout(),
            .ltout(\pid_side.N_1578_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNID3MD1_9_LC_23_11_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNID3MD1_9_LC_23_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNID3MD1_9_LC_23_11_7 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \pid_side.error_d_reg_esr_RNID3MD1_9_LC_23_11_7  (
            .in0(N__54057),
            .in1(N__54489),
            .in2(N__53760),
            .in3(N__53691),
            .lcout(\pid_side.error_d_reg_esr_RNID3MD1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI11FQ_9_LC_23_12_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI11FQ_9_LC_23_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI11FQ_9_LC_23_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_esr_RNI11FQ_9_LC_23_12_0  (
            .in0(N__54052),
            .in1(N__54346),
            .in2(_gnd_net_),
            .in3(N__54140),
            .lcout(\pid_side.un1_pid_prereg_80_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_8_LC_23_12_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_23_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_23_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_8_LC_23_12_1  (
            .in0(N__54777),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59224),
            .ce(N__57961),
            .sr(N__57623));
    defparam \pid_side.error_p_reg_esr_RNIC27J_8_LC_23_12_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIC27J_8_LC_23_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIC27J_8_LC_23_12_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIC27J_8_LC_23_12_2  (
            .in0(N__53689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54493),
            .lcout(),
            .ltout(\pid_side.N_1574_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI8ULD1_8_LC_23_12_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI8ULD1_8_LC_23_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI8ULD1_8_LC_23_12_3 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \pid_side.error_d_reg_esr_RNI8ULD1_8_LC_23_12_3  (
            .in0(N__54776),
            .in1(N__54570),
            .in2(N__53730),
            .in3(N__54960),
            .lcout(\pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8 ),
            .ltout(\pid_side.error_d_reg_esr_RNI8ULD1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIL1CR2_8_LC_23_12_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIL1CR2_8_LC_23_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIL1CR2_8_LC_23_12_4 .LUT_INIT=16'b0011001110011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIL1CR2_8_LC_23_12_4  (
            .in0(N__53690),
            .in1(N__53712),
            .in2(N__53706),
            .in3(N__54494),
            .lcout(\pid_side.error_p_reg_esr_RNIL1CR2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNIUTEQ_8_LC_23_12_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNIUTEQ_8_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNIUTEQ_8_LC_23_12_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_d_reg_esr_RNIUTEQ_8_LC_23_12_5  (
            .in0(N__54775),
            .in1(_gnd_net_),
            .in2(N__54495),
            .in3(N__53688),
            .lcout(\pid_side.un1_pid_prereg_70_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_9_LC_23_12_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_23_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_23_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_9_LC_23_12_6  (
            .in0(N__54053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59224),
            .ce(N__57961),
            .sr(N__57623));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_3 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_3  (
            .in0(N__54836),
            .in1(_gnd_net_),
            .in2(N__54081),
            .in3(N__54153),
            .lcout(\pid_side.un1_pid_prereg_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4  (
            .in0(N__54152),
            .in1(N__54077),
            .in2(_gnd_net_),
            .in3(N__54835),
            .lcout(\pid_side.un1_pid_prereg_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_17_LC_23_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54837),
            .lcout(\pid_side.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59257),
            .ce(N__57965),
            .sr(N__57635));
    defparam \pid_side.error_d_reg_esr_9_LC_23_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_9_LC_23_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_9_LC_23_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_9_LC_23_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54069),
            .lcout(\pid_side.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59272),
            .ce(N__56598),
            .sr(N__58190));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_16_0 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_16_0  (
            .in0(N__57980),
            .in1(N__54458),
            .in2(_gnd_net_),
            .in3(N__57997),
            .lcout(\pid_side.un1_pid_prereg_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_23_17_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_23_17_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_23_17_3  (
            .in0(N__54462),
            .in1(N__57981),
            .in2(_gnd_net_),
            .in3(N__58004),
            .lcout(\pid_side.un1_pid_prereg_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_8_LC_23_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_8_LC_23_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_8_LC_23_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_8_LC_23_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53928),
            .lcout(\pid_front.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59327),
            .ce(N__58523),
            .sr(N__58183));
    defparam \pid_front.error_d_reg_esr_12_LC_23_23_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_12_LC_23_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_12_LC_23_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_12_LC_23_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53865),
            .lcout(\pid_front.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59327),
            .ce(N__58523),
            .sr(N__58183));
    defparam \pid_front.error_d_reg_esr_10_LC_23_23_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_10_LC_23_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_10_LC_23_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_10_LC_23_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54327),
            .lcout(\pid_front.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59327),
            .ce(N__58523),
            .sr(N__58183));
    defparam \pid_side.error_p_reg_esr_4_LC_24_9_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_4_LC_24_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_4_LC_24_9_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_p_reg_esr_4_LC_24_9_1  (
            .in0(_gnd_net_),
            .in1(N__54288),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59197),
            .ce(N__56603),
            .sr(N__58204));
    defparam \pid_side.error_p_reg_esr_1_LC_24_9_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_1_LC_24_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_1_LC_24_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_1_LC_24_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54267),
            .lcout(\pid_side.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59197),
            .ce(N__56603),
            .sr(N__58204));
    defparam \pid_side.error_p_reg_esr_3_LC_24_9_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_3_LC_24_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_3_LC_24_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_3_LC_24_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54246),
            .lcout(\pid_side.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59197),
            .ce(N__56603),
            .sr(N__58204));
    defparam \pid_side.error_p_reg_esr_18_LC_24_9_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_18_LC_24_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_18_LC_24_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_18_LC_24_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54231),
            .lcout(\pid_side.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59197),
            .ce(N__56603),
            .sr(N__58204));
    defparam \pid_side.error_p_reg_esr_2_LC_24_9_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_2_LC_24_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_2_LC_24_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_2_LC_24_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54204),
            .lcout(\pid_side.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59197),
            .ce(N__56603),
            .sr(N__58204));
    defparam \pid_side.error_p_reg_esr_16_LC_24_10_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_16_LC_24_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_16_LC_24_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_16_LC_24_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54189),
            .lcout(\pid_side.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59209),
            .ce(N__56608),
            .sr(N__58202));
    defparam \pid_side.error_p_reg_esr_17_LC_24_10_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_17_LC_24_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_17_LC_24_10_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_p_reg_esr_17_LC_24_10_2  (
            .in0(_gnd_net_),
            .in1(N__54162),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59209),
            .ce(N__56608),
            .sr(N__58202));
    defparam \pid_side.error_d_reg_esr_2_LC_24_10_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_2_LC_24_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_2_LC_24_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_2_LC_24_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54549),
            .lcout(\pid_side.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59209),
            .ce(N__56608),
            .sr(N__58202));
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_13_LC_24_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54522),
            .lcout(\pid_side.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59209),
            .ce(N__56608),
            .sr(N__58202));
    defparam \pid_side.error_p_reg_esr_8_LC_24_10_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_8_LC_24_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_8_LC_24_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_8_LC_24_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54501),
            .lcout(\pid_side.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59209),
            .ce(N__56608),
            .sr(N__58202));
    defparam \pid_side.error_p_reg_esr_20_LC_24_10_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_20_LC_24_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_20_LC_24_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_20_LC_24_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54471),
            .lcout(\pid_side.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59209),
            .ce(N__56608),
            .sr(N__58202));
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_14_LC_24_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54441),
            .lcout(\pid_side.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59209),
            .ce(N__56608),
            .sr(N__58202));
    defparam \pid_side.error_p_reg_esr_10_LC_24_11_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_10_LC_24_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_10_LC_24_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_10_LC_24_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54411),
            .lcout(\pid_side.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59225),
            .ce(N__56564),
            .sr(N__58199));
    defparam \pid_side.error_p_reg_esr_15_LC_24_11_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_15_LC_24_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_15_LC_24_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_15_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54384),
            .lcout(\pid_side.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59225),
            .ce(N__56564),
            .sr(N__58199));
    defparam \pid_side.error_p_reg_esr_6_LC_24_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_6_LC_24_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_6_LC_24_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_6_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54360),
            .lcout(\pid_side.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59225),
            .ce(N__56564),
            .sr(N__58199));
    defparam \pid_side.error_p_reg_esr_9_LC_24_11_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_9_LC_24_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_9_LC_24_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_9_LC_24_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54354),
            .lcout(\pid_side.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59225),
            .ce(N__56564),
            .sr(N__58199));
    defparam \pid_side.error_p_reg_esr_7_LC_24_11_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_7_LC_24_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_7_LC_24_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_7_LC_24_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54693),
            .lcout(\pid_side.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59225),
            .ce(N__56564),
            .sr(N__58199));
    defparam \pid_side.error_p_reg_esr_19_LC_24_11_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_19_LC_24_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_19_LC_24_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_19_LC_24_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54687),
            .lcout(\pid_side.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59225),
            .ce(N__56564),
            .sr(N__58199));
    defparam \pid_side.error_p_reg_esr_12_LC_24_11_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_12_LC_24_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_12_LC_24_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_12_LC_24_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54663),
            .lcout(\pid_side.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59225),
            .ce(N__56564),
            .sr(N__58199));
    defparam \pid_side.error_d_reg_prev_esr_7_LC_24_12_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_24_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_24_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_7_LC_24_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56649),
            .lcout(\pid_side.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59241),
            .ce(N__57964),
            .sr(N__57631));
    defparam \pid_side.error_d_reg_esr_RNIRQEQ_7_LC_24_12_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNIRQEQ_7_LC_24_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNIRQEQ_7_LC_24_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_esr_RNIRQEQ_7_LC_24_12_1  (
            .in0(N__56647),
            .in1(N__54567),
            .in2(_gnd_net_),
            .in3(N__54957),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_60_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI1DBR2_6_LC_24_12_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI1DBR2_6_LC_24_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI1DBR2_6_LC_24_12_2 .LUT_INIT=16'b0000111110100101;
    LogicCell40 \pid_side.error_p_reg_esr_RNI1DBR2_6_LC_24_12_2  (
            .in0(N__54910),
            .in1(N__54629),
            .in2(N__54615),
            .in3(N__54928),
            .lcout(\pid_side.error_p_reg_esr_RNI1DBR2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIA07J_7_LC_24_12_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIA07J_7_LC_24_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIA07J_7_LC_24_12_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIA07J_7_LC_24_12_3  (
            .in0(_gnd_net_),
            .in1(N__54568),
            .in2(_gnd_net_),
            .in3(N__54958),
            .lcout(),
            .ltout(\pid_side.N_1570_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_RNI3PLD1_7_LC_24_12_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNI3PLD1_7_LC_24_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNI3PLD1_7_LC_24_12_4 .LUT_INIT=16'b1100111101001101;
    LogicCell40 \pid_side.error_d_reg_esr_RNI3PLD1_7_LC_24_12_4  (
            .in0(N__54911),
            .in1(N__56648),
            .in2(N__54594),
            .in3(N__54929),
            .lcout(\pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7 ),
            .ltout(\pid_side.error_d_reg_esr_RNI3PLD1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIBNBR2_7_LC_24_12_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIBNBR2_7_LC_24_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIBNBR2_7_LC_24_12_5 .LUT_INIT=16'b0110011001010101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIBNBR2_7_LC_24_12_5  (
            .in0(N__54576),
            .in1(N__54569),
            .in2(N__54552),
            .in3(N__54959),
            .lcout(\pid_side.error_p_reg_esr_RNIBNBR2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_6_LC_24_12_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_24_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_24_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_6_LC_24_12_6  (
            .in0(N__55010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59241),
            .ce(N__57964),
            .sr(N__57631));
    defparam \pid_side.error_d_reg_esr_RNIONEQ_6_LC_24_12_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_RNIONEQ_6_LC_24_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_esr_RNIONEQ_6_LC_24_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_esr_RNIONEQ_6_LC_24_12_7  (
            .in0(N__54927),
            .in1(N__54909),
            .in2(_gnd_net_),
            .in3(N__55009),
            .lcout(\pid_side.un1_pid_prereg_50_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_11_LC_24_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_11_LC_24_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_11_LC_24_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_11_LC_24_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54882),
            .lcout(\pid_side.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59258),
            .ce(N__56597),
            .sr(N__58195));
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_17_LC_24_14_0  (
            .in0(N__54846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_15_LC_24_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_15_LC_24_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_15_LC_24_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_15_LC_24_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54822),
            .lcout(\pid_side.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_8_LC_24_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_8_LC_24_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_8_LC_24_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_8_LC_24_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54786),
            .lcout(\pid_side.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_5_LC_24_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_5_LC_24_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_5_LC_24_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_5_LC_24_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54762),
            .lcout(\pid_side.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_12_LC_24_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_12_LC_24_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_12_LC_24_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_12_LC_24_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54720),
            .lcout(\pid_side.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_14_LC_24_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_14_LC_24_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_14_LC_24_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_14_LC_24_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55179),
            .lcout(\pid_side.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_3_LC_24_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_3_LC_24_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_3_LC_24_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_3_LC_24_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55140),
            .lcout(\pid_side.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_13_LC_24_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_13_LC_24_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_13_LC_24_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_13_LC_24_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55116),
            .lcout(\pid_side.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59273),
            .ce(N__56610),
            .sr(N__58194));
    defparam \pid_side.error_d_reg_esr_10_LC_24_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_10_LC_24_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_10_LC_24_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_10_LC_24_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55086),
            .lcout(\pid_side.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59286),
            .ce(N__56599),
            .sr(N__58192));
    defparam \pid_side.error_d_reg_esr_19_LC_24_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_19_LC_24_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_19_LC_24_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_19_LC_24_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55053),
            .lcout(\pid_side.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59286),
            .ce(N__56599),
            .sr(N__58192));
    defparam \pid_side.error_d_reg_esr_20_LC_24_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_20_LC_24_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_20_LC_24_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_20_LC_24_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55029),
            .lcout(\pid_side.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59286),
            .ce(N__56599),
            .sr(N__58192));
    defparam \pid_side.error_d_reg_esr_6_LC_24_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_6_LC_24_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_6_LC_24_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_6_LC_24_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55020),
            .lcout(\pid_side.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59286),
            .ce(N__56599),
            .sr(N__58192));
    defparam \pid_side.error_d_reg_esr_18_LC_24_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_18_LC_24_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_18_LC_24_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_18_LC_24_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54993),
            .lcout(\pid_side.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59286),
            .ce(N__56599),
            .sr(N__58192));
    defparam \pid_side.error_d_reg_esr_7_LC_24_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_7_LC_24_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_7_LC_24_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_7_LC_24_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54966),
            .lcout(\pid_side.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59286),
            .ce(N__56599),
            .sr(N__58192));
    defparam \pid_side.error_d_reg_esr_16_LC_24_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_16_LC_24_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_16_LC_24_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_16_LC_24_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56634),
            .lcout(\pid_side.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59296),
            .ce(N__56609),
            .sr(N__58191));
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_24_17_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_24_17_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_24_17_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_0_LC_24_17_0  (
            .in0(_gnd_net_),
            .in1(N__56508),
            .in2(_gnd_net_),
            .in3(N__58323),
            .lcout(xy_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59304),
            .ce(N__55212),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_24_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_24_17_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_24_17_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_1_LC_24_17_1  (
            .in0(N__58324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56313),
            .lcout(xy_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59304),
            .ce(N__55212),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_24_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_24_17_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_24_17_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_2_LC_24_17_2  (
            .in0(_gnd_net_),
            .in1(N__56140),
            .in2(_gnd_net_),
            .in3(N__58325),
            .lcout(xy_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59304),
            .ce(N__55212),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_24_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_24_17_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_24_17_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_5_LC_24_17_4  (
            .in0(_gnd_net_),
            .in1(N__55931),
            .in2(_gnd_net_),
            .in3(N__58327),
            .lcout(xy_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59304),
            .ce(N__55212),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_24_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_24_17_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_24_17_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_6_LC_24_17_5  (
            .in0(N__58328),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55754),
            .lcout(xy_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59304),
            .ce(N__55212),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_17_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_7_LC_24_17_6  (
            .in0(_gnd_net_),
            .in1(N__55582),
            .in2(_gnd_net_),
            .in3(N__58329),
            .lcout(xy_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59304),
            .ce(N__55212),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_24_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_24_17_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_24_17_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_3_LC_24_17_7  (
            .in0(N__58326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55362),
            .lcout(xy_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59304),
            .ce(N__55212),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_20_LC_24_19_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_24_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_24_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_20_LC_24_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58005),
            .lcout(\pid_side.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59316),
            .ce(N__57966),
            .sr(N__57650));
    defparam \pid_front.error_d_reg_esr_0_LC_24_21_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_0_LC_24_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_0_LC_24_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_0_LC_24_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56949),
            .lcout(\pid_front.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59323),
            .ce(N__58536),
            .sr(N__58187));
    defparam \pid_front.error_d_reg_esr_1_LC_24_22_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_1_LC_24_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_1_LC_24_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_1_LC_24_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56901),
            .lcout(\pid_front.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59328),
            .ce(N__58534),
            .sr(N__58186));
    defparam \pid_front.error_d_reg_esr_13_LC_24_22_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_13_LC_24_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_13_LC_24_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_13_LC_24_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56859),
            .lcout(\pid_front.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59328),
            .ce(N__58534),
            .sr(N__58186));
    defparam \pid_front.error_d_reg_esr_11_LC_24_22_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_11_LC_24_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_11_LC_24_22_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_11_LC_24_22_4  (
            .in0(N__56832),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59328),
            .ce(N__58534),
            .sr(N__58186));
    defparam \pid_front.error_d_reg_esr_9_LC_24_22_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_9_LC_24_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_9_LC_24_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_9_LC_24_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56784),
            .lcout(\pid_front.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59328),
            .ce(N__58534),
            .sr(N__58186));
    defparam \pid_front.error_d_reg_esr_16_LC_24_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_16_LC_24_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_16_LC_24_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_16_LC_24_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56736),
            .lcout(\pid_front.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59332),
            .ce(N__58524),
            .sr(N__58185));
    defparam \pid_front.error_d_reg_esr_17_LC_24_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_17_LC_24_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_17_LC_24_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_17_LC_24_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56682),
            .lcout(\pid_front.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59332),
            .ce(N__58524),
            .sr(N__58185));
    defparam \pid_front.error_d_reg_esr_18_LC_24_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_18_LC_24_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_18_LC_24_23_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_18_LC_24_23_2  (
            .in0(N__59583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59332),
            .ce(N__58524),
            .sr(N__58185));
    defparam \pid_front.error_d_reg_esr_19_LC_24_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_19_LC_24_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_19_LC_24_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_19_LC_24_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59538),
            .lcout(\pid_front.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59332),
            .ce(N__58524),
            .sr(N__58185));
    defparam \pid_front.error_d_reg_esr_20_LC_24_23_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_20_LC_24_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_20_LC_24_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_20_LC_24_23_5  (
            .in0(N__59511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59332),
            .ce(N__58524),
            .sr(N__58185));
    defparam \pid_front.error_d_reg_esr_14_LC_24_23_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_14_LC_24_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_14_LC_24_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_14_LC_24_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59475),
            .lcout(\pid_front.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59332),
            .ce(N__58524),
            .sr(N__58185));
    defparam \pid_front.error_d_reg_esr_4_LC_24_23_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_4_LC_24_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_4_LC_24_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_4_LC_24_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59433),
            .lcout(\pid_front.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59332),
            .ce(N__58524),
            .sr(N__58185));
    defparam \pid_front.error_d_reg_esr_7_LC_24_24_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_7_LC_24_24_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_7_LC_24_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_7_LC_24_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59403),
            .lcout(\pid_front.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59335),
            .ce(N__58535),
            .sr(N__58184));
    defparam \pid_front.error_d_reg_esr_15_LC_24_24_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_15_LC_24_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_15_LC_24_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_15_LC_24_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59367),
            .lcout(\pid_front.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__59335),
            .ce(N__58535),
            .sr(N__58184));
endmodule // Pc2drone
