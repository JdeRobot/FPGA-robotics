-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Apr 6 2019 11:52:24

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2drone
entity Pc2drone is
port (
    uart_input_drone : in std_logic;
    uart_drone_data_rdy_debug : out std_logic;
    uart_commands_input_debug : out std_logic;
    ppm_output : out std_logic;
    uart_input_pc : in std_logic;
    uart_drone_input_debug : out std_logic;
    drone_frame_decoder_data_rdy_debug : out std_logic;
    clk_system : in std_logic);
end Pc2drone;

-- Architecture of Pc2drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2drone is

signal \N__29944\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \pid_alt.O_17\ : std_logic;
signal \pid_alt.O_6\ : std_logic;
signal \pid_alt.O_7\ : std_logic;
signal \pid_alt.O_10\ : std_logic;
signal \pid_alt.O_16\ : std_logic;
signal \pid_alt.O_12\ : std_logic;
signal \pid_alt.O_11\ : std_logic;
signal \pid_alt.O_13\ : std_logic;
signal \pid_alt.O_18\ : std_logic;
signal \pid_alt.O_14\ : std_logic;
signal \pid_alt.O_4\ : std_logic;
signal \pid_alt.O_5\ : std_logic;
signal \pid_alt.O_9\ : std_logic;
signal \pid_alt.O_15\ : std_logic;
signal \pid_alt.O_8\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_0\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_1\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_2\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_3\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_4\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_5\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_7\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_8\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_9\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_10\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_11\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_12\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_14\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pid_alt.error_1\ : std_logic;
signal \pid_alt.error_cry_0\ : std_logic;
signal \pid_alt.error_2\ : std_logic;
signal \pid_alt.error_cry_1\ : std_logic;
signal \pid_alt.error_3\ : std_logic;
signal \pid_alt.error_cry_2\ : std_logic;
signal \pid_alt.error_4\ : std_logic;
signal \pid_alt.error_cry_3\ : std_logic;
signal \pid_alt.error_5\ : std_logic;
signal \pid_alt.error_cry_4\ : std_logic;
signal \pid_alt.error_6\ : std_logic;
signal \pid_alt.error_cry_5\ : std_logic;
signal \pid_alt.error_7\ : std_logic;
signal \pid_alt.error_cry_6\ : std_logic;
signal \pid_alt.error_cry_7\ : std_logic;
signal \pid_alt.error_8\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pid_alt.error_9\ : std_logic;
signal \pid_alt.error_cry_8\ : std_logic;
signal \pid_alt.error_10\ : std_logic;
signal \pid_alt.error_cry_9\ : std_logic;
signal \pid_alt.error_11\ : std_logic;
signal \pid_alt.error_cry_10\ : std_logic;
signal \pid_alt.error_12\ : std_logic;
signal \pid_alt.error_cry_11\ : std_logic;
signal \pid_alt.error_13\ : std_logic;
signal \pid_alt.error_cry_12\ : std_logic;
signal \pid_alt.error_14\ : std_logic;
signal \pid_alt.error_cry_13\ : std_logic;
signal \pid_alt.error_cry_14\ : std_logic;
signal \pid_alt.error_15\ : std_logic;
signal drone_altitude_i_10 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_10\ : std_logic;
signal drone_altitude_i_11 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_11\ : std_logic;
signal \pid_alt.error_axbZ0Z_12\ : std_logic;
signal drone_altitude_12 : std_logic;
signal \pid_alt.error_axbZ0Z_13\ : std_logic;
signal drone_altitude_13 : std_logic;
signal \pid_alt.error_axbZ0Z_14\ : std_logic;
signal drone_altitude_15 : std_logic;
signal drone_altitude_i_7 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_7\ : std_logic;
signal \ppm_encoder_1.N_297_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_13_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_13\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_6\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_6\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\ : std_logic;
signal \bfn_1_28_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_7\ : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_15\ : std_logic;
signal \bfn_1_30_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_17\ : std_logic;
signal alt_kp_0 : std_logic;
signal alt_kp_2 : std_logic;
signal alt_kp_1 : std_logic;
signal \pid_alt.source_p_enZ0\ : std_logic;
signal alt_kp_3 : std_logic;
signal alt_kp_6 : std_logic;
signal \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_8\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_9\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_12\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_10\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_13\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_11\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT10lto13_1\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_15\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_14\ : std_logic;
signal \dron_frame_decoder_1.WDT10_0_i\ : std_logic;
signal drone_altitude_0 : std_logic;
signal \pid_alt.drone_altitude_i_0\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_4\ : std_logic;
signal drone_altitude_i_4 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_5\ : std_logic;
signal drone_altitude_i_5 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_6\ : std_logic;
signal drone_altitude_i_6 : std_logic;
signal drone_altitude_1 : std_logic;
signal \pid_alt.error_axbZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.source_Altitude8lto3Z0Z_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.source_Altitude8lt7_0_cascade_\ : std_logic;
signal drone_altitude_2 : std_logic;
signal \pid_alt.error_axbZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.source_Altitude8lt7_0\ : std_logic;
signal drone_altitude_3 : std_logic;
signal \pid_alt.error_axbZ0Z_3\ : std_logic;
signal alt_command_3 : std_logic;
signal alt_command_1 : std_logic;
signal \Commands_frame_decoder.source_CH1data8lto7Z0Z_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8_cascade_\ : std_logic;
signal alt_command_0 : std_logic;
signal \Commands_frame_decoder.source_CH1data8\ : std_logic;
signal alt_command_2 : std_logic;
signal \Commands_frame_decoder.source_CH1data8lt7_0\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_8\ : std_logic;
signal drone_altitude_i_8 : std_logic;
signal drone_altitude_i_9 : std_logic;
signal drone_altitude_14 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_9\ : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1\ : std_logic;
signal throttle_command_3 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4\ : std_logic;
signal throttle_command_6 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7\ : std_logic;
signal \bfn_2_20_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12\ : std_logic;
signal throttle_command_14 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_13\ : std_logic;
signal throttle_command_1 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\ : std_logic;
signal throttle_command_10 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\ : std_logic;
signal throttle_command_13 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\ : std_logic;
signal throttle_command_4 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\ : std_logic;
signal throttle_command_5 : std_logic;
signal throttle_command_8 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\ : std_logic;
signal throttle_command_7 : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_7\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_7\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_7\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_58_d_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\ : std_logic;
signal throttle_command_2 : std_logic;
signal \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\ : std_logic;
signal throttle_command_0 : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_8\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_9\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_299\ : std_logic;
signal alt_kp_7 : std_logic;
signal alt_kp_5 : std_logic;
signal \dron_frame_decoder_1.state_ns_0_a3_0_0_3_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_a3_0_0_1_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_a3_0_3_1\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_a3_0_3_3\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.N_217_cascade_\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.N_219\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_a2_1_1_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_239\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_0\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_a2_0_2_0\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_243\ : std_logic;
signal alt_command_4 : std_logic;
signal alt_command_5 : std_logic;
signal alt_command_6 : std_logic;
signal alt_command_7 : std_logic;
signal \dron_frame_decoder_1.N_238_0\ : std_logic;
signal \dron_frame_decoder_1.N_237\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.un1_sink_data_valid_5_0_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.un1_sink_data_valid_5_0_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_230_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_6\ : std_logic;
signal uart_drone_data_rdy_debug_c : std_logic;
signal drone_frame_decoder_data_rdy_debug_c : std_logic;
signal \uart_pc.N_152_cascade_\ : std_logic;
signal \uart_pc.CO0_cascade_\ : std_logic;
signal \uart_pc.un1_state_7_0\ : std_logic;
signal throttle_command_9 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\ : std_logic;
signal throttle_command_11 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\ : std_logic;
signal throttle_command_12 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_12\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_303_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_12\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_8\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_9\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_4\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_4\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_5\ : std_logic;
signal \ppm_encoder_1.throttle_RNIN3352Z0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0\ : std_logic;
signal \bfn_3_25_0_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIALN65Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_2\ : std_logic;
signal \ppm_encoder_1.throttle_RNI5V123Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_3\ : std_logic;
signal \ppm_encoder_1.throttle_RNI82223Z0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_2\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_3\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_4\ : std_logic;
signal \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_7\ : std_logic;
signal \ppm_encoder_1.throttle_RNIJII96Z0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_8\ : std_logic;
signal \ppm_encoder_1.throttle_RNIONI96Z0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_8\ : std_logic;
signal \bfn_3_26_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_9\ : std_logic;
signal \ppm_encoder_1.throttle_RNITSI96Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_12\ : std_logic;
signal \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_11\ : std_logic;
signal \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_15\ : std_logic;
signal \bfn_3_27_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_17\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_16\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_9\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_295\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_4\ : std_logic;
signal \reset_module_System.count_1_1_cascade_\ : std_logic;
signal \reset_module_System.reset6_13_cascade_\ : std_logic;
signal \reset_module_System.reset6_3\ : std_logic;
signal \reset_module_System.reset6_17_cascade_\ : std_logic;
signal \reset_module_System.reset6_19_cascade_\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.reset6_11\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_a2_0_3_0\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_0_a4_0_0_2\ : std_logic;
signal uart_drone_data_0 : std_logic;
signal uart_drone_data_1 : std_logic;
signal uart_drone_data_2 : std_logic;
signal uart_drone_data_3 : std_logic;
signal uart_drone_data_4 : std_logic;
signal uart_drone_data_5 : std_logic;
signal uart_drone_data_6 : std_logic;
signal uart_drone_data_7 : std_logic;
signal \uart_drone.state_1_sqmuxa_0\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \bfn_4_19_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\ : std_logic;
signal \Commands_frame_decoder.WDT8lto13_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\ : std_logic;
signal ppm_output_c : std_logic;
signal \ppm_encoder_1.aileronZ0Z_8\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_300_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\ : std_logic;
signal \ppm_encoder_1.N_139_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_14\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_11\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_2_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_11\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_10\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_10\ : std_logic;
signal \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\ : std_logic;
signal \ppm_encoder_1.N_318\ : std_logic;
signal \ppm_encoder_1.N_226\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_10\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_11\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_12\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_18\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\ : std_logic;
signal \bfn_4_29_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_4\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_7\ : std_logic;
signal \bfn_4_30_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \Commands_frame_decoder.state_1_RNIVM1OZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\ : std_logic;
signal alt_kp_4 : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_5\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_i_a2_3_1Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_0_a4_0_3_2\ : std_logic;
signal \Commands_frame_decoder.N_323_cascade_\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_0\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_3\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_4\ : std_logic;
signal \uart_drone.data_AuxZ0Z_5\ : std_logic;
signal \uart_drone.data_AuxZ0Z_6\ : std_logic;
signal \uart_drone.data_AuxZ0Z_7\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_1_cascade_\ : std_logic;
signal \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2\ : std_logic;
signal \uart_drone.state_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.un1_state49_iZ0\ : std_logic;
signal \uart_drone.N_126_li_cascade_\ : std_logic;
signal \uart_drone.N_143_cascade_\ : std_logic;
signal \uart_drone.timer_CountZ1Z_1\ : std_logic;
signal \uart_drone.timer_CountZ0Z_0\ : std_logic;
signal \uart_drone.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_5_19_0_\ : std_logic;
signal \uart_drone.timer_CountZ1Z_2\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_3\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_4\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxa\ : std_logic;
signal \uart_pc.bit_CountZ0Z_2\ : std_logic;
signal \uart_pc.bit_CountZ0Z_1\ : std_logic;
signal \uart_pc.bit_CountZ0Z_0\ : std_logic;
signal \uart_pc.data_Auxce_0_0_0\ : std_logic;
signal \uart_pc.data_AuxZ1Z_0\ : std_logic;
signal \uart_pc.data_Auxce_0_1\ : std_logic;
signal \uart_pc.data_AuxZ1Z_1\ : std_logic;
signal \uart_pc.data_Auxce_0_0_2\ : std_logic;
signal \uart_pc.data_AuxZ1Z_2\ : std_logic;
signal \uart_pc.data_Auxce_0_3\ : std_logic;
signal \uart_pc.data_AuxZ0Z_3\ : std_logic;
signal \uart_pc.data_Auxce_0_0_4\ : std_logic;
signal \uart_pc.data_AuxZ0Z_4\ : std_logic;
signal \uart_pc.data_Auxce_0_5\ : std_logic;
signal \uart_pc.data_AuxZ0Z_5\ : std_logic;
signal \uart_pc.data_AuxZ0Z_7\ : std_logic;
signal \uart_pc.data_Auxce_0_6\ : std_logic;
signal \uart_pc.data_AuxZ0Z_6\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_18\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_1\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_11\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_302_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_5\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_16\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_4\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_4\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_3\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_5\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_5\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.N_296_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_11\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_12\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_\ : std_logic;
signal \ppm_encoder_1.N_237\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.N_237_cascade_\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\ : std_logic;
signal \uart_pc_sync.aux_2__0__0_0\ : std_logic;
signal \uart_pc_sync.aux_3__0__0_0\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa\ : std_logic;
signal \uart_drone.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_1\ : std_logic;
signal \uart_drone.data_Auxce_0_6\ : std_logic;
signal \uart_pc.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_0\ : std_logic;
signal \uart_drone.N_126_li\ : std_logic;
signal \uart_drone.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_0\ : std_logic;
signal \uart_drone.data_Auxce_0_5\ : std_logic;
signal uart_commands_input_debug_c : std_logic;
signal \uart_pc.stateZ0Z_1\ : std_logic;
signal \uart_pc.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_pc.N_152\ : std_logic;
signal \uart_pc.N_144_1\ : std_logic;
signal \uart_pc.N_144_1_cascade_\ : std_logic;
signal \uart_pc.state_1_sqmuxa\ : std_logic;
signal \uart_pc.N_145\ : std_logic;
signal \uart_drone.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_pc.stateZ0Z_2\ : std_logic;
signal \uart_pc.N_143_cascade_\ : std_logic;
signal \uart_pc.state_RNIEAGSZ0Z_4\ : std_logic;
signal \uart_pc.un1_state_4_0\ : std_logic;
signal \uart_pc.N_126_li\ : std_logic;
signal \uart_pc.stateZ0Z_4\ : std_logic;
signal \uart_pc.stateZ0Z_3\ : std_logic;
signal \uart_pc.N_126_li_cascade_\ : std_logic;
signal \uart_pc.un1_state_2_0\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_13\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_10\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_9\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_8\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_14\ : std_logic;
signal \ppm_encoder_1.N_305_cascade_\ : std_logic;
signal \ppm_encoder_1.N_298\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_7\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_13\ : std_logic;
signal \ppm_encoder_1.N_304_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_13\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_12\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux\ : std_logic;
signal \ppm_encoder_1.N_319_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_14\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_6\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_6\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_13\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_13\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_7\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_7\ : std_logic;
signal \ppm_encoder_1.N_590_i\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_0\ : std_logic;
signal \bfn_7_28_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_7\ : std_logic;
signal \bfn_7_29_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_8\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_9\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_15\ : std_logic;
signal \bfn_7_30_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_17\ : std_logic;
signal \ppm_encoder_1.N_168_g\ : std_logic;
signal uart_input_drone_c : std_logic;
signal \uart_drone_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \uart_drone_sync.aux_1__0_Z0Z_0\ : std_logic;
signal \uart_drone_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \uart_drone_sync.aux_3__0_Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\ : std_logic;
signal \frame_decoder_CH2data_7\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \frame_decoder_CH2data_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH2data_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH2data_3\ : std_logic;
signal \frame_decoder_OFF2data_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH2data_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH2data_5\ : std_logic;
signal \frame_decoder_OFF2data_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH2data_6\ : std_logic;
signal \frame_decoder_OFF2data_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7\ : std_logic;
signal \scaler_2.N_521_i_l_ofxZ0\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8\ : std_logic;
signal \uart_drone.data_AuxZ0Z_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_1\ : std_logic;
signal \uart_drone.data_Auxce_0_0_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_2\ : std_logic;
signal \uart_drone.data_Auxce_0_3\ : std_logic;
signal \uart_drone.data_AuxZ0Z_3\ : std_logic;
signal \uart_drone.un1_state_2_0\ : std_logic;
signal uart_drone_input_debug_c : std_logic;
signal \uart_drone.data_AuxZ0Z_4\ : std_logic;
signal \uart_drone.data_Auxce_0_0_4\ : std_logic;
signal \uart_drone.stateZ0Z_2\ : std_logic;
signal \uart_drone.N_145\ : std_logic;
signal \uart_drone.state_RNIOU0NZ0Z_4\ : std_logic;
signal \uart_drone.N_143\ : std_logic;
signal \uart_drone.N_144_1\ : std_logic;
signal \Commands_frame_decoder.state_1_RNO_4Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.WDT8lt14_0\ : std_logic;
signal \uart_pc.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \uart_pc.timer_CountZ1Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_2\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_pc.timer_CountZ0Z_4\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_4\ : std_logic;
signal \uart_pc.timer_CountZ0Z_0\ : std_logic;
signal \uart_pc.timer_CountZ1Z_1\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_1\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_3\ : std_logic;
signal \uart_pc.N_143\ : std_logic;
signal \uart_pc.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_pc.timer_CountZ1Z_3\ : std_logic;
signal \uart_drone.timer_CountZ0Z_4\ : std_logic;
signal \uart_drone.timer_CountZ1Z_3\ : std_logic;
signal \uart_drone.stateZ0Z_4\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_13\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_14\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_12\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_10\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_10\ : std_logic;
signal \ppm_encoder_1.N_301\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_5\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_4\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_8\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_12\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\ : std_logic;
signal \ppm_encoder_1.N_144_17\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\ : std_logic;
signal \ppm_encoder_1.N_144_17_cascade_\ : std_logic;
signal \ppm_encoder_1.N_144\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_13\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_11_mux\ : std_logic;
signal \ppm_encoder_1.N_590_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_14\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_14\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_16\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_16\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_17\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_17\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_15\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_158_d\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_58_d\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_15\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_17\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_16\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_15\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\ : std_logic;
signal uart_input_pc_c : std_logic;
signal \uart_pc_sync.aux_0__0__0_0\ : std_logic;
signal \uart_pc_sync.aux_1__0__0_0\ : std_logic;
signal \frame_decoder_OFF2data_7\ : std_logic;
signal \frame_decoder_OFF2data_1\ : std_logic;
signal \frame_decoder_OFF2data_4\ : std_logic;
signal \frame_decoder_OFF2data_2\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal scaler_2_data_6 : std_logic;
signal \scaler_2.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\ : std_logic;
signal scaler_2_data_7 : std_logic;
signal \scaler_2.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\ : std_logic;
signal scaler_2_data_8 : std_logic;
signal \scaler_2.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\ : std_logic;
signal scaler_2_data_9 : std_logic;
signal \scaler_2.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\ : std_logic;
signal scaler_2_data_10 : std_logic;
signal \scaler_2.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\ : std_logic;
signal scaler_2_data_11 : std_logic;
signal \scaler_2.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\ : std_logic;
signal scaler_2_data_12 : std_logic;
signal \scaler_2.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\ : std_logic;
signal scaler_2_data_13 : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_9\ : std_logic;
signal scaler_2_data_14 : std_logic;
signal scaler_2_data_5 : std_logic;
signal scaler_3_data_5 : std_logic;
signal scaler_4_data_5 : std_logic;
signal \uart_drone.data_Auxce_0_0_0\ : std_logic;
signal scaler_2_data_4 : std_logic;
signal scaler_3_data_4 : std_logic;
signal scaler_4_data_4 : std_logic;
signal \Commands_frame_decoder.N_282_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_0_a4_0_0Z0Z_1\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8lto7Z0Z_1\ : std_logic;
signal \Commands_frame_decoder.N_319_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_318\ : std_logic;
signal \Commands_frame_decoder.N_282_0\ : std_logic;
signal \Commands_frame_decoder.state_1_RNO_1Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_i_0_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.N_323\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_0_a4_0_2_1\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_1\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_13\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pid_altitude_dv_0\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\ : std_logic;
signal pid_altitude_dv : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa\ : std_logic;
signal \frame_decoder_CH4data_7\ : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\ : std_logic;
signal \scaler_2.un2_source_data_0\ : std_logic;
signal \frame_decoder_OFF2data_0\ : std_logic;
signal \frame_decoder_CH2data_0\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\ : std_logic;
signal \frame_decoder_OFF4data_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1_c_RNO_1\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal scaler_4_data_6 : std_logic;
signal \scaler_4.un2_source_data_0_cry_1\ : std_logic;
signal scaler_4_data_7 : std_logic;
signal \scaler_4.un2_source_data_0_cry_2\ : std_logic;
signal scaler_4_data_8 : std_logic;
signal \scaler_4.un2_source_data_0_cry_3\ : std_logic;
signal scaler_4_data_9 : std_logic;
signal \scaler_4.un2_source_data_0_cry_4\ : std_logic;
signal scaler_4_data_10 : std_logic;
signal \scaler_4.un2_source_data_0_cry_5\ : std_logic;
signal scaler_4_data_11 : std_logic;
signal \scaler_4.un2_source_data_0_cry_6\ : std_logic;
signal scaler_4_data_12 : std_logic;
signal \scaler_4.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_8\ : std_logic;
signal scaler_4_data_13 : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_9\ : std_logic;
signal scaler_4_data_14 : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_6\ : std_logic;
signal \uart_drone.stateZ0Z_3\ : std_logic;
signal \uart_drone.N_152\ : std_logic;
signal \uart_drone.un1_state_7_0\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_7\ : std_logic;
signal \frame_decoder_OFF4data_0\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \frame_decoder_OFF4data_1\ : std_logic;
signal \scaler_4.un2_source_data_0\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH4data_2\ : std_logic;
signal \frame_decoder_OFF4data_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH4data_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH4data_4\ : std_logic;
signal \frame_decoder_OFF4data_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH4data_5\ : std_logic;
signal \frame_decoder_OFF4data_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH4data_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7\ : std_logic;
signal \scaler_4.N_545_i_l_ofxZ0\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8_c_RNIS918\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal scaler_3_data_6 : std_logic;
signal \scaler_3.un2_source_data_0_cry_1\ : std_logic;
signal scaler_3_data_7 : std_logic;
signal \scaler_3.un2_source_data_0_cry_2\ : std_logic;
signal scaler_3_data_8 : std_logic;
signal \scaler_3.un2_source_data_0_cry_3\ : std_logic;
signal scaler_3_data_9 : std_logic;
signal \scaler_3.un2_source_data_0_cry_4\ : std_logic;
signal scaler_3_data_10 : std_logic;
signal \scaler_3.un2_source_data_0_cry_5\ : std_logic;
signal scaler_3_data_11 : std_logic;
signal \scaler_3.un2_source_data_0_cry_6\ : std_logic;
signal scaler_3_data_12 : std_logic;
signal \scaler_3.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_8\ : std_logic;
signal scaler_3_data_13 : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_9\ : std_logic;
signal scaler_3_data_14 : std_logic;
signal pc_frame_decoder_dv_0_g : std_logic;
signal \uart_drone.bit_CountZ0Z_2\ : std_logic;
signal \uart_drone.bit_CountZ0Z_1\ : std_logic;
signal \uart_drone.data_Auxce_0_1\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_10\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_i_a4_2_0_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_292\ : std_logic;
signal \uart_drone.un1_state_4_0\ : std_logic;
signal \uart_drone.bit_CountZ0Z_0\ : std_logic;
signal \uart_drone.CO0\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \Commands_frame_decoder.count8_axb_1\ : std_logic;
signal \Commands_frame_decoder.count8_cry_0\ : std_logic;
signal \Commands_frame_decoder.count_i_2\ : std_logic;
signal \Commands_frame_decoder.count8_cry_1\ : std_logic;
signal \Commands_frame_decoder.count8\ : std_logic;
signal \Commands_frame_decoder.count8_THRU_CO\ : std_logic;
signal reset_system : std_logic;
signal \Commands_frame_decoder.count8_THRU_CO_cascade_\ : std_logic;
signal \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0_cascade_\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.CO0\ : std_logic;
signal \Commands_frame_decoder.CO0_cascade_\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_1\ : std_logic;
signal pc_frame_decoder_dv_0 : std_logic;
signal \frame_decoder_CH4data_1\ : std_logic;
signal \frame_decoder_CH4data_0\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH3data_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH3data_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2_c_RNI780L\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH3data_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH3data_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH3data_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\ : std_logic;
signal \scaler_3.N_533_i_l_ofxZ0\ : std_logic;
signal \scaler_3.un2_source_data_0\ : std_logic;
signal \frame_decoder_CH3data_0\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1_c_RNO_0\ : std_logic;
signal \scaler_3.un3_source_data_0_axb_7\ : std_logic;
signal \frame_decoder_CH3data_1\ : std_logic;
signal \frame_decoder_CH3data_7\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\ : std_logic;
signal \Commands_frame_decoder.preinitZ0\ : std_logic;
signal \Commands_frame_decoder.count_1_sqmuxa\ : std_logic;
signal pc_frame_decoder_dv : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Commands_frame_decoder.count8_0_i\ : std_logic;
signal \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0\ : std_logic;
signal \Commands_frame_decoder.state_1_ns_i_a4_2_0_0\ : std_logic;
signal \Commands_frame_decoder.count8_0\ : std_logic;
signal \frame_decoder_OFF4data_3\ : std_logic;
signal \frame_decoder_OFF4data_6\ : std_logic;
signal uart_pc_data_2 : std_logic;
signal \frame_decoder_OFF3data_2\ : std_logic;
signal uart_pc_data_6 : std_logic;
signal \frame_decoder_OFF3data_6\ : std_logic;
signal uart_pc_data_3 : std_logic;
signal \frame_decoder_OFF3data_3\ : std_logic;
signal uart_pc_data_4 : std_logic;
signal \frame_decoder_OFF3data_4\ : std_logic;
signal uart_pc_data_5 : std_logic;
signal \frame_decoder_OFF3data_5\ : std_logic;
signal uart_pc_data_1 : std_logic;
signal \frame_decoder_OFF3data_1\ : std_logic;
signal uart_pc_data_7 : std_logic;
signal \frame_decoder_OFF3data_7\ : std_logic;
signal uart_pc_data_0 : std_logic;
signal \frame_decoder_OFF3data_0\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\ : std_logic;
signal uart_pc_data_rdy : std_logic;
signal \Commands_frame_decoder.source_offset3data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\ : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_8\ : std_logic;
signal \Commands_frame_decoder.N_316\ : std_logic;
signal \Commands_frame_decoder.source_offset3data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.state_1Z0Z_9\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_system_c_g : std_logic;
signal reset_system_g : std_logic;

signal clk_system_wire : std_logic;
signal uart_input_drone_wire : std_logic;
signal uart_input_pc_wire : std_logic;
signal ppm_output_wire : std_logic;
signal uart_drone_data_rdy_debug_wire : std_logic;
signal uart_commands_input_debug_wire : std_logic;
signal drone_frame_decoder_data_rdy_debug_wire : std_logic;
signal uart_drone_input_debug_wire : std_logic;
signal \pid_alt.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    clk_system_wire <= clk_system;
    uart_input_drone_wire <= uart_input_drone;
    uart_input_pc_wire <= uart_input_pc;
    ppm_output <= ppm_output_wire;
    uart_drone_data_rdy_debug <= uart_drone_data_rdy_debug_wire;
    uart_commands_input_debug <= uart_commands_input_debug_wire;
    drone_frame_decoder_data_rdy_debug <= drone_frame_decoder_data_rdy_debug_wire;
    uart_drone_input_debug <= uart_drone_input_debug_wire;
    \pid_alt.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_A_wire\ <= \N__11359\&\N__11377\&\N__11392\&\N__11407\&\N__11422\&\N__11437\&\N__11227\&\N__11242\&\N__11257\&\N__11272\&\N__11284\&\N__11299\&\N__11314\&\N__11329\&\N__11188\&\N__12091\;
    \pid_alt.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__13195\&\N__12018\&\N__13174\&\N__16630\&\N__12037\&\N__11806\&\N__11785\&\N__11824\;
    \pid_alt.O_18\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_17\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_16\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_15\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_14\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_13\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_12\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_11\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_10\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_9\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_8\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_7\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_6\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_5\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_4\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(4);

    \pid_alt.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__27295\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__27264\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_mulonly_0_24_0_O_wire\
        );

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__29942\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29944\,
            DIN => \N__29943\,
            DOUT => \N__29942\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__29944\,
            PADOUT => \N__29943\,
            PADIN => \N__29942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_drone_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29933\,
            DIN => \N__29932\,
            DOUT => \N__29931\,
            PACKAGEPIN => uart_input_drone_wire
        );

    \uart_input_drone_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__29933\,
            PADOUT => \N__29932\,
            PADIN => \N__29931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_drone_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_pc_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29924\,
            DIN => \N__29923\,
            DOUT => \N__29922\,
            PACKAGEPIN => uart_input_pc_wire
        );

    \uart_input_pc_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__29924\,
            PADOUT => \N__29923\,
            PADIN => \N__29922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_pc_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ppm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29915\,
            DIN => \N__29914\,
            DOUT => \N__29913\,
            PACKAGEPIN => ppm_output_wire
        );

    \ppm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__29915\,
            PADOUT => \N__29914\,
            PADIN => \N__29913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15523\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_drone_data_rdy_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29906\,
            DIN => \N__29905\,
            DOUT => \N__29904\,
            PACKAGEPIN => uart_drone_data_rdy_debug_wire
        );

    \uart_drone_data_rdy_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__29906\,
            PADOUT => \N__29905\,
            PADIN => \N__29904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13492\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_commands_input_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29897\,
            DIN => \N__29896\,
            DOUT => \N__29895\,
            PACKAGEPIN => uart_commands_input_debug_wire
        );

    \uart_commands_input_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__29897\,
            PADOUT => \N__29896\,
            PADIN => \N__29895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19151\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \drone_frame_decoder_data_rdy_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29888\,
            DIN => \N__29887\,
            DOUT => \N__29886\,
            PACKAGEPIN => drone_frame_decoder_data_rdy_debug_wire
        );

    \drone_frame_decoder_data_rdy_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__29888\,
            PADOUT => \N__29887\,
            PADIN => \N__29886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13846\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_drone_input_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__29879\,
            DIN => \N__29878\,
            DOUT => \N__29877\,
            PACKAGEPIN => uart_drone_input_debug_wire
        );

    \uart_drone_input_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__29879\,
            PADOUT => \N__29878\,
            PADIN => \N__29877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21749\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__7203\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29857\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__29857\,
            I => \N__29853\
        );

    \I__7201\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29850\
        );

    \I__7200\ : Span4Mux_h
    port map (
            O => \N__29853\,
            I => \N__29840\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__29850\,
            I => \N__29840\
        );

    \I__7198\ : InMux
    port map (
            O => \N__29849\,
            I => \N__29835\
        );

    \I__7197\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29832\
        );

    \I__7196\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29828\
        );

    \I__7195\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29823\
        );

    \I__7194\ : InMux
    port map (
            O => \N__29845\,
            I => \N__29820\
        );

    \I__7193\ : Span4Mux_v
    port map (
            O => \N__29840\,
            I => \N__29817\
        );

    \I__7192\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29814\
        );

    \I__7191\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29811\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__29835\,
            I => \N__29808\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29805\
        );

    \I__7188\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29802\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29799\
        );

    \I__7186\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29796\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__29826\,
            I => \N__29793\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__29823\,
            I => \N__29790\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29787\
        );

    \I__7182\ : Sp12to4
    port map (
            O => \N__29817\,
            I => \N__29782\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__29814\,
            I => \N__29782\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__29811\,
            I => \N__29779\
        );

    \I__7179\ : Span4Mux_v
    port map (
            O => \N__29808\,
            I => \N__29774\
        );

    \I__7178\ : Span4Mux_h
    port map (
            O => \N__29805\,
            I => \N__29774\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__29802\,
            I => \N__29771\
        );

    \I__7176\ : Span4Mux_h
    port map (
            O => \N__29799\,
            I => \N__29766\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__29796\,
            I => \N__29766\
        );

    \I__7174\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29763\
        );

    \I__7173\ : Span4Mux_h
    port map (
            O => \N__29790\,
            I => \N__29760\
        );

    \I__7172\ : Span4Mux_h
    port map (
            O => \N__29787\,
            I => \N__29757\
        );

    \I__7171\ : Span12Mux_h
    port map (
            O => \N__29782\,
            I => \N__29754\
        );

    \I__7170\ : Span4Mux_v
    port map (
            O => \N__29779\,
            I => \N__29745\
        );

    \I__7169\ : Span4Mux_h
    port map (
            O => \N__29774\,
            I => \N__29745\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__29771\,
            I => \N__29745\
        );

    \I__7167\ : Span4Mux_v
    port map (
            O => \N__29766\,
            I => \N__29745\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__29763\,
            I => uart_pc_data_0
        );

    \I__7165\ : Odrv4
    port map (
            O => \N__29760\,
            I => uart_pc_data_0
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__29757\,
            I => uart_pc_data_0
        );

    \I__7163\ : Odrv12
    port map (
            O => \N__29754\,
            I => uart_pc_data_0
        );

    \I__7162\ : Odrv4
    port map (
            O => \N__29745\,
            I => uart_pc_data_0
        );

    \I__7161\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29731\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29726\
        );

    \I__7159\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29723\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__29729\,
            I => \N__29719\
        );

    \I__7157\ : Span4Mux_h
    port map (
            O => \N__29726\,
            I => \N__29716\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29713\
        );

    \I__7155\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29710\
        );

    \I__7154\ : InMux
    port map (
            O => \N__29719\,
            I => \N__29707\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__29716\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__7152\ : Odrv12
    port map (
            O => \N__29713\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__29710\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__29707\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__7149\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29695\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29692\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__29692\,
            I => \N__29689\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__29689\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__7145\ : CascadeMux
    port map (
            O => \N__29686\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_\
        );

    \I__7144\ : CEMux
    port map (
            O => \N__29683\,
            I => \N__29679\
        );

    \I__7143\ : CEMux
    port map (
            O => \N__29682\,
            I => \N__29676\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__29679\,
            I => \N__29673\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__29676\,
            I => \N__29670\
        );

    \I__7140\ : Span4Mux_v
    port map (
            O => \N__29673\,
            I => \N__29667\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__29670\,
            I => \N__29664\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__29667\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__29664\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__7136\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29653\
        );

    \I__7135\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29650\
        );

    \I__7134\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29644\
        );

    \I__7133\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29641\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__29653\,
            I => \N__29637\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__29650\,
            I => \N__29634\
        );

    \I__7130\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29631\
        );

    \I__7129\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29628\
        );

    \I__7128\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29625\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__29644\,
            I => \N__29622\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29619\
        );

    \I__7125\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29615\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__29637\,
            I => \N__29610\
        );

    \I__7123\ : Span4Mux_h
    port map (
            O => \N__29634\,
            I => \N__29601\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__29631\,
            I => \N__29601\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__29628\,
            I => \N__29601\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__29625\,
            I => \N__29601\
        );

    \I__7119\ : Span4Mux_v
    port map (
            O => \N__29622\,
            I => \N__29595\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__29619\,
            I => \N__29595\
        );

    \I__7117\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29592\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__29615\,
            I => \N__29584\
        );

    \I__7115\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29579\
        );

    \I__7114\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29579\
        );

    \I__7113\ : Span4Mux_h
    port map (
            O => \N__29610\,
            I => \N__29574\
        );

    \I__7112\ : Span4Mux_v
    port map (
            O => \N__29601\,
            I => \N__29574\
        );

    \I__7111\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29571\
        );

    \I__7110\ : Span4Mux_h
    port map (
            O => \N__29595\,
            I => \N__29568\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__29592\,
            I => \N__29565\
        );

    \I__7108\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29558\
        );

    \I__7107\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29558\
        );

    \I__7106\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29558\
        );

    \I__7105\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29553\
        );

    \I__7104\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29553\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__29584\,
            I => \N__29548\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29548\
        );

    \I__7101\ : Span4Mux_h
    port map (
            O => \N__29574\,
            I => \N__29545\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__29571\,
            I => uart_pc_data_rdy
        );

    \I__7099\ : Odrv4
    port map (
            O => \N__29568\,
            I => uart_pc_data_rdy
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__29565\,
            I => uart_pc_data_rdy
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__29558\,
            I => uart_pc_data_rdy
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__29553\,
            I => uart_pc_data_rdy
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__29548\,
            I => uart_pc_data_rdy
        );

    \I__7094\ : Odrv4
    port map (
            O => \N__29545\,
            I => uart_pc_data_rdy
        );

    \I__7093\ : CascadeMux
    port map (
            O => \N__29530\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa_cascade_\
        );

    \I__7092\ : CEMux
    port map (
            O => \N__29527\,
            I => \N__29524\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29520\
        );

    \I__7090\ : CEMux
    port map (
            O => \N__29523\,
            I => \N__29517\
        );

    \I__7089\ : Span4Mux_h
    port map (
            O => \N__29520\,
            I => \N__29514\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__29517\,
            I => \N__29511\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__29514\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__7086\ : Odrv12
    port map (
            O => \N__29511\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__7085\ : InMux
    port map (
            O => \N__29506\,
            I => \N__29502\
        );

    \I__7084\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29499\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__29502\,
            I => \N__29496\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__29499\,
            I => \N__29493\
        );

    \I__7081\ : Span4Mux_h
    port map (
            O => \N__29496\,
            I => \N__29490\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__29493\,
            I => \N__29487\
        );

    \I__7079\ : Odrv4
    port map (
            O => \N__29490\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa\
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__29487\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa\
        );

    \I__7077\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29478\
        );

    \I__7076\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29475\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__29478\,
            I => \Commands_frame_decoder.state_1Z0Z_8\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__29475\,
            I => \Commands_frame_decoder.state_1Z0Z_8\
        );

    \I__7073\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29464\
        );

    \I__7072\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29464\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__29464\,
            I => \N__29452\
        );

    \I__7070\ : InMux
    port map (
            O => \N__29463\,
            I => \N__29449\
        );

    \I__7069\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29442\
        );

    \I__7068\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29442\
        );

    \I__7067\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29442\
        );

    \I__7066\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29437\
        );

    \I__7065\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29437\
        );

    \I__7064\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29430\
        );

    \I__7063\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29430\
        );

    \I__7062\ : InMux
    port map (
            O => \N__29455\,
            I => \N__29430\
        );

    \I__7061\ : Span12Mux_h
    port map (
            O => \N__29452\,
            I => \N__29423\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__29449\,
            I => \N__29423\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29423\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29420\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29417\
        );

    \I__7056\ : Odrv12
    port map (
            O => \N__29423\,
            I => \Commands_frame_decoder.N_316\
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__29420\,
            I => \Commands_frame_decoder.N_316\
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__29417\,
            I => \Commands_frame_decoder.N_316\
        );

    \I__7053\ : InMux
    port map (
            O => \N__29410\,
            I => \N__29407\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__29407\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa\
        );

    \I__7051\ : InMux
    port map (
            O => \N__29404\,
            I => \N__29400\
        );

    \I__7050\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29397\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__29400\,
            I => \Commands_frame_decoder.state_1Z0Z_9\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__29397\,
            I => \Commands_frame_decoder.state_1Z0Z_9\
        );

    \I__7047\ : ClkMux
    port map (
            O => \N__29392\,
            I => \N__28987\
        );

    \I__7046\ : ClkMux
    port map (
            O => \N__29391\,
            I => \N__28987\
        );

    \I__7045\ : ClkMux
    port map (
            O => \N__29390\,
            I => \N__28987\
        );

    \I__7044\ : ClkMux
    port map (
            O => \N__29389\,
            I => \N__28987\
        );

    \I__7043\ : ClkMux
    port map (
            O => \N__29388\,
            I => \N__28987\
        );

    \I__7042\ : ClkMux
    port map (
            O => \N__29387\,
            I => \N__28987\
        );

    \I__7041\ : ClkMux
    port map (
            O => \N__29386\,
            I => \N__28987\
        );

    \I__7040\ : ClkMux
    port map (
            O => \N__29385\,
            I => \N__28987\
        );

    \I__7039\ : ClkMux
    port map (
            O => \N__29384\,
            I => \N__28987\
        );

    \I__7038\ : ClkMux
    port map (
            O => \N__29383\,
            I => \N__28987\
        );

    \I__7037\ : ClkMux
    port map (
            O => \N__29382\,
            I => \N__28987\
        );

    \I__7036\ : ClkMux
    port map (
            O => \N__29381\,
            I => \N__28987\
        );

    \I__7035\ : ClkMux
    port map (
            O => \N__29380\,
            I => \N__28987\
        );

    \I__7034\ : ClkMux
    port map (
            O => \N__29379\,
            I => \N__28987\
        );

    \I__7033\ : ClkMux
    port map (
            O => \N__29378\,
            I => \N__28987\
        );

    \I__7032\ : ClkMux
    port map (
            O => \N__29377\,
            I => \N__28987\
        );

    \I__7031\ : ClkMux
    port map (
            O => \N__29376\,
            I => \N__28987\
        );

    \I__7030\ : ClkMux
    port map (
            O => \N__29375\,
            I => \N__28987\
        );

    \I__7029\ : ClkMux
    port map (
            O => \N__29374\,
            I => \N__28987\
        );

    \I__7028\ : ClkMux
    port map (
            O => \N__29373\,
            I => \N__28987\
        );

    \I__7027\ : ClkMux
    port map (
            O => \N__29372\,
            I => \N__28987\
        );

    \I__7026\ : ClkMux
    port map (
            O => \N__29371\,
            I => \N__28987\
        );

    \I__7025\ : ClkMux
    port map (
            O => \N__29370\,
            I => \N__28987\
        );

    \I__7024\ : ClkMux
    port map (
            O => \N__29369\,
            I => \N__28987\
        );

    \I__7023\ : ClkMux
    port map (
            O => \N__29368\,
            I => \N__28987\
        );

    \I__7022\ : ClkMux
    port map (
            O => \N__29367\,
            I => \N__28987\
        );

    \I__7021\ : ClkMux
    port map (
            O => \N__29366\,
            I => \N__28987\
        );

    \I__7020\ : ClkMux
    port map (
            O => \N__29365\,
            I => \N__28987\
        );

    \I__7019\ : ClkMux
    port map (
            O => \N__29364\,
            I => \N__28987\
        );

    \I__7018\ : ClkMux
    port map (
            O => \N__29363\,
            I => \N__28987\
        );

    \I__7017\ : ClkMux
    port map (
            O => \N__29362\,
            I => \N__28987\
        );

    \I__7016\ : ClkMux
    port map (
            O => \N__29361\,
            I => \N__28987\
        );

    \I__7015\ : ClkMux
    port map (
            O => \N__29360\,
            I => \N__28987\
        );

    \I__7014\ : ClkMux
    port map (
            O => \N__29359\,
            I => \N__28987\
        );

    \I__7013\ : ClkMux
    port map (
            O => \N__29358\,
            I => \N__28987\
        );

    \I__7012\ : ClkMux
    port map (
            O => \N__29357\,
            I => \N__28987\
        );

    \I__7011\ : ClkMux
    port map (
            O => \N__29356\,
            I => \N__28987\
        );

    \I__7010\ : ClkMux
    port map (
            O => \N__29355\,
            I => \N__28987\
        );

    \I__7009\ : ClkMux
    port map (
            O => \N__29354\,
            I => \N__28987\
        );

    \I__7008\ : ClkMux
    port map (
            O => \N__29353\,
            I => \N__28987\
        );

    \I__7007\ : ClkMux
    port map (
            O => \N__29352\,
            I => \N__28987\
        );

    \I__7006\ : ClkMux
    port map (
            O => \N__29351\,
            I => \N__28987\
        );

    \I__7005\ : ClkMux
    port map (
            O => \N__29350\,
            I => \N__28987\
        );

    \I__7004\ : ClkMux
    port map (
            O => \N__29349\,
            I => \N__28987\
        );

    \I__7003\ : ClkMux
    port map (
            O => \N__29348\,
            I => \N__28987\
        );

    \I__7002\ : ClkMux
    port map (
            O => \N__29347\,
            I => \N__28987\
        );

    \I__7001\ : ClkMux
    port map (
            O => \N__29346\,
            I => \N__28987\
        );

    \I__7000\ : ClkMux
    port map (
            O => \N__29345\,
            I => \N__28987\
        );

    \I__6999\ : ClkMux
    port map (
            O => \N__29344\,
            I => \N__28987\
        );

    \I__6998\ : ClkMux
    port map (
            O => \N__29343\,
            I => \N__28987\
        );

    \I__6997\ : ClkMux
    port map (
            O => \N__29342\,
            I => \N__28987\
        );

    \I__6996\ : ClkMux
    port map (
            O => \N__29341\,
            I => \N__28987\
        );

    \I__6995\ : ClkMux
    port map (
            O => \N__29340\,
            I => \N__28987\
        );

    \I__6994\ : ClkMux
    port map (
            O => \N__29339\,
            I => \N__28987\
        );

    \I__6993\ : ClkMux
    port map (
            O => \N__29338\,
            I => \N__28987\
        );

    \I__6992\ : ClkMux
    port map (
            O => \N__29337\,
            I => \N__28987\
        );

    \I__6991\ : ClkMux
    port map (
            O => \N__29336\,
            I => \N__28987\
        );

    \I__6990\ : ClkMux
    port map (
            O => \N__29335\,
            I => \N__28987\
        );

    \I__6989\ : ClkMux
    port map (
            O => \N__29334\,
            I => \N__28987\
        );

    \I__6988\ : ClkMux
    port map (
            O => \N__29333\,
            I => \N__28987\
        );

    \I__6987\ : ClkMux
    port map (
            O => \N__29332\,
            I => \N__28987\
        );

    \I__6986\ : ClkMux
    port map (
            O => \N__29331\,
            I => \N__28987\
        );

    \I__6985\ : ClkMux
    port map (
            O => \N__29330\,
            I => \N__28987\
        );

    \I__6984\ : ClkMux
    port map (
            O => \N__29329\,
            I => \N__28987\
        );

    \I__6983\ : ClkMux
    port map (
            O => \N__29328\,
            I => \N__28987\
        );

    \I__6982\ : ClkMux
    port map (
            O => \N__29327\,
            I => \N__28987\
        );

    \I__6981\ : ClkMux
    port map (
            O => \N__29326\,
            I => \N__28987\
        );

    \I__6980\ : ClkMux
    port map (
            O => \N__29325\,
            I => \N__28987\
        );

    \I__6979\ : ClkMux
    port map (
            O => \N__29324\,
            I => \N__28987\
        );

    \I__6978\ : ClkMux
    port map (
            O => \N__29323\,
            I => \N__28987\
        );

    \I__6977\ : ClkMux
    port map (
            O => \N__29322\,
            I => \N__28987\
        );

    \I__6976\ : ClkMux
    port map (
            O => \N__29321\,
            I => \N__28987\
        );

    \I__6975\ : ClkMux
    port map (
            O => \N__29320\,
            I => \N__28987\
        );

    \I__6974\ : ClkMux
    port map (
            O => \N__29319\,
            I => \N__28987\
        );

    \I__6973\ : ClkMux
    port map (
            O => \N__29318\,
            I => \N__28987\
        );

    \I__6972\ : ClkMux
    port map (
            O => \N__29317\,
            I => \N__28987\
        );

    \I__6971\ : ClkMux
    port map (
            O => \N__29316\,
            I => \N__28987\
        );

    \I__6970\ : ClkMux
    port map (
            O => \N__29315\,
            I => \N__28987\
        );

    \I__6969\ : ClkMux
    port map (
            O => \N__29314\,
            I => \N__28987\
        );

    \I__6968\ : ClkMux
    port map (
            O => \N__29313\,
            I => \N__28987\
        );

    \I__6967\ : ClkMux
    port map (
            O => \N__29312\,
            I => \N__28987\
        );

    \I__6966\ : ClkMux
    port map (
            O => \N__29311\,
            I => \N__28987\
        );

    \I__6965\ : ClkMux
    port map (
            O => \N__29310\,
            I => \N__28987\
        );

    \I__6964\ : ClkMux
    port map (
            O => \N__29309\,
            I => \N__28987\
        );

    \I__6963\ : ClkMux
    port map (
            O => \N__29308\,
            I => \N__28987\
        );

    \I__6962\ : ClkMux
    port map (
            O => \N__29307\,
            I => \N__28987\
        );

    \I__6961\ : ClkMux
    port map (
            O => \N__29306\,
            I => \N__28987\
        );

    \I__6960\ : ClkMux
    port map (
            O => \N__29305\,
            I => \N__28987\
        );

    \I__6959\ : ClkMux
    port map (
            O => \N__29304\,
            I => \N__28987\
        );

    \I__6958\ : ClkMux
    port map (
            O => \N__29303\,
            I => \N__28987\
        );

    \I__6957\ : ClkMux
    port map (
            O => \N__29302\,
            I => \N__28987\
        );

    \I__6956\ : ClkMux
    port map (
            O => \N__29301\,
            I => \N__28987\
        );

    \I__6955\ : ClkMux
    port map (
            O => \N__29300\,
            I => \N__28987\
        );

    \I__6954\ : ClkMux
    port map (
            O => \N__29299\,
            I => \N__28987\
        );

    \I__6953\ : ClkMux
    port map (
            O => \N__29298\,
            I => \N__28987\
        );

    \I__6952\ : ClkMux
    port map (
            O => \N__29297\,
            I => \N__28987\
        );

    \I__6951\ : ClkMux
    port map (
            O => \N__29296\,
            I => \N__28987\
        );

    \I__6950\ : ClkMux
    port map (
            O => \N__29295\,
            I => \N__28987\
        );

    \I__6949\ : ClkMux
    port map (
            O => \N__29294\,
            I => \N__28987\
        );

    \I__6948\ : ClkMux
    port map (
            O => \N__29293\,
            I => \N__28987\
        );

    \I__6947\ : ClkMux
    port map (
            O => \N__29292\,
            I => \N__28987\
        );

    \I__6946\ : ClkMux
    port map (
            O => \N__29291\,
            I => \N__28987\
        );

    \I__6945\ : ClkMux
    port map (
            O => \N__29290\,
            I => \N__28987\
        );

    \I__6944\ : ClkMux
    port map (
            O => \N__29289\,
            I => \N__28987\
        );

    \I__6943\ : ClkMux
    port map (
            O => \N__29288\,
            I => \N__28987\
        );

    \I__6942\ : ClkMux
    port map (
            O => \N__29287\,
            I => \N__28987\
        );

    \I__6941\ : ClkMux
    port map (
            O => \N__29286\,
            I => \N__28987\
        );

    \I__6940\ : ClkMux
    port map (
            O => \N__29285\,
            I => \N__28987\
        );

    \I__6939\ : ClkMux
    port map (
            O => \N__29284\,
            I => \N__28987\
        );

    \I__6938\ : ClkMux
    port map (
            O => \N__29283\,
            I => \N__28987\
        );

    \I__6937\ : ClkMux
    port map (
            O => \N__29282\,
            I => \N__28987\
        );

    \I__6936\ : ClkMux
    port map (
            O => \N__29281\,
            I => \N__28987\
        );

    \I__6935\ : ClkMux
    port map (
            O => \N__29280\,
            I => \N__28987\
        );

    \I__6934\ : ClkMux
    port map (
            O => \N__29279\,
            I => \N__28987\
        );

    \I__6933\ : ClkMux
    port map (
            O => \N__29278\,
            I => \N__28987\
        );

    \I__6932\ : ClkMux
    port map (
            O => \N__29277\,
            I => \N__28987\
        );

    \I__6931\ : ClkMux
    port map (
            O => \N__29276\,
            I => \N__28987\
        );

    \I__6930\ : ClkMux
    port map (
            O => \N__29275\,
            I => \N__28987\
        );

    \I__6929\ : ClkMux
    port map (
            O => \N__29274\,
            I => \N__28987\
        );

    \I__6928\ : ClkMux
    port map (
            O => \N__29273\,
            I => \N__28987\
        );

    \I__6927\ : ClkMux
    port map (
            O => \N__29272\,
            I => \N__28987\
        );

    \I__6926\ : ClkMux
    port map (
            O => \N__29271\,
            I => \N__28987\
        );

    \I__6925\ : ClkMux
    port map (
            O => \N__29270\,
            I => \N__28987\
        );

    \I__6924\ : ClkMux
    port map (
            O => \N__29269\,
            I => \N__28987\
        );

    \I__6923\ : ClkMux
    port map (
            O => \N__29268\,
            I => \N__28987\
        );

    \I__6922\ : ClkMux
    port map (
            O => \N__29267\,
            I => \N__28987\
        );

    \I__6921\ : ClkMux
    port map (
            O => \N__29266\,
            I => \N__28987\
        );

    \I__6920\ : ClkMux
    port map (
            O => \N__29265\,
            I => \N__28987\
        );

    \I__6919\ : ClkMux
    port map (
            O => \N__29264\,
            I => \N__28987\
        );

    \I__6918\ : ClkMux
    port map (
            O => \N__29263\,
            I => \N__28987\
        );

    \I__6917\ : ClkMux
    port map (
            O => \N__29262\,
            I => \N__28987\
        );

    \I__6916\ : ClkMux
    port map (
            O => \N__29261\,
            I => \N__28987\
        );

    \I__6915\ : ClkMux
    port map (
            O => \N__29260\,
            I => \N__28987\
        );

    \I__6914\ : ClkMux
    port map (
            O => \N__29259\,
            I => \N__28987\
        );

    \I__6913\ : ClkMux
    port map (
            O => \N__29258\,
            I => \N__28987\
        );

    \I__6912\ : GlobalMux
    port map (
            O => \N__28987\,
            I => \N__28984\
        );

    \I__6911\ : gio2CtrlBuf
    port map (
            O => \N__28984\,
            I => clk_system_c_g
        );

    \I__6910\ : CascadeMux
    port map (
            O => \N__28981\,
            I => \N__28973\
        );

    \I__6909\ : CascadeMux
    port map (
            O => \N__28980\,
            I => \N__28969\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__28979\,
            I => \N__28965\
        );

    \I__6907\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28921\
        );

    \I__6906\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28916\
        );

    \I__6905\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28916\
        );

    \I__6904\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28913\
        );

    \I__6903\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28908\
        );

    \I__6902\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28908\
        );

    \I__6901\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28905\
        );

    \I__6900\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28900\
        );

    \I__6899\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28900\
        );

    \I__6898\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28897\
        );

    \I__6897\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28892\
        );

    \I__6896\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28892\
        );

    \I__6895\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28889\
        );

    \I__6894\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28878\
        );

    \I__6893\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28878\
        );

    \I__6892\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28878\
        );

    \I__6891\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28878\
        );

    \I__6890\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28878\
        );

    \I__6889\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28867\
        );

    \I__6888\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28867\
        );

    \I__6887\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28867\
        );

    \I__6886\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28867\
        );

    \I__6885\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28867\
        );

    \I__6884\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28862\
        );

    \I__6883\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28862\
        );

    \I__6882\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28855\
        );

    \I__6881\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28855\
        );

    \I__6880\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28855\
        );

    \I__6879\ : InMux
    port map (
            O => \N__28944\,
            I => \N__28844\
        );

    \I__6878\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28844\
        );

    \I__6877\ : InMux
    port map (
            O => \N__28942\,
            I => \N__28844\
        );

    \I__6876\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28844\
        );

    \I__6875\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28844\
        );

    \I__6874\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28841\
        );

    \I__6873\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28838\
        );

    \I__6872\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28835\
        );

    \I__6871\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28830\
        );

    \I__6870\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28830\
        );

    \I__6869\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28827\
        );

    \I__6868\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28824\
        );

    \I__6867\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28821\
        );

    \I__6866\ : InMux
    port map (
            O => \N__28931\,
            I => \N__28818\
        );

    \I__6865\ : InMux
    port map (
            O => \N__28930\,
            I => \N__28815\
        );

    \I__6864\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28812\
        );

    \I__6863\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28809\
        );

    \I__6862\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28806\
        );

    \I__6861\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28803\
        );

    \I__6860\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28800\
        );

    \I__6859\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28797\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__28921\,
            I => \N__28708\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__28916\,
            I => \N__28705\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28702\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__28908\,
            I => \N__28699\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28696\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__28900\,
            I => \N__28693\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__28897\,
            I => \N__28690\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__28892\,
            I => \N__28687\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__28889\,
            I => \N__28684\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__28878\,
            I => \N__28681\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28678\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__28862\,
            I => \N__28675\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__28855\,
            I => \N__28672\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28669\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28666\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__28838\,
            I => \N__28663\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28660\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__28830\,
            I => \N__28657\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__28827\,
            I => \N__28654\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28651\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__28821\,
            I => \N__28648\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28645\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__28815\,
            I => \N__28642\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__28812\,
            I => \N__28639\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28636\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__28806\,
            I => \N__28633\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28630\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__28800\,
            I => \N__28627\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28624\
        );

    \I__6829\ : SRMux
    port map (
            O => \N__28796\,
            I => \N__28393\
        );

    \I__6828\ : SRMux
    port map (
            O => \N__28795\,
            I => \N__28393\
        );

    \I__6827\ : SRMux
    port map (
            O => \N__28794\,
            I => \N__28393\
        );

    \I__6826\ : SRMux
    port map (
            O => \N__28793\,
            I => \N__28393\
        );

    \I__6825\ : SRMux
    port map (
            O => \N__28792\,
            I => \N__28393\
        );

    \I__6824\ : SRMux
    port map (
            O => \N__28791\,
            I => \N__28393\
        );

    \I__6823\ : SRMux
    port map (
            O => \N__28790\,
            I => \N__28393\
        );

    \I__6822\ : SRMux
    port map (
            O => \N__28789\,
            I => \N__28393\
        );

    \I__6821\ : SRMux
    port map (
            O => \N__28788\,
            I => \N__28393\
        );

    \I__6820\ : SRMux
    port map (
            O => \N__28787\,
            I => \N__28393\
        );

    \I__6819\ : SRMux
    port map (
            O => \N__28786\,
            I => \N__28393\
        );

    \I__6818\ : SRMux
    port map (
            O => \N__28785\,
            I => \N__28393\
        );

    \I__6817\ : SRMux
    port map (
            O => \N__28784\,
            I => \N__28393\
        );

    \I__6816\ : SRMux
    port map (
            O => \N__28783\,
            I => \N__28393\
        );

    \I__6815\ : SRMux
    port map (
            O => \N__28782\,
            I => \N__28393\
        );

    \I__6814\ : SRMux
    port map (
            O => \N__28781\,
            I => \N__28393\
        );

    \I__6813\ : SRMux
    port map (
            O => \N__28780\,
            I => \N__28393\
        );

    \I__6812\ : SRMux
    port map (
            O => \N__28779\,
            I => \N__28393\
        );

    \I__6811\ : SRMux
    port map (
            O => \N__28778\,
            I => \N__28393\
        );

    \I__6810\ : SRMux
    port map (
            O => \N__28777\,
            I => \N__28393\
        );

    \I__6809\ : SRMux
    port map (
            O => \N__28776\,
            I => \N__28393\
        );

    \I__6808\ : SRMux
    port map (
            O => \N__28775\,
            I => \N__28393\
        );

    \I__6807\ : SRMux
    port map (
            O => \N__28774\,
            I => \N__28393\
        );

    \I__6806\ : SRMux
    port map (
            O => \N__28773\,
            I => \N__28393\
        );

    \I__6805\ : SRMux
    port map (
            O => \N__28772\,
            I => \N__28393\
        );

    \I__6804\ : SRMux
    port map (
            O => \N__28771\,
            I => \N__28393\
        );

    \I__6803\ : SRMux
    port map (
            O => \N__28770\,
            I => \N__28393\
        );

    \I__6802\ : SRMux
    port map (
            O => \N__28769\,
            I => \N__28393\
        );

    \I__6801\ : SRMux
    port map (
            O => \N__28768\,
            I => \N__28393\
        );

    \I__6800\ : SRMux
    port map (
            O => \N__28767\,
            I => \N__28393\
        );

    \I__6799\ : SRMux
    port map (
            O => \N__28766\,
            I => \N__28393\
        );

    \I__6798\ : SRMux
    port map (
            O => \N__28765\,
            I => \N__28393\
        );

    \I__6797\ : SRMux
    port map (
            O => \N__28764\,
            I => \N__28393\
        );

    \I__6796\ : SRMux
    port map (
            O => \N__28763\,
            I => \N__28393\
        );

    \I__6795\ : SRMux
    port map (
            O => \N__28762\,
            I => \N__28393\
        );

    \I__6794\ : SRMux
    port map (
            O => \N__28761\,
            I => \N__28393\
        );

    \I__6793\ : SRMux
    port map (
            O => \N__28760\,
            I => \N__28393\
        );

    \I__6792\ : SRMux
    port map (
            O => \N__28759\,
            I => \N__28393\
        );

    \I__6791\ : SRMux
    port map (
            O => \N__28758\,
            I => \N__28393\
        );

    \I__6790\ : SRMux
    port map (
            O => \N__28757\,
            I => \N__28393\
        );

    \I__6789\ : SRMux
    port map (
            O => \N__28756\,
            I => \N__28393\
        );

    \I__6788\ : SRMux
    port map (
            O => \N__28755\,
            I => \N__28393\
        );

    \I__6787\ : SRMux
    port map (
            O => \N__28754\,
            I => \N__28393\
        );

    \I__6786\ : SRMux
    port map (
            O => \N__28753\,
            I => \N__28393\
        );

    \I__6785\ : SRMux
    port map (
            O => \N__28752\,
            I => \N__28393\
        );

    \I__6784\ : SRMux
    port map (
            O => \N__28751\,
            I => \N__28393\
        );

    \I__6783\ : SRMux
    port map (
            O => \N__28750\,
            I => \N__28393\
        );

    \I__6782\ : SRMux
    port map (
            O => \N__28749\,
            I => \N__28393\
        );

    \I__6781\ : SRMux
    port map (
            O => \N__28748\,
            I => \N__28393\
        );

    \I__6780\ : SRMux
    port map (
            O => \N__28747\,
            I => \N__28393\
        );

    \I__6779\ : SRMux
    port map (
            O => \N__28746\,
            I => \N__28393\
        );

    \I__6778\ : SRMux
    port map (
            O => \N__28745\,
            I => \N__28393\
        );

    \I__6777\ : SRMux
    port map (
            O => \N__28744\,
            I => \N__28393\
        );

    \I__6776\ : SRMux
    port map (
            O => \N__28743\,
            I => \N__28393\
        );

    \I__6775\ : SRMux
    port map (
            O => \N__28742\,
            I => \N__28393\
        );

    \I__6774\ : SRMux
    port map (
            O => \N__28741\,
            I => \N__28393\
        );

    \I__6773\ : SRMux
    port map (
            O => \N__28740\,
            I => \N__28393\
        );

    \I__6772\ : SRMux
    port map (
            O => \N__28739\,
            I => \N__28393\
        );

    \I__6771\ : SRMux
    port map (
            O => \N__28738\,
            I => \N__28393\
        );

    \I__6770\ : SRMux
    port map (
            O => \N__28737\,
            I => \N__28393\
        );

    \I__6769\ : SRMux
    port map (
            O => \N__28736\,
            I => \N__28393\
        );

    \I__6768\ : SRMux
    port map (
            O => \N__28735\,
            I => \N__28393\
        );

    \I__6767\ : SRMux
    port map (
            O => \N__28734\,
            I => \N__28393\
        );

    \I__6766\ : SRMux
    port map (
            O => \N__28733\,
            I => \N__28393\
        );

    \I__6765\ : SRMux
    port map (
            O => \N__28732\,
            I => \N__28393\
        );

    \I__6764\ : SRMux
    port map (
            O => \N__28731\,
            I => \N__28393\
        );

    \I__6763\ : SRMux
    port map (
            O => \N__28730\,
            I => \N__28393\
        );

    \I__6762\ : SRMux
    port map (
            O => \N__28729\,
            I => \N__28393\
        );

    \I__6761\ : SRMux
    port map (
            O => \N__28728\,
            I => \N__28393\
        );

    \I__6760\ : SRMux
    port map (
            O => \N__28727\,
            I => \N__28393\
        );

    \I__6759\ : SRMux
    port map (
            O => \N__28726\,
            I => \N__28393\
        );

    \I__6758\ : SRMux
    port map (
            O => \N__28725\,
            I => \N__28393\
        );

    \I__6757\ : SRMux
    port map (
            O => \N__28724\,
            I => \N__28393\
        );

    \I__6756\ : SRMux
    port map (
            O => \N__28723\,
            I => \N__28393\
        );

    \I__6755\ : SRMux
    port map (
            O => \N__28722\,
            I => \N__28393\
        );

    \I__6754\ : SRMux
    port map (
            O => \N__28721\,
            I => \N__28393\
        );

    \I__6753\ : SRMux
    port map (
            O => \N__28720\,
            I => \N__28393\
        );

    \I__6752\ : SRMux
    port map (
            O => \N__28719\,
            I => \N__28393\
        );

    \I__6751\ : SRMux
    port map (
            O => \N__28718\,
            I => \N__28393\
        );

    \I__6750\ : SRMux
    port map (
            O => \N__28717\,
            I => \N__28393\
        );

    \I__6749\ : SRMux
    port map (
            O => \N__28716\,
            I => \N__28393\
        );

    \I__6748\ : SRMux
    port map (
            O => \N__28715\,
            I => \N__28393\
        );

    \I__6747\ : SRMux
    port map (
            O => \N__28714\,
            I => \N__28393\
        );

    \I__6746\ : SRMux
    port map (
            O => \N__28713\,
            I => \N__28393\
        );

    \I__6745\ : SRMux
    port map (
            O => \N__28712\,
            I => \N__28393\
        );

    \I__6744\ : SRMux
    port map (
            O => \N__28711\,
            I => \N__28393\
        );

    \I__6743\ : Glb2LocalMux
    port map (
            O => \N__28708\,
            I => \N__28393\
        );

    \I__6742\ : Glb2LocalMux
    port map (
            O => \N__28705\,
            I => \N__28393\
        );

    \I__6741\ : Glb2LocalMux
    port map (
            O => \N__28702\,
            I => \N__28393\
        );

    \I__6740\ : Glb2LocalMux
    port map (
            O => \N__28699\,
            I => \N__28393\
        );

    \I__6739\ : Glb2LocalMux
    port map (
            O => \N__28696\,
            I => \N__28393\
        );

    \I__6738\ : Glb2LocalMux
    port map (
            O => \N__28693\,
            I => \N__28393\
        );

    \I__6737\ : Glb2LocalMux
    port map (
            O => \N__28690\,
            I => \N__28393\
        );

    \I__6736\ : Glb2LocalMux
    port map (
            O => \N__28687\,
            I => \N__28393\
        );

    \I__6735\ : Glb2LocalMux
    port map (
            O => \N__28684\,
            I => \N__28393\
        );

    \I__6734\ : Glb2LocalMux
    port map (
            O => \N__28681\,
            I => \N__28393\
        );

    \I__6733\ : Glb2LocalMux
    port map (
            O => \N__28678\,
            I => \N__28393\
        );

    \I__6732\ : Glb2LocalMux
    port map (
            O => \N__28675\,
            I => \N__28393\
        );

    \I__6731\ : Glb2LocalMux
    port map (
            O => \N__28672\,
            I => \N__28393\
        );

    \I__6730\ : Glb2LocalMux
    port map (
            O => \N__28669\,
            I => \N__28393\
        );

    \I__6729\ : Glb2LocalMux
    port map (
            O => \N__28666\,
            I => \N__28393\
        );

    \I__6728\ : Glb2LocalMux
    port map (
            O => \N__28663\,
            I => \N__28393\
        );

    \I__6727\ : Glb2LocalMux
    port map (
            O => \N__28660\,
            I => \N__28393\
        );

    \I__6726\ : Glb2LocalMux
    port map (
            O => \N__28657\,
            I => \N__28393\
        );

    \I__6725\ : Glb2LocalMux
    port map (
            O => \N__28654\,
            I => \N__28393\
        );

    \I__6724\ : Glb2LocalMux
    port map (
            O => \N__28651\,
            I => \N__28393\
        );

    \I__6723\ : Glb2LocalMux
    port map (
            O => \N__28648\,
            I => \N__28393\
        );

    \I__6722\ : Glb2LocalMux
    port map (
            O => \N__28645\,
            I => \N__28393\
        );

    \I__6721\ : Glb2LocalMux
    port map (
            O => \N__28642\,
            I => \N__28393\
        );

    \I__6720\ : Glb2LocalMux
    port map (
            O => \N__28639\,
            I => \N__28393\
        );

    \I__6719\ : Glb2LocalMux
    port map (
            O => \N__28636\,
            I => \N__28393\
        );

    \I__6718\ : Glb2LocalMux
    port map (
            O => \N__28633\,
            I => \N__28393\
        );

    \I__6717\ : Glb2LocalMux
    port map (
            O => \N__28630\,
            I => \N__28393\
        );

    \I__6716\ : Glb2LocalMux
    port map (
            O => \N__28627\,
            I => \N__28393\
        );

    \I__6715\ : Glb2LocalMux
    port map (
            O => \N__28624\,
            I => \N__28393\
        );

    \I__6714\ : GlobalMux
    port map (
            O => \N__28393\,
            I => \N__28390\
        );

    \I__6713\ : gio2CtrlBuf
    port map (
            O => \N__28390\,
            I => reset_system_g
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__28387\,
            I => \N__28384\
        );

    \I__6711\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28381\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__28381\,
            I => \N__28378\
        );

    \I__6709\ : Odrv12
    port map (
            O => \N__28378\,
            I => \frame_decoder_OFF4data_3\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__28375\,
            I => \N__28372\
        );

    \I__6707\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28369\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__28369\,
            I => \N__28366\
        );

    \I__6705\ : Odrv4
    port map (
            O => \N__28366\,
            I => \frame_decoder_OFF4data_6\
        );

    \I__6704\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28357\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__28362\,
            I => \N__28350\
        );

    \I__6702\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28347\
        );

    \I__6701\ : InMux
    port map (
            O => \N__28360\,
            I => \N__28344\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__28357\,
            I => \N__28341\
        );

    \I__6699\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28338\
        );

    \I__6698\ : InMux
    port map (
            O => \N__28355\,
            I => \N__28335\
        );

    \I__6697\ : InMux
    port map (
            O => \N__28354\,
            I => \N__28332\
        );

    \I__6696\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28329\
        );

    \I__6695\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28326\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__28347\,
            I => \N__28323\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__28344\,
            I => \N__28316\
        );

    \I__6692\ : Span4Mux_v
    port map (
            O => \N__28341\,
            I => \N__28316\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__28338\,
            I => \N__28316\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__28335\,
            I => \N__28313\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__28332\,
            I => \N__28302\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__28329\,
            I => \N__28302\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__28326\,
            I => \N__28299\
        );

    \I__6686\ : Span4Mux_v
    port map (
            O => \N__28323\,
            I => \N__28294\
        );

    \I__6685\ : Span4Mux_h
    port map (
            O => \N__28316\,
            I => \N__28294\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__28313\,
            I => \N__28291\
        );

    \I__6683\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28288\
        );

    \I__6682\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28285\
        );

    \I__6681\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28282\
        );

    \I__6680\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28279\
        );

    \I__6679\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28276\
        );

    \I__6678\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28273\
        );

    \I__6677\ : Span12Mux_h
    port map (
            O => \N__28302\,
            I => \N__28270\
        );

    \I__6676\ : Span4Mux_v
    port map (
            O => \N__28299\,
            I => \N__28267\
        );

    \I__6675\ : Span4Mux_h
    port map (
            O => \N__28294\,
            I => \N__28260\
        );

    \I__6674\ : Span4Mux_v
    port map (
            O => \N__28291\,
            I => \N__28260\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__28288\,
            I => \N__28260\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__28285\,
            I => \N__28251\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__28282\,
            I => \N__28251\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__28279\,
            I => \N__28251\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__28276\,
            I => \N__28251\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__28273\,
            I => uart_pc_data_2
        );

    \I__6667\ : Odrv12
    port map (
            O => \N__28270\,
            I => uart_pc_data_2
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__28267\,
            I => uart_pc_data_2
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__28260\,
            I => uart_pc_data_2
        );

    \I__6664\ : Odrv12
    port map (
            O => \N__28251\,
            I => uart_pc_data_2
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__28240\,
            I => \N__28237\
        );

    \I__6662\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__28234\,
            I => \frame_decoder_OFF3data_2\
        );

    \I__6660\ : InMux
    port map (
            O => \N__28231\,
            I => \N__28225\
        );

    \I__6659\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28222\
        );

    \I__6658\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28217\
        );

    \I__6657\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28214\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__28225\,
            I => \N__28210\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__28222\,
            I => \N__28207\
        );

    \I__6654\ : InMux
    port map (
            O => \N__28221\,
            I => \N__28204\
        );

    \I__6653\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28200\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__28217\,
            I => \N__28195\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__28214\,
            I => \N__28195\
        );

    \I__6650\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28191\
        );

    \I__6649\ : Span4Mux_v
    port map (
            O => \N__28210\,
            I => \N__28188\
        );

    \I__6648\ : Span4Mux_s3_h
    port map (
            O => \N__28207\,
            I => \N__28185\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28182\
        );

    \I__6646\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28179\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__28200\,
            I => \N__28176\
        );

    \I__6644\ : Span4Mux_v
    port map (
            O => \N__28195\,
            I => \N__28172\
        );

    \I__6643\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28169\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__28191\,
            I => \N__28165\
        );

    \I__6641\ : Span4Mux_h
    port map (
            O => \N__28188\,
            I => \N__28154\
        );

    \I__6640\ : Span4Mux_v
    port map (
            O => \N__28185\,
            I => \N__28154\
        );

    \I__6639\ : Span4Mux_v
    port map (
            O => \N__28182\,
            I => \N__28154\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__28179\,
            I => \N__28154\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__28176\,
            I => \N__28154\
        );

    \I__6636\ : CascadeMux
    port map (
            O => \N__28175\,
            I => \N__28151\
        );

    \I__6635\ : Sp12to4
    port map (
            O => \N__28172\,
            I => \N__28146\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__28169\,
            I => \N__28146\
        );

    \I__6633\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28143\
        );

    \I__6632\ : Span12Mux_v
    port map (
            O => \N__28165\,
            I => \N__28138\
        );

    \I__6631\ : Sp12to4
    port map (
            O => \N__28154\,
            I => \N__28138\
        );

    \I__6630\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28135\
        );

    \I__6629\ : Odrv12
    port map (
            O => \N__28146\,
            I => uart_pc_data_6
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__28143\,
            I => uart_pc_data_6
        );

    \I__6627\ : Odrv12
    port map (
            O => \N__28138\,
            I => uart_pc_data_6
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__28135\,
            I => uart_pc_data_6
        );

    \I__6625\ : CascadeMux
    port map (
            O => \N__28126\,
            I => \N__28123\
        );

    \I__6624\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28120\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__28120\,
            I => \frame_decoder_OFF3data_6\
        );

    \I__6622\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28110\
        );

    \I__6621\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28107\
        );

    \I__6620\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28102\
        );

    \I__6619\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28099\
        );

    \I__6618\ : InMux
    port map (
            O => \N__28113\,
            I => \N__28095\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__28110\,
            I => \N__28092\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__28107\,
            I => \N__28089\
        );

    \I__6615\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28086\
        );

    \I__6614\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28083\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28080\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28099\,
            I => \N__28077\
        );

    \I__6611\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28073\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__28095\,
            I => \N__28070\
        );

    \I__6609\ : Span4Mux_v
    port map (
            O => \N__28092\,
            I => \N__28065\
        );

    \I__6608\ : Span4Mux_v
    port map (
            O => \N__28089\,
            I => \N__28065\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__28086\,
            I => \N__28060\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__28083\,
            I => \N__28053\
        );

    \I__6605\ : Span4Mux_h
    port map (
            O => \N__28080\,
            I => \N__28053\
        );

    \I__6604\ : Span4Mux_v
    port map (
            O => \N__28077\,
            I => \N__28053\
        );

    \I__6603\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28050\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__28073\,
            I => \N__28045\
        );

    \I__6601\ : Span4Mux_v
    port map (
            O => \N__28070\,
            I => \N__28045\
        );

    \I__6600\ : Span4Mux_h
    port map (
            O => \N__28065\,
            I => \N__28042\
        );

    \I__6599\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28039\
        );

    \I__6598\ : InMux
    port map (
            O => \N__28063\,
            I => \N__28036\
        );

    \I__6597\ : Span12Mux_v
    port map (
            O => \N__28060\,
            I => \N__28033\
        );

    \I__6596\ : Span4Mux_h
    port map (
            O => \N__28053\,
            I => \N__28028\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__28050\,
            I => \N__28028\
        );

    \I__6594\ : Span4Mux_v
    port map (
            O => \N__28045\,
            I => \N__28021\
        );

    \I__6593\ : Span4Mux_h
    port map (
            O => \N__28042\,
            I => \N__28021\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__28039\,
            I => \N__28021\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__28036\,
            I => uart_pc_data_3
        );

    \I__6590\ : Odrv12
    port map (
            O => \N__28033\,
            I => uart_pc_data_3
        );

    \I__6589\ : Odrv4
    port map (
            O => \N__28028\,
            I => uart_pc_data_3
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__28021\,
            I => uart_pc_data_3
        );

    \I__6587\ : CascadeMux
    port map (
            O => \N__28012\,
            I => \N__28009\
        );

    \I__6586\ : InMux
    port map (
            O => \N__28009\,
            I => \N__28006\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__28006\,
            I => \frame_decoder_OFF3data_3\
        );

    \I__6584\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27997\
        );

    \I__6583\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27994\
        );

    \I__6582\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27990\
        );

    \I__6581\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27986\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__27997\,
            I => \N__27981\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__27994\,
            I => \N__27981\
        );

    \I__6578\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27978\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__27990\,
            I => \N__27973\
        );

    \I__6576\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27969\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__27986\,
            I => \N__27964\
        );

    \I__6574\ : Span4Mux_v
    port map (
            O => \N__27981\,
            I => \N__27964\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__27978\,
            I => \N__27961\
        );

    \I__6572\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27958\
        );

    \I__6571\ : CascadeMux
    port map (
            O => \N__27976\,
            I => \N__27953\
        );

    \I__6570\ : Span4Mux_v
    port map (
            O => \N__27973\,
            I => \N__27950\
        );

    \I__6569\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27947\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N__27940\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__27964\,
            I => \N__27940\
        );

    \I__6566\ : Span4Mux_v
    port map (
            O => \N__27961\,
            I => \N__27940\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__27958\,
            I => \N__27937\
        );

    \I__6564\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27934\
        );

    \I__6563\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27931\
        );

    \I__6562\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27928\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__27950\,
            I => \N__27925\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__27947\,
            I => \N__27920\
        );

    \I__6559\ : Span4Mux_h
    port map (
            O => \N__27940\,
            I => \N__27920\
        );

    \I__6558\ : Span4Mux_h
    port map (
            O => \N__27937\,
            I => \N__27917\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__27934\,
            I => \N__27914\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__27931\,
            I => uart_pc_data_4
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__27928\,
            I => uart_pc_data_4
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__27925\,
            I => uart_pc_data_4
        );

    \I__6553\ : Odrv4
    port map (
            O => \N__27920\,
            I => uart_pc_data_4
        );

    \I__6552\ : Odrv4
    port map (
            O => \N__27917\,
            I => uart_pc_data_4
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__27914\,
            I => uart_pc_data_4
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__27901\,
            I => \N__27898\
        );

    \I__6549\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27895\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__27895\,
            I => \frame_decoder_OFF3data_4\
        );

    \I__6547\ : InMux
    port map (
            O => \N__27892\,
            I => \N__27887\
        );

    \I__6546\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27884\
        );

    \I__6545\ : InMux
    port map (
            O => \N__27890\,
            I => \N__27880\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__27887\,
            I => \N__27875\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__27884\,
            I => \N__27875\
        );

    \I__6542\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27872\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__27880\,
            I => \N__27864\
        );

    \I__6540\ : Span4Mux_v
    port map (
            O => \N__27875\,
            I => \N__27864\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__27872\,
            I => \N__27861\
        );

    \I__6538\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27858\
        );

    \I__6537\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27854\
        );

    \I__6536\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27849\
        );

    \I__6535\ : Span4Mux_h
    port map (
            O => \N__27864\,
            I => \N__27842\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__27861\,
            I => \N__27842\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27842\
        );

    \I__6532\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27839\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__27854\,
            I => \N__27836\
        );

    \I__6530\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27833\
        );

    \I__6529\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27830\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__27849\,
            I => \N__27827\
        );

    \I__6527\ : Span4Mux_h
    port map (
            O => \N__27842\,
            I => \N__27820\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__27839\,
            I => \N__27820\
        );

    \I__6525\ : Span4Mux_v
    port map (
            O => \N__27836\,
            I => \N__27813\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__27833\,
            I => \N__27813\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__27830\,
            I => \N__27813\
        );

    \I__6522\ : Span4Mux_v
    port map (
            O => \N__27827\,
            I => \N__27809\
        );

    \I__6521\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27806\
        );

    \I__6520\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27803\
        );

    \I__6519\ : Span4Mux_v
    port map (
            O => \N__27820\,
            I => \N__27800\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__27813\,
            I => \N__27797\
        );

    \I__6517\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27794\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__27809\,
            I => uart_pc_data_5
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__27806\,
            I => uart_pc_data_5
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__27803\,
            I => uart_pc_data_5
        );

    \I__6513\ : Odrv4
    port map (
            O => \N__27800\,
            I => uart_pc_data_5
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__27797\,
            I => uart_pc_data_5
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__27794\,
            I => uart_pc_data_5
        );

    \I__6510\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27778\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__27778\,
            I => \frame_decoder_OFF3data_5\
        );

    \I__6508\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27771\
        );

    \I__6507\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27764\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__27771\,
            I => \N__27760\
        );

    \I__6505\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27757\
        );

    \I__6504\ : CascadeMux
    port map (
            O => \N__27769\,
            I => \N__27754\
        );

    \I__6503\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27751\
        );

    \I__6502\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27748\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__27764\,
            I => \N__27745\
        );

    \I__6500\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27742\
        );

    \I__6499\ : Span4Mux_v
    port map (
            O => \N__27760\,
            I => \N__27737\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__27757\,
            I => \N__27737\
        );

    \I__6497\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27733\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__27751\,
            I => \N__27730\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__27748\,
            I => \N__27727\
        );

    \I__6494\ : Span4Mux_v
    port map (
            O => \N__27745\,
            I => \N__27724\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__27742\,
            I => \N__27719\
        );

    \I__6492\ : Span4Mux_v
    port map (
            O => \N__27737\,
            I => \N__27719\
        );

    \I__6491\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27715\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__27733\,
            I => \N__27710\
        );

    \I__6489\ : Span4Mux_h
    port map (
            O => \N__27730\,
            I => \N__27707\
        );

    \I__6488\ : Span4Mux_h
    port map (
            O => \N__27727\,
            I => \N__27704\
        );

    \I__6487\ : Span4Mux_v
    port map (
            O => \N__27724\,
            I => \N__27699\
        );

    \I__6486\ : Span4Mux_h
    port map (
            O => \N__27719\,
            I => \N__27699\
        );

    \I__6485\ : InMux
    port map (
            O => \N__27718\,
            I => \N__27696\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__27715\,
            I => \N__27693\
        );

    \I__6483\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27690\
        );

    \I__6482\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27687\
        );

    \I__6481\ : Span4Mux_h
    port map (
            O => \N__27710\,
            I => \N__27684\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__27707\,
            I => \N__27679\
        );

    \I__6479\ : Span4Mux_v
    port map (
            O => \N__27704\,
            I => \N__27679\
        );

    \I__6478\ : Span4Mux_h
    port map (
            O => \N__27699\,
            I => \N__27674\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__27696\,
            I => \N__27674\
        );

    \I__6476\ : Span4Mux_h
    port map (
            O => \N__27693\,
            I => \N__27669\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__27690\,
            I => \N__27669\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__27687\,
            I => uart_pc_data_1
        );

    \I__6473\ : Odrv4
    port map (
            O => \N__27684\,
            I => uart_pc_data_1
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__27679\,
            I => uart_pc_data_1
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__27674\,
            I => uart_pc_data_1
        );

    \I__6470\ : Odrv4
    port map (
            O => \N__27669\,
            I => uart_pc_data_1
        );

    \I__6469\ : CascadeMux
    port map (
            O => \N__27658\,
            I => \N__27655\
        );

    \I__6468\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27652\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__27652\,
            I => \frame_decoder_OFF3data_1\
        );

    \I__6466\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27643\
        );

    \I__6465\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27640\
        );

    \I__6464\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27636\
        );

    \I__6463\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27633\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__27643\,
            I => \N__27627\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__27640\,
            I => \N__27627\
        );

    \I__6460\ : InMux
    port map (
            O => \N__27639\,
            I => \N__27624\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__27636\,
            I => \N__27618\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__27633\,
            I => \N__27614\
        );

    \I__6457\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27611\
        );

    \I__6456\ : Span4Mux_v
    port map (
            O => \N__27627\,
            I => \N__27606\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__27624\,
            I => \N__27606\
        );

    \I__6454\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27602\
        );

    \I__6453\ : InMux
    port map (
            O => \N__27622\,
            I => \N__27599\
        );

    \I__6452\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27596\
        );

    \I__6451\ : Span4Mux_v
    port map (
            O => \N__27618\,
            I => \N__27593\
        );

    \I__6450\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27590\
        );

    \I__6449\ : Span4Mux_v
    port map (
            O => \N__27614\,
            I => \N__27587\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__27611\,
            I => \N__27584\
        );

    \I__6447\ : Span4Mux_v
    port map (
            O => \N__27606\,
            I => \N__27581\
        );

    \I__6446\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27578\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__27602\,
            I => \N__27572\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__27599\,
            I => \N__27572\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__27596\,
            I => \N__27569\
        );

    \I__6442\ : Span4Mux_v
    port map (
            O => \N__27593\,
            I => \N__27564\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__27590\,
            I => \N__27564\
        );

    \I__6440\ : Sp12to4
    port map (
            O => \N__27587\,
            I => \N__27555\
        );

    \I__6439\ : Span12Mux_v
    port map (
            O => \N__27584\,
            I => \N__27555\
        );

    \I__6438\ : Sp12to4
    port map (
            O => \N__27581\,
            I => \N__27555\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__27578\,
            I => \N__27555\
        );

    \I__6436\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27552\
        );

    \I__6435\ : Span4Mux_h
    port map (
            O => \N__27572\,
            I => \N__27549\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__27569\,
            I => \N__27544\
        );

    \I__6433\ : Span4Mux_h
    port map (
            O => \N__27564\,
            I => \N__27544\
        );

    \I__6432\ : Odrv12
    port map (
            O => \N__27555\,
            I => uart_pc_data_7
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__27552\,
            I => uart_pc_data_7
        );

    \I__6430\ : Odrv4
    port map (
            O => \N__27549\,
            I => uart_pc_data_7
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__27544\,
            I => uart_pc_data_7
        );

    \I__6428\ : CascadeMux
    port map (
            O => \N__27535\,
            I => \N__27532\
        );

    \I__6427\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27526\
        );

    \I__6426\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27526\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__27526\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__6424\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27520\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__27520\,
            I => \scaler_3.N_533_i_l_ofxZ0\
        );

    \I__6422\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27512\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__27516\,
            I => \N__27509\
        );

    \I__6420\ : InMux
    port map (
            O => \N__27515\,
            I => \N__27505\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__27512\,
            I => \N__27502\
        );

    \I__6418\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27497\
        );

    \I__6417\ : InMux
    port map (
            O => \N__27508\,
            I => \N__27497\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__27505\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__6415\ : Odrv12
    port map (
            O => \N__27502\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__27497\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__6413\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27484\
        );

    \I__6412\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27481\
        );

    \I__6411\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27478\
        );

    \I__6410\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27475\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__27484\,
            I => \N__27470\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__27481\,
            I => \N__27470\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__27478\,
            I => \N__27465\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__27475\,
            I => \N__27465\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__27470\,
            I => \N__27462\
        );

    \I__6404\ : Span4Mux_v
    port map (
            O => \N__27465\,
            I => \N__27459\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__27462\,
            I => \frame_decoder_CH3data_0\
        );

    \I__6402\ : Odrv4
    port map (
            O => \N__27459\,
            I => \frame_decoder_CH3data_0\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__27454\,
            I => \N__27451\
        );

    \I__6400\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27448\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__27448\,
            I => \scaler_3.un2_source_data_0_cry_1_c_RNO_0\
        );

    \I__6398\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27442\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__27442\,
            I => \scaler_3.un3_source_data_0_axb_7\
        );

    \I__6396\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27436\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27433\
        );

    \I__6394\ : Odrv4
    port map (
            O => \N__27433\,
            I => \frame_decoder_CH3data_1\
        );

    \I__6393\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27424\
        );

    \I__6392\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27424\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__27424\,
            I => \frame_decoder_CH3data_7\
        );

    \I__6390\ : CEMux
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__27418\,
            I => \N__27414\
        );

    \I__6388\ : CEMux
    port map (
            O => \N__27417\,
            I => \N__27411\
        );

    \I__6387\ : Span4Mux_v
    port map (
            O => \N__27414\,
            I => \N__27408\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__27411\,
            I => \N__27405\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__27408\,
            I => \N__27401\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__27405\,
            I => \N__27398\
        );

    \I__6383\ : CEMux
    port map (
            O => \N__27404\,
            I => \N__27395\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__27401\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6381\ : Odrv4
    port map (
            O => \N__27398\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__27395\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__27388\,
            I => \N__27384\
        );

    \I__6378\ : InMux
    port map (
            O => \N__27387\,
            I => \N__27381\
        );

    \I__6377\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27378\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__27381\,
            I => \N__27375\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__27378\,
            I => \N__27371\
        );

    \I__6374\ : Span4Mux_v
    port map (
            O => \N__27375\,
            I => \N__27368\
        );

    \I__6373\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27365\
        );

    \I__6372\ : Span4Mux_h
    port map (
            O => \N__27371\,
            I => \N__27362\
        );

    \I__6371\ : Odrv4
    port map (
            O => \N__27368\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__27365\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__27362\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__6368\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27352\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__27352\,
            I => \Commands_frame_decoder.count_1_sqmuxa\
        );

    \I__6366\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27343\
        );

    \I__6365\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27338\
        );

    \I__6364\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27338\
        );

    \I__6363\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27334\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__27343\,
            I => \N__27329\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__27338\,
            I => \N__27329\
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__27337\,
            I => \N__27326\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__27334\,
            I => \N__27323\
        );

    \I__6358\ : Span4Mux_h
    port map (
            O => \N__27329\,
            I => \N__27320\
        );

    \I__6357\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27317\
        );

    \I__6356\ : Span12Mux_v
    port map (
            O => \N__27323\,
            I => \N__27314\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__27320\,
            I => pc_frame_decoder_dv
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__27317\,
            I => pc_frame_decoder_dv
        );

    \I__6353\ : Odrv12
    port map (
            O => \N__27314\,
            I => pc_frame_decoder_dv
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__27307\,
            I => \N__27303\
        );

    \I__6351\ : CascadeMux
    port map (
            O => \N__27306\,
            I => \N__27300\
        );

    \I__6350\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27292\
        );

    \I__6349\ : InMux
    port map (
            O => \N__27300\,
            I => \N__27289\
        );

    \I__6348\ : CascadeMux
    port map (
            O => \N__27299\,
            I => \N__27286\
        );

    \I__6347\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27283\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__27297\,
            I => \N__27280\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__27296\,
            I => \N__27277\
        );

    \I__6344\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27261\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__27292\,
            I => \N__27258\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27255\
        );

    \I__6341\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27252\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__27283\,
            I => \N__27249\
        );

    \I__6339\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27246\
        );

    \I__6338\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27243\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__27276\,
            I => \N__27240\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__27275\,
            I => \N__27237\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__27274\,
            I => \N__27234\
        );

    \I__6334\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27231\
        );

    \I__6333\ : CascadeMux
    port map (
            O => \N__27272\,
            I => \N__27228\
        );

    \I__6332\ : CascadeMux
    port map (
            O => \N__27271\,
            I => \N__27225\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__27270\,
            I => \N__27222\
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__27269\,
            I => \N__27219\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__27268\,
            I => \N__27216\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__27267\,
            I => \N__27213\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__27266\,
            I => \N__27210\
        );

    \I__6326\ : CascadeMux
    port map (
            O => \N__27265\,
            I => \N__27203\
        );

    \I__6325\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27200\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__27261\,
            I => \N__27197\
        );

    \I__6323\ : Span4Mux_h
    port map (
            O => \N__27258\,
            I => \N__27194\
        );

    \I__6322\ : Span4Mux_v
    port map (
            O => \N__27255\,
            I => \N__27189\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__27252\,
            I => \N__27189\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__27249\,
            I => \N__27182\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__27246\,
            I => \N__27182\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__27243\,
            I => \N__27182\
        );

    \I__6317\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27179\
        );

    \I__6316\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27176\
        );

    \I__6315\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27173\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__27231\,
            I => \N__27170\
        );

    \I__6313\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27161\
        );

    \I__6312\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27161\
        );

    \I__6311\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27161\
        );

    \I__6310\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27161\
        );

    \I__6309\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27154\
        );

    \I__6308\ : InMux
    port map (
            O => \N__27213\,
            I => \N__27154\
        );

    \I__6307\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27154\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__27209\,
            I => \N__27151\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__27208\,
            I => \N__27148\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__27207\,
            I => \N__27145\
        );

    \I__6303\ : CascadeMux
    port map (
            O => \N__27206\,
            I => \N__27142\
        );

    \I__6302\ : InMux
    port map (
            O => \N__27203\,
            I => \N__27139\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__27200\,
            I => \N__27136\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__27197\,
            I => \N__27133\
        );

    \I__6299\ : Span4Mux_v
    port map (
            O => \N__27194\,
            I => \N__27124\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__27189\,
            I => \N__27124\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__27182\,
            I => \N__27124\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__27179\,
            I => \N__27124\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__27176\,
            I => \N__27119\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__27173\,
            I => \N__27119\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__27170\,
            I => \N__27116\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__27161\,
            I => \N__27111\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__27154\,
            I => \N__27111\
        );

    \I__6290\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27108\
        );

    \I__6289\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27103\
        );

    \I__6288\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27103\
        );

    \I__6287\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27100\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__27139\,
            I => \N__27097\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__27136\,
            I => \N__27094\
        );

    \I__6284\ : Span4Mux_v
    port map (
            O => \N__27133\,
            I => \N__27091\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__27124\,
            I => \N__27088\
        );

    \I__6282\ : Span4Mux_s3_v
    port map (
            O => \N__27119\,
            I => \N__27085\
        );

    \I__6281\ : Span4Mux_v
    port map (
            O => \N__27116\,
            I => \N__27082\
        );

    \I__6280\ : Span4Mux_h
    port map (
            O => \N__27111\,
            I => \N__27079\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__27108\,
            I => \N__27072\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__27103\,
            I => \N__27072\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27072\
        );

    \I__6276\ : Span12Mux_v
    port map (
            O => \N__27097\,
            I => \N__27069\
        );

    \I__6275\ : Sp12to4
    port map (
            O => \N__27094\,
            I => \N__27066\
        );

    \I__6274\ : Span4Mux_v
    port map (
            O => \N__27091\,
            I => \N__27059\
        );

    \I__6273\ : Span4Mux_v
    port map (
            O => \N__27088\,
            I => \N__27059\
        );

    \I__6272\ : Span4Mux_v
    port map (
            O => \N__27085\,
            I => \N__27059\
        );

    \I__6271\ : Span4Mux_h
    port map (
            O => \N__27082\,
            I => \N__27052\
        );

    \I__6270\ : Span4Mux_v
    port map (
            O => \N__27079\,
            I => \N__27052\
        );

    \I__6269\ : Span4Mux_v
    port map (
            O => \N__27072\,
            I => \N__27052\
        );

    \I__6268\ : Odrv12
    port map (
            O => \N__27069\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6267\ : Odrv12
    port map (
            O => \N__27066\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6266\ : Odrv4
    port map (
            O => \N__27059\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6265\ : Odrv4
    port map (
            O => \N__27052\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6264\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27039\
        );

    \I__6263\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27036\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__27039\,
            I => \Commands_frame_decoder.count8_0_i\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__27036\,
            I => \Commands_frame_decoder.count8_0_i\
        );

    \I__6260\ : InMux
    port map (
            O => \N__27031\,
            I => \N__27027\
        );

    \I__6259\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27024\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__27027\,
            I => \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__27024\,
            I => \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0\
        );

    \I__6256\ : InMux
    port map (
            O => \N__27019\,
            I => \N__27014\
        );

    \I__6255\ : InMux
    port map (
            O => \N__27018\,
            I => \N__27009\
        );

    \I__6254\ : InMux
    port map (
            O => \N__27017\,
            I => \N__27009\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__27014\,
            I => \Commands_frame_decoder.state_1_ns_i_a4_2_0_0\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__27009\,
            I => \Commands_frame_decoder.state_1_ns_i_a4_2_0_0\
        );

    \I__6251\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26998\
        );

    \I__6250\ : InMux
    port map (
            O => \N__27003\,
            I => \N__26995\
        );

    \I__6249\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26990\
        );

    \I__6248\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26990\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__26998\,
            I => \Commands_frame_decoder.count8_0\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__26995\,
            I => \Commands_frame_decoder.count8_0\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__26990\,
            I => \Commands_frame_decoder.count8_0\
        );

    \I__6244\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26980\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__26980\,
            I => \frame_decoder_CH3data_2\
        );

    \I__6242\ : CascadeMux
    port map (
            O => \N__26977\,
            I => \N__26974\
        );

    \I__6241\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26968\
        );

    \I__6240\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26968\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__26968\,
            I => \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\
        );

    \I__6238\ : InMux
    port map (
            O => \N__26965\,
            I => \scaler_3.un3_source_data_0_cry_1\
        );

    \I__6237\ : InMux
    port map (
            O => \N__26962\,
            I => \N__26959\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__26959\,
            I => \frame_decoder_CH3data_3\
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__26956\,
            I => \N__26953\
        );

    \I__6234\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26947\
        );

    \I__6233\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26947\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__26947\,
            I => \scaler_3.un3_source_data_0_cry_2_c_RNI780L\
        );

    \I__6231\ : InMux
    port map (
            O => \N__26944\,
            I => \scaler_3.un3_source_data_0_cry_2\
        );

    \I__6230\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26938\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__26938\,
            I => \frame_decoder_CH3data_4\
        );

    \I__6228\ : CascadeMux
    port map (
            O => \N__26935\,
            I => \N__26932\
        );

    \I__6227\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26926\
        );

    \I__6226\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26926\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__26926\,
            I => \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\
        );

    \I__6224\ : InMux
    port map (
            O => \N__26923\,
            I => \scaler_3.un3_source_data_0_cry_3\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__26920\,
            I => \N__26917\
        );

    \I__6222\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26914\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__26914\,
            I => \frame_decoder_CH3data_5\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__6219\ : InMux
    port map (
            O => \N__26908\,
            I => \N__26902\
        );

    \I__6218\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26902\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__26902\,
            I => \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\
        );

    \I__6216\ : InMux
    port map (
            O => \N__26899\,
            I => \scaler_3.un3_source_data_0_cry_4\
        );

    \I__6215\ : InMux
    port map (
            O => \N__26896\,
            I => \N__26893\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__26893\,
            I => \frame_decoder_CH3data_6\
        );

    \I__6213\ : CascadeMux
    port map (
            O => \N__26890\,
            I => \N__26887\
        );

    \I__6212\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26881\
        );

    \I__6211\ : InMux
    port map (
            O => \N__26886\,
            I => \N__26881\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__26881\,
            I => \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\
        );

    \I__6209\ : InMux
    port map (
            O => \N__26878\,
            I => \scaler_3.un3_source_data_0_cry_5\
        );

    \I__6208\ : CascadeMux
    port map (
            O => \N__26875\,
            I => \N__26872\
        );

    \I__6207\ : InMux
    port map (
            O => \N__26872\,
            I => \N__26866\
        );

    \I__6206\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26866\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__26866\,
            I => \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\
        );

    \I__6204\ : InMux
    port map (
            O => \N__26863\,
            I => \scaler_3.un3_source_data_0_cry_6\
        );

    \I__6203\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26856\
        );

    \I__6202\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26853\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__26856\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__26853\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\
        );

    \I__6199\ : InMux
    port map (
            O => \N__26848\,
            I => \bfn_12_16_0_\
        );

    \I__6198\ : InMux
    port map (
            O => \N__26845\,
            I => \scaler_3.un3_source_data_0_cry_8\
        );

    \I__6197\ : CascadeMux
    port map (
            O => \N__26842\,
            I => \N__26839\
        );

    \I__6196\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26836\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__26836\,
            I => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\
        );

    \I__6194\ : IoInMux
    port map (
            O => \N__26833\,
            I => \N__26830\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__26830\,
            I => \N__26827\
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__26827\,
            I => pc_frame_decoder_dv_0
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__26824\,
            I => \N__26821\
        );

    \I__6190\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26818\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__26818\,
            I => \N__26815\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__26815\,
            I => \frame_decoder_CH4data_1\
        );

    \I__6187\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26807\
        );

    \I__6186\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26804\
        );

    \I__6185\ : InMux
    port map (
            O => \N__26810\,
            I => \N__26801\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__26807\,
            I => \N__26794\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__26804\,
            I => \N__26794\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26794\
        );

    \I__6181\ : Span4Mux_v
    port map (
            O => \N__26794\,
            I => \N__26790\
        );

    \I__6180\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26787\
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__26790\,
            I => \frame_decoder_CH4data_0\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__26787\,
            I => \frame_decoder_CH4data_0\
        );

    \I__6177\ : CEMux
    port map (
            O => \N__26782\,
            I => \N__26778\
        );

    \I__6176\ : CEMux
    port map (
            O => \N__26781\,
            I => \N__26775\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__26778\,
            I => \N__26770\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__26775\,
            I => \N__26767\
        );

    \I__6173\ : CEMux
    port map (
            O => \N__26774\,
            I => \N__26764\
        );

    \I__6172\ : CEMux
    port map (
            O => \N__26773\,
            I => \N__26761\
        );

    \I__6171\ : Span4Mux_v
    port map (
            O => \N__26770\,
            I => \N__26754\
        );

    \I__6170\ : Span4Mux_h
    port map (
            O => \N__26767\,
            I => \N__26754\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__26764\,
            I => \N__26754\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__26761\,
            I => \N__26751\
        );

    \I__6167\ : Span4Mux_h
    port map (
            O => \N__26754\,
            I => \N__26748\
        );

    \I__6166\ : Span4Mux_v
    port map (
            O => \N__26751\,
            I => \N__26745\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__26748\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__6164\ : Odrv4
    port map (
            O => \N__26745\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__6163\ : InMux
    port map (
            O => \N__26740\,
            I => \scaler_3.un3_source_data_0_cry_0\
        );

    \I__6162\ : InMux
    port map (
            O => \N__26737\,
            I => \N__26734\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__26734\,
            I => \N__26731\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__26731\,
            I => \uart_drone.CO0\
        );

    \I__6159\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26725\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__26725\,
            I => \Commands_frame_decoder.count8_axb_1\
        );

    \I__6157\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26719\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__26719\,
            I => \Commands_frame_decoder.count_i_2\
        );

    \I__6155\ : InMux
    port map (
            O => \N__26716\,
            I => \Commands_frame_decoder.count8\
        );

    \I__6154\ : InMux
    port map (
            O => \N__26713\,
            I => \N__26710\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__26710\,
            I => \Commands_frame_decoder.count8_THRU_CO\
        );

    \I__6152\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26704\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__26704\,
            I => \N__26701\
        );

    \I__6150\ : Span4Mux_v
    port map (
            O => \N__26701\,
            I => \N__26698\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__26698\,
            I => \N__26688\
        );

    \I__6148\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26680\
        );

    \I__6147\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26676\
        );

    \I__6146\ : InMux
    port map (
            O => \N__26695\,
            I => \N__26671\
        );

    \I__6145\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26671\
        );

    \I__6144\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26664\
        );

    \I__6143\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26664\
        );

    \I__6142\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26664\
        );

    \I__6141\ : Span4Mux_v
    port map (
            O => \N__26688\,
            I => \N__26661\
        );

    \I__6140\ : InMux
    port map (
            O => \N__26687\,
            I => \N__26658\
        );

    \I__6139\ : InMux
    port map (
            O => \N__26686\,
            I => \N__26648\
        );

    \I__6138\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26648\
        );

    \I__6137\ : InMux
    port map (
            O => \N__26684\,
            I => \N__26648\
        );

    \I__6136\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26648\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__26680\,
            I => \N__26643\
        );

    \I__6134\ : IoInMux
    port map (
            O => \N__26679\,
            I => \N__26639\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__26676\,
            I => \N__26632\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__26671\,
            I => \N__26632\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__26664\,
            I => \N__26632\
        );

    \I__6130\ : Span4Mux_h
    port map (
            O => \N__26661\,
            I => \N__26627\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__26658\,
            I => \N__26627\
        );

    \I__6128\ : InMux
    port map (
            O => \N__26657\,
            I => \N__26618\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__26648\,
            I => \N__26615\
        );

    \I__6126\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26612\
        );

    \I__6125\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26609\
        );

    \I__6124\ : Span4Mux_h
    port map (
            O => \N__26643\,
            I => \N__26605\
        );

    \I__6123\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26602\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__26639\,
            I => \N__26599\
        );

    \I__6121\ : Span4Mux_v
    port map (
            O => \N__26632\,
            I => \N__26596\
        );

    \I__6120\ : Span4Mux_v
    port map (
            O => \N__26627\,
            I => \N__26593\
        );

    \I__6119\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26590\
        );

    \I__6118\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26585\
        );

    \I__6117\ : InMux
    port map (
            O => \N__26624\,
            I => \N__26585\
        );

    \I__6116\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26578\
        );

    \I__6115\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26578\
        );

    \I__6114\ : InMux
    port map (
            O => \N__26621\,
            I => \N__26578\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__26618\,
            I => \N__26575\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__26615\,
            I => \N__26568\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__26612\,
            I => \N__26568\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__26609\,
            I => \N__26568\
        );

    \I__6109\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26565\
        );

    \I__6108\ : Sp12to4
    port map (
            O => \N__26605\,
            I => \N__26560\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__26602\,
            I => \N__26560\
        );

    \I__6106\ : Span4Mux_s1_v
    port map (
            O => \N__26599\,
            I => \N__26557\
        );

    \I__6105\ : Span4Mux_v
    port map (
            O => \N__26596\,
            I => \N__26552\
        );

    \I__6104\ : Span4Mux_v
    port map (
            O => \N__26593\,
            I => \N__26552\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__26590\,
            I => \N__26537\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__26585\,
            I => \N__26537\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26537\
        );

    \I__6100\ : Span12Mux_h
    port map (
            O => \N__26575\,
            I => \N__26537\
        );

    \I__6099\ : Sp12to4
    port map (
            O => \N__26568\,
            I => \N__26537\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__26565\,
            I => \N__26537\
        );

    \I__6097\ : Span12Mux_s11_v
    port map (
            O => \N__26560\,
            I => \N__26537\
        );

    \I__6096\ : Span4Mux_v
    port map (
            O => \N__26557\,
            I => \N__26534\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__26552\,
            I => reset_system
        );

    \I__6094\ : Odrv12
    port map (
            O => \N__26537\,
            I => reset_system
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__26534\,
            I => reset_system
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__26527\,
            I => \Commands_frame_decoder.count8_THRU_CO_cascade_\
        );

    \I__6091\ : CascadeMux
    port map (
            O => \N__26524\,
            I => \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0_cascade_\
        );

    \I__6090\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26516\
        );

    \I__6089\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26511\
        );

    \I__6088\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26511\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__26516\,
            I => \Commands_frame_decoder.countZ0Z_2\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__26511\,
            I => \Commands_frame_decoder.countZ0Z_2\
        );

    \I__6085\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26503\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__26503\,
            I => \Commands_frame_decoder.CO0\
        );

    \I__6083\ : CascadeMux
    port map (
            O => \N__26500\,
            I => \Commands_frame_decoder.CO0_cascade_\
        );

    \I__6082\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26491\
        );

    \I__6081\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26484\
        );

    \I__6080\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26484\
        );

    \I__6079\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26484\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__26491\,
            I => \Commands_frame_decoder.countZ0Z_1\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__26484\,
            I => \Commands_frame_decoder.countZ0Z_1\
        );

    \I__6076\ : InMux
    port map (
            O => \N__26479\,
            I => \N__26475\
        );

    \I__6075\ : InMux
    port map (
            O => \N__26478\,
            I => \N__26472\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__26475\,
            I => \N__26469\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__26472\,
            I => \N__26466\
        );

    \I__6072\ : Span12Mux_v
    port map (
            O => \N__26469\,
            I => \N__26463\
        );

    \I__6071\ : Span4Mux_h
    port map (
            O => \N__26466\,
            I => \N__26460\
        );

    \I__6070\ : Odrv12
    port map (
            O => \N__26463\,
            I => scaler_3_data_11
        );

    \I__6069\ : Odrv4
    port map (
            O => \N__26460\,
            I => scaler_3_data_11
        );

    \I__6068\ : InMux
    port map (
            O => \N__26455\,
            I => \scaler_3.un2_source_data_0_cry_6\
        );

    \I__6067\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26448\
        );

    \I__6066\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26445\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__26448\,
            I => \N__26442\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26439\
        );

    \I__6063\ : Span12Mux_v
    port map (
            O => \N__26442\,
            I => \N__26436\
        );

    \I__6062\ : Span4Mux_h
    port map (
            O => \N__26439\,
            I => \N__26433\
        );

    \I__6061\ : Odrv12
    port map (
            O => \N__26436\,
            I => scaler_3_data_12
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__26433\,
            I => scaler_3_data_12
        );

    \I__6059\ : InMux
    port map (
            O => \N__26428\,
            I => \scaler_3.un2_source_data_0_cry_7\
        );

    \I__6058\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26422\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__26422\,
            I => \N__26418\
        );

    \I__6056\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26415\
        );

    \I__6055\ : Span4Mux_h
    port map (
            O => \N__26418\,
            I => \N__26412\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__26415\,
            I => \N__26409\
        );

    \I__6053\ : Span4Mux_v
    port map (
            O => \N__26412\,
            I => \N__26406\
        );

    \I__6052\ : Span4Mux_h
    port map (
            O => \N__26409\,
            I => \N__26403\
        );

    \I__6051\ : Odrv4
    port map (
            O => \N__26406\,
            I => scaler_3_data_13
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__26403\,
            I => scaler_3_data_13
        );

    \I__6049\ : InMux
    port map (
            O => \N__26398\,
            I => \bfn_11_17_0_\
        );

    \I__6048\ : InMux
    port map (
            O => \N__26395\,
            I => \scaler_3.un2_source_data_0_cry_9\
        );

    \I__6047\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26389\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__26389\,
            I => \N__26386\
        );

    \I__6045\ : Span4Mux_v
    port map (
            O => \N__26386\,
            I => \N__26383\
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__26383\,
            I => scaler_3_data_14
        );

    \I__6043\ : CEMux
    port map (
            O => \N__26380\,
            I => \N__26359\
        );

    \I__6042\ : CEMux
    port map (
            O => \N__26379\,
            I => \N__26359\
        );

    \I__6041\ : CEMux
    port map (
            O => \N__26378\,
            I => \N__26359\
        );

    \I__6040\ : CEMux
    port map (
            O => \N__26377\,
            I => \N__26359\
        );

    \I__6039\ : CEMux
    port map (
            O => \N__26376\,
            I => \N__26359\
        );

    \I__6038\ : CEMux
    port map (
            O => \N__26375\,
            I => \N__26359\
        );

    \I__6037\ : CEMux
    port map (
            O => \N__26374\,
            I => \N__26359\
        );

    \I__6036\ : GlobalMux
    port map (
            O => \N__26359\,
            I => \N__26356\
        );

    \I__6035\ : gio2CtrlBuf
    port map (
            O => \N__26356\,
            I => pc_frame_decoder_dv_0_g
        );

    \I__6034\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26350\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__26350\,
            I => \N__26345\
        );

    \I__6032\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26342\
        );

    \I__6031\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26337\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__26345\,
            I => \N__26329\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__26342\,
            I => \N__26329\
        );

    \I__6028\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26326\
        );

    \I__6027\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26323\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__26337\,
            I => \N__26320\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \N__26317\
        );

    \I__6024\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26314\
        );

    \I__6023\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26310\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__26329\,
            I => \N__26301\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__26326\,
            I => \N__26301\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__26323\,
            I => \N__26301\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__26320\,
            I => \N__26301\
        );

    \I__6018\ : InMux
    port map (
            O => \N__26317\,
            I => \N__26298\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__26314\,
            I => \N__26295\
        );

    \I__6016\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26292\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__26310\,
            I => \N__26287\
        );

    \I__6014\ : Span4Mux_v
    port map (
            O => \N__26301\,
            I => \N__26287\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__26298\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6012\ : Odrv12
    port map (
            O => \N__26295\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__26292\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6010\ : Odrv4
    port map (
            O => \N__26287\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__6009\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26275\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__26275\,
            I => \N__26268\
        );

    \I__6007\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26265\
        );

    \I__6006\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26260\
        );

    \I__6005\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26257\
        );

    \I__6004\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26254\
        );

    \I__6003\ : Span4Mux_h
    port map (
            O => \N__26268\,
            I => \N__26247\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__26265\,
            I => \N__26247\
        );

    \I__6001\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26244\
        );

    \I__6000\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26240\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__26260\,
            I => \N__26233\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__26257\,
            I => \N__26233\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26233\
        );

    \I__5996\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26228\
        );

    \I__5995\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26228\
        );

    \I__5994\ : Sp12to4
    port map (
            O => \N__26247\,
            I => \N__26223\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__26244\,
            I => \N__26223\
        );

    \I__5992\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26220\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__26240\,
            I => \N__26215\
        );

    \I__5990\ : Span12Mux_v
    port map (
            O => \N__26233\,
            I => \N__26215\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__26228\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5988\ : Odrv12
    port map (
            O => \N__26223\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__26220\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5986\ : Odrv12
    port map (
            O => \N__26215\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5985\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26203\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__26203\,
            I => \N__26200\
        );

    \I__5983\ : Span4Mux_h
    port map (
            O => \N__26200\,
            I => \N__26197\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__26197\,
            I => \uart_drone.data_Auxce_0_1\
        );

    \I__5981\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26188\
        );

    \I__5980\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26188\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__26188\,
            I => \N__26185\
        );

    \I__5978\ : Span4Mux_h
    port map (
            O => \N__26185\,
            I => \N__26180\
        );

    \I__5977\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26175\
        );

    \I__5976\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26175\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__26180\,
            I => \Commands_frame_decoder.state_1Z0Z_10\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__26175\,
            I => \Commands_frame_decoder.state_1Z0Z_10\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__26170\,
            I => \Commands_frame_decoder.state_1_ns_i_a4_2_0_0_cascade_\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__26167\,
            I => \N__26164\
        );

    \I__5971\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26158\
        );

    \I__5970\ : InMux
    port map (
            O => \N__26163\,
            I => \N__26158\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__26158\,
            I => \N__26155\
        );

    \I__5968\ : Span4Mux_h
    port map (
            O => \N__26155\,
            I => \N__26152\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__26152\,
            I => \Commands_frame_decoder.N_292\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__26149\,
            I => \N__26144\
        );

    \I__5965\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26141\
        );

    \I__5964\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26138\
        );

    \I__5963\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26134\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__26141\,
            I => \N__26131\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__26138\,
            I => \N__26128\
        );

    \I__5960\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26125\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__26134\,
            I => \N__26116\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__26131\,
            I => \N__26116\
        );

    \I__5957\ : Span4Mux_h
    port map (
            O => \N__26128\,
            I => \N__26116\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__26125\,
            I => \N__26116\
        );

    \I__5955\ : Odrv4
    port map (
            O => \N__26116\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__5954\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26105\
        );

    \I__5953\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26102\
        );

    \I__5952\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26099\
        );

    \I__5951\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26096\
        );

    \I__5950\ : InMux
    port map (
            O => \N__26109\,
            I => \N__26091\
        );

    \I__5949\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26087\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__26105\,
            I => \N__26082\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26082\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__26099\,
            I => \N__26077\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__26096\,
            I => \N__26077\
        );

    \I__5944\ : InMux
    port map (
            O => \N__26095\,
            I => \N__26074\
        );

    \I__5943\ : InMux
    port map (
            O => \N__26094\,
            I => \N__26069\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__26091\,
            I => \N__26066\
        );

    \I__5941\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26063\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__26087\,
            I => \N__26058\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__26082\,
            I => \N__26058\
        );

    \I__5938\ : Span4Mux_v
    port map (
            O => \N__26077\,
            I => \N__26053\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__26074\,
            I => \N__26053\
        );

    \I__5936\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26048\
        );

    \I__5935\ : InMux
    port map (
            O => \N__26072\,
            I => \N__26048\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__26069\,
            I => \N__26043\
        );

    \I__5933\ : Span4Mux_h
    port map (
            O => \N__26066\,
            I => \N__26043\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__26063\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__26058\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__5930\ : Odrv4
    port map (
            O => \N__26053\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__26048\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__5928\ : Odrv4
    port map (
            O => \N__26043\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__5927\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__26029\,
            I => \N__26026\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__26026\,
            I => \scaler_4.N_545_i_l_ofxZ0\
        );

    \I__5924\ : InMux
    port map (
            O => \N__26023\,
            I => \N__26019\
        );

    \I__5923\ : InMux
    port map (
            O => \N__26022\,
            I => \N__26016\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__26019\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__26016\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__5920\ : InMux
    port map (
            O => \N__26011\,
            I => \bfn_11_15_0_\
        );

    \I__5919\ : InMux
    port map (
            O => \N__26008\,
            I => \scaler_4.un3_source_data_0_cry_8\
        );

    \I__5918\ : CascadeMux
    port map (
            O => \N__26005\,
            I => \N__26002\
        );

    \I__5917\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25999\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__25999\,
            I => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\
        );

    \I__5915\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25993\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__5913\ : Span4Mux_v
    port map (
            O => \N__25990\,
            I => \N__25987\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__25987\,
            I => \N__25983\
        );

    \I__5911\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25980\
        );

    \I__5910\ : Span4Mux_h
    port map (
            O => \N__25983\,
            I => \N__25975\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__25980\,
            I => \N__25975\
        );

    \I__5908\ : Span4Mux_v
    port map (
            O => \N__25975\,
            I => \N__25972\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__25972\,
            I => scaler_3_data_6
        );

    \I__5906\ : InMux
    port map (
            O => \N__25969\,
            I => \scaler_3.un2_source_data_0_cry_1\
        );

    \I__5905\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25963\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__25963\,
            I => \N__25960\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__25960\,
            I => \N__25956\
        );

    \I__5902\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25953\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__25956\,
            I => \N__25948\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__25953\,
            I => \N__25948\
        );

    \I__5899\ : Span4Mux_h
    port map (
            O => \N__25948\,
            I => \N__25945\
        );

    \I__5898\ : Odrv4
    port map (
            O => \N__25945\,
            I => scaler_3_data_7
        );

    \I__5897\ : InMux
    port map (
            O => \N__25942\,
            I => \scaler_3.un2_source_data_0_cry_2\
        );

    \I__5896\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25936\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__25936\,
            I => \N__25932\
        );

    \I__5894\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25929\
        );

    \I__5893\ : Span4Mux_v
    port map (
            O => \N__25932\,
            I => \N__25924\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__25929\,
            I => \N__25924\
        );

    \I__5891\ : Span4Mux_h
    port map (
            O => \N__25924\,
            I => \N__25921\
        );

    \I__5890\ : Odrv4
    port map (
            O => \N__25921\,
            I => scaler_3_data_8
        );

    \I__5889\ : InMux
    port map (
            O => \N__25918\,
            I => \scaler_3.un2_source_data_0_cry_3\
        );

    \I__5888\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25912\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25908\
        );

    \I__5886\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25905\
        );

    \I__5885\ : Span4Mux_v
    port map (
            O => \N__25908\,
            I => \N__25902\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__25905\,
            I => \N__25899\
        );

    \I__5883\ : Span4Mux_h
    port map (
            O => \N__25902\,
            I => \N__25894\
        );

    \I__5882\ : Span4Mux_h
    port map (
            O => \N__25899\,
            I => \N__25894\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__25894\,
            I => scaler_3_data_9
        );

    \I__5880\ : InMux
    port map (
            O => \N__25891\,
            I => \scaler_3.un2_source_data_0_cry_4\
        );

    \I__5879\ : InMux
    port map (
            O => \N__25888\,
            I => \N__25884\
        );

    \I__5878\ : InMux
    port map (
            O => \N__25887\,
            I => \N__25881\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__25884\,
            I => \N__25878\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__25881\,
            I => \N__25875\
        );

    \I__5875\ : Span12Mux_s11_h
    port map (
            O => \N__25878\,
            I => \N__25872\
        );

    \I__5874\ : Span4Mux_h
    port map (
            O => \N__25875\,
            I => \N__25869\
        );

    \I__5873\ : Odrv12
    port map (
            O => \N__25872\,
            I => scaler_3_data_10
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__25869\,
            I => scaler_3_data_10
        );

    \I__5871\ : InMux
    port map (
            O => \N__25864\,
            I => \scaler_3.un2_source_data_0_cry_5\
        );

    \I__5870\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25857\
        );

    \I__5869\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25853\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__25857\,
            I => \N__25849\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__25856\,
            I => \N__25846\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__25853\,
            I => \N__25843\
        );

    \I__5865\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25840\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__25849\,
            I => \N__25837\
        );

    \I__5863\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25834\
        );

    \I__5862\ : Odrv4
    port map (
            O => \N__25843\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__25840\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__25837\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__25834\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5858\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25822\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__25822\,
            I => \frame_decoder_OFF4data_1\
        );

    \I__5856\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25815\
        );

    \I__5855\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25812\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__25815\,
            I => \N__25806\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__25812\,
            I => \N__25806\
        );

    \I__5852\ : CascadeMux
    port map (
            O => \N__25811\,
            I => \N__25803\
        );

    \I__5851\ : Span4Mux_h
    port map (
            O => \N__25806\,
            I => \N__25799\
        );

    \I__5850\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25794\
        );

    \I__5849\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25794\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__25799\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__25794\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__5846\ : InMux
    port map (
            O => \N__25789\,
            I => \scaler_4.un3_source_data_0_cry_0\
        );

    \I__5845\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25783\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__25783\,
            I => \frame_decoder_CH4data_2\
        );

    \I__5843\ : CascadeMux
    port map (
            O => \N__25780\,
            I => \N__25777\
        );

    \I__5842\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25774\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__25774\,
            I => \frame_decoder_OFF4data_2\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__25771\,
            I => \N__25768\
        );

    \I__5839\ : InMux
    port map (
            O => \N__25768\,
            I => \N__25762\
        );

    \I__5838\ : InMux
    port map (
            O => \N__25767\,
            I => \N__25762\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__25762\,
            I => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\
        );

    \I__5836\ : InMux
    port map (
            O => \N__25759\,
            I => \scaler_4.un3_source_data_0_cry_1\
        );

    \I__5835\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25753\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__25753\,
            I => \frame_decoder_CH4data_3\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__25750\,
            I => \N__25747\
        );

    \I__5832\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25741\
        );

    \I__5831\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25741\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__25741\,
            I => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\
        );

    \I__5829\ : InMux
    port map (
            O => \N__25738\,
            I => \scaler_4.un3_source_data_0_cry_2\
        );

    \I__5828\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25732\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__25732\,
            I => \frame_decoder_CH4data_4\
        );

    \I__5826\ : CascadeMux
    port map (
            O => \N__25729\,
            I => \N__25726\
        );

    \I__5825\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25723\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__25723\,
            I => \N__25720\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__25720\,
            I => \frame_decoder_OFF4data_4\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__25717\,
            I => \N__25714\
        );

    \I__5821\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25708\
        );

    \I__5820\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25708\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__25708\,
            I => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\
        );

    \I__5818\ : InMux
    port map (
            O => \N__25705\,
            I => \scaler_4.un3_source_data_0_cry_3\
        );

    \I__5817\ : InMux
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__25699\,
            I => \frame_decoder_CH4data_5\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__25696\,
            I => \N__25693\
        );

    \I__5814\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25690\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__25690\,
            I => \frame_decoder_OFF4data_5\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__5811\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25678\
        );

    \I__5810\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25678\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__25678\,
            I => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\
        );

    \I__5808\ : InMux
    port map (
            O => \N__25675\,
            I => \scaler_4.un3_source_data_0_cry_4\
        );

    \I__5807\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25669\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25666\
        );

    \I__5805\ : Odrv4
    port map (
            O => \N__25666\,
            I => \frame_decoder_CH4data_6\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__25663\,
            I => \N__25660\
        );

    \I__5803\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25654\
        );

    \I__5802\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25654\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__25654\,
            I => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\
        );

    \I__5800\ : InMux
    port map (
            O => \N__25651\,
            I => \scaler_4.un3_source_data_0_cry_5\
        );

    \I__5799\ : InMux
    port map (
            O => \N__25648\,
            I => \N__25645\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__25645\,
            I => \scaler_4.un3_source_data_0_axb_7\
        );

    \I__5797\ : CascadeMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__5796\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25633\
        );

    \I__5795\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25633\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__25633\,
            I => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\
        );

    \I__5793\ : InMux
    port map (
            O => \N__25630\,
            I => \scaler_4.un3_source_data_0_cry_6\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__25627\,
            I => \N__25624\
        );

    \I__5791\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25621\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__25621\,
            I => \N__25618\
        );

    \I__5789\ : Span4Mux_v
    port map (
            O => \N__25618\,
            I => \N__25613\
        );

    \I__5788\ : CascadeMux
    port map (
            O => \N__25617\,
            I => \N__25609\
        );

    \I__5787\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25606\
        );

    \I__5786\ : Span4Mux_h
    port map (
            O => \N__25613\,
            I => \N__25603\
        );

    \I__5785\ : InMux
    port map (
            O => \N__25612\,
            I => \N__25598\
        );

    \I__5784\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25598\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__25606\,
            I => \N__25595\
        );

    \I__5782\ : Odrv4
    port map (
            O => \N__25603\,
            I => \Commands_frame_decoder.state_1Z0Z_6\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__25598\,
            I => \Commands_frame_decoder.state_1Z0Z_6\
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__25595\,
            I => \Commands_frame_decoder.state_1Z0Z_6\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__25588\,
            I => \N__25584\
        );

    \I__5778\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25579\
        );

    \I__5777\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25575\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__25583\,
            I => \N__25572\
        );

    \I__5775\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25568\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__25579\,
            I => \N__25563\
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__25578\,
            I => \N__25560\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__25575\,
            I => \N__25557\
        );

    \I__5771\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25552\
        );

    \I__5770\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25552\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__25568\,
            I => \N__25549\
        );

    \I__5768\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25544\
        );

    \I__5767\ : InMux
    port map (
            O => \N__25566\,
            I => \N__25544\
        );

    \I__5766\ : Span4Mux_h
    port map (
            O => \N__25563\,
            I => \N__25541\
        );

    \I__5765\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25538\
        );

    \I__5764\ : Odrv12
    port map (
            O => \N__25557\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__25552\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__25549\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__25544\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__25541\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__25538\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__5758\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25519\
        );

    \I__5757\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25516\
        );

    \I__5756\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25513\
        );

    \I__5755\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25510\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__25519\,
            I => \N__25507\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__25516\,
            I => \N__25502\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__25513\,
            I => \N__25502\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__25510\,
            I => \N__25499\
        );

    \I__5750\ : Span4Mux_v
    port map (
            O => \N__25507\,
            I => \N__25494\
        );

    \I__5749\ : Span4Mux_v
    port map (
            O => \N__25502\,
            I => \N__25494\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__25499\,
            I => \uart_drone.N_152\
        );

    \I__5747\ : Odrv4
    port map (
            O => \N__25494\,
            I => \uart_drone.N_152\
        );

    \I__5746\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__5745\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25483\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__25483\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__5743\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25476\
        );

    \I__5742\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25473\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__25476\,
            I => \Commands_frame_decoder.state_1Z0Z_7\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__25473\,
            I => \Commands_frame_decoder.state_1Z0Z_7\
        );

    \I__5739\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25465\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__25465\,
            I => \N__25462\
        );

    \I__5737\ : Span4Mux_h
    port map (
            O => \N__25462\,
            I => \N__25458\
        );

    \I__5736\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25455\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__25458\,
            I => \N__25450\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__25455\,
            I => \N__25450\
        );

    \I__5733\ : Span4Mux_v
    port map (
            O => \N__25450\,
            I => \N__25447\
        );

    \I__5732\ : Odrv4
    port map (
            O => \N__25447\,
            I => scaler_4_data_7
        );

    \I__5731\ : InMux
    port map (
            O => \N__25444\,
            I => \scaler_4.un2_source_data_0_cry_2\
        );

    \I__5730\ : InMux
    port map (
            O => \N__25441\,
            I => \N__25438\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__25438\,
            I => \N__25434\
        );

    \I__5728\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25431\
        );

    \I__5727\ : Span4Mux_v
    port map (
            O => \N__25434\,
            I => \N__25426\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25426\
        );

    \I__5725\ : Span4Mux_v
    port map (
            O => \N__25426\,
            I => \N__25423\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__25423\,
            I => scaler_4_data_8
        );

    \I__5723\ : InMux
    port map (
            O => \N__25420\,
            I => \scaler_4.un2_source_data_0_cry_3\
        );

    \I__5722\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25414\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__25414\,
            I => \N__25410\
        );

    \I__5720\ : InMux
    port map (
            O => \N__25413\,
            I => \N__25407\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__25410\,
            I => \N__25402\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__25407\,
            I => \N__25402\
        );

    \I__5717\ : Span4Mux_v
    port map (
            O => \N__25402\,
            I => \N__25399\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__25399\,
            I => scaler_4_data_9
        );

    \I__5715\ : InMux
    port map (
            O => \N__25396\,
            I => \scaler_4.un2_source_data_0_cry_4\
        );

    \I__5714\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25390\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25386\
        );

    \I__5712\ : InMux
    port map (
            O => \N__25389\,
            I => \N__25383\
        );

    \I__5711\ : Span4Mux_v
    port map (
            O => \N__25386\,
            I => \N__25378\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__25383\,
            I => \N__25378\
        );

    \I__5709\ : Span4Mux_v
    port map (
            O => \N__25378\,
            I => \N__25375\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__25375\,
            I => scaler_4_data_10
        );

    \I__5707\ : InMux
    port map (
            O => \N__25372\,
            I => \scaler_4.un2_source_data_0_cry_5\
        );

    \I__5706\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25366\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__25366\,
            I => \N__25362\
        );

    \I__5704\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25359\
        );

    \I__5703\ : Span4Mux_v
    port map (
            O => \N__25362\,
            I => \N__25354\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__25359\,
            I => \N__25354\
        );

    \I__5701\ : Span4Mux_v
    port map (
            O => \N__25354\,
            I => \N__25351\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__25351\,
            I => scaler_4_data_11
        );

    \I__5699\ : InMux
    port map (
            O => \N__25348\,
            I => \scaler_4.un2_source_data_0_cry_6\
        );

    \I__5698\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25342\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25338\
        );

    \I__5696\ : InMux
    port map (
            O => \N__25341\,
            I => \N__25335\
        );

    \I__5695\ : Span4Mux_v
    port map (
            O => \N__25338\,
            I => \N__25330\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__25335\,
            I => \N__25330\
        );

    \I__5693\ : Span4Mux_v
    port map (
            O => \N__25330\,
            I => \N__25327\
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__25327\,
            I => scaler_4_data_12
        );

    \I__5691\ : InMux
    port map (
            O => \N__25324\,
            I => \scaler_4.un2_source_data_0_cry_7\
        );

    \I__5690\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25318\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__25318\,
            I => \N__25315\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__25315\,
            I => \N__25311\
        );

    \I__5687\ : InMux
    port map (
            O => \N__25314\,
            I => \N__25308\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__25311\,
            I => \N__25303\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__25308\,
            I => \N__25303\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__25303\,
            I => \N__25300\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__25300\,
            I => scaler_4_data_13
        );

    \I__5682\ : InMux
    port map (
            O => \N__25297\,
            I => \bfn_10_16_0_\
        );

    \I__5681\ : InMux
    port map (
            O => \N__25294\,
            I => \scaler_4.un2_source_data_0_cry_9\
        );

    \I__5680\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25288\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__25288\,
            I => \N__25285\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__25285\,
            I => \N__25282\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__25282\,
            I => \N__25279\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__25279\,
            I => scaler_4_data_14
        );

    \I__5675\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25272\
        );

    \I__5674\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25268\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__25272\,
            I => \N__25265\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__25271\,
            I => \N__25262\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__25268\,
            I => \N__25258\
        );

    \I__5670\ : Span4Mux_h
    port map (
            O => \N__25265\,
            I => \N__25255\
        );

    \I__5669\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25250\
        );

    \I__5668\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25250\
        );

    \I__5667\ : Odrv4
    port map (
            O => \N__25258\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__25255\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__25250\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__5664\ : InMux
    port map (
            O => \N__25243\,
            I => \N__25238\
        );

    \I__5663\ : InMux
    port map (
            O => \N__25242\,
            I => \N__25235\
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__25241\,
            I => \N__25231\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__25238\,
            I => \N__25228\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__25235\,
            I => \N__25225\
        );

    \I__5659\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25222\
        );

    \I__5658\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25219\
        );

    \I__5657\ : Odrv12
    port map (
            O => \N__25228\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__25225\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__25222\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__25219\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5653\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25205\
        );

    \I__5652\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25202\
        );

    \I__5651\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25199\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__25205\,
            I => \N__25195\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__25202\,
            I => \N__25192\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__25199\,
            I => \N__25189\
        );

    \I__5647\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25186\
        );

    \I__5646\ : Span4Mux_v
    port map (
            O => \N__25195\,
            I => \N__25183\
        );

    \I__5645\ : Span12Mux_h
    port map (
            O => \N__25192\,
            I => \N__25180\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__25189\,
            I => \N__25177\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__25186\,
            I => \N__25174\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__25183\,
            I => \frame_decoder_CH2data_0\
        );

    \I__5641\ : Odrv12
    port map (
            O => \N__25180\,
            I => \frame_decoder_CH2data_0\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__25177\,
            I => \frame_decoder_CH2data_0\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__25174\,
            I => \frame_decoder_CH2data_0\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__25165\,
            I => \N__25162\
        );

    \I__5637\ : InMux
    port map (
            O => \N__25162\,
            I => \N__25159\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__25159\,
            I => \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\
        );

    \I__5635\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25150\
        );

    \I__5634\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25150\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__25150\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__25147\,
            I => \N__25144\
        );

    \I__5631\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25141\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__25141\,
            I => \N__25138\
        );

    \I__5629\ : Span4Mux_h
    port map (
            O => \N__25138\,
            I => \N__25135\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__25135\,
            I => \scaler_4.un2_source_data_0_cry_1_c_RNO_1\
        );

    \I__5627\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25128\
        );

    \I__5626\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25125\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__25128\,
            I => \N__25122\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__25125\,
            I => \N__25119\
        );

    \I__5623\ : Span12Mux_v
    port map (
            O => \N__25122\,
            I => \N__25116\
        );

    \I__5622\ : Span4Mux_v
    port map (
            O => \N__25119\,
            I => \N__25113\
        );

    \I__5621\ : Odrv12
    port map (
            O => \N__25116\,
            I => scaler_4_data_6
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__25113\,
            I => scaler_4_data_6
        );

    \I__5619\ : InMux
    port map (
            O => \N__25108\,
            I => \scaler_4.un2_source_data_0_cry_1\
        );

    \I__5618\ : InMux
    port map (
            O => \N__25105\,
            I => \ppm_encoder_1.un1_elevator_cry_12\
        );

    \I__5617\ : InMux
    port map (
            O => \N__25102\,
            I => \bfn_9_20_0_\
        );

    \I__5616\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25095\
        );

    \I__5615\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25092\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25089\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__25092\,
            I => \N__25084\
        );

    \I__5612\ : Span4Mux_h
    port map (
            O => \N__25089\,
            I => \N__25084\
        );

    \I__5611\ : Span4Mux_v
    port map (
            O => \N__25084\,
            I => \N__25081\
        );

    \I__5610\ : Odrv4
    port map (
            O => \N__25081\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__5609\ : CEMux
    port map (
            O => \N__25078\,
            I => \N__25073\
        );

    \I__5608\ : CEMux
    port map (
            O => \N__25077\,
            I => \N__25070\
        );

    \I__5607\ : CEMux
    port map (
            O => \N__25076\,
            I => \N__25067\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__25073\,
            I => \N__25062\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__25070\,
            I => \N__25057\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25057\
        );

    \I__5603\ : CEMux
    port map (
            O => \N__25066\,
            I => \N__25054\
        );

    \I__5602\ : CEMux
    port map (
            O => \N__25065\,
            I => \N__25051\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__25062\,
            I => \N__25043\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__25057\,
            I => \N__25043\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__25054\,
            I => \N__25043\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__25051\,
            I => \N__25039\
        );

    \I__5597\ : CEMux
    port map (
            O => \N__25050\,
            I => \N__25036\
        );

    \I__5596\ : Sp12to4
    port map (
            O => \N__25043\,
            I => \N__25033\
        );

    \I__5595\ : CEMux
    port map (
            O => \N__25042\,
            I => \N__25030\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__25039\,
            I => \N__25025\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__25036\,
            I => \N__25025\
        );

    \I__5592\ : Span12Mux_s4_h
    port map (
            O => \N__25033\,
            I => \N__25020\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__25020\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__25025\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__5589\ : Odrv12
    port map (
            O => \N__25020\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__5588\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25012\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__25012\,
            I => \N__25009\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__25009\,
            I => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\
        );

    \I__5585\ : InMux
    port map (
            O => \N__25006\,
            I => \N__25002\
        );

    \I__5584\ : InMux
    port map (
            O => \N__25005\,
            I => \N__24998\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__25002\,
            I => \N__24995\
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__25001\,
            I => \N__24992\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__24998\,
            I => \N__24987\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__24995\,
            I => \N__24987\
        );

    \I__5579\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24984\
        );

    \I__5578\ : Span4Mux_h
    port map (
            O => \N__24987\,
            I => \N__24981\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__24984\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__24981\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__5575\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24973\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__24973\,
            I => \N__24970\
        );

    \I__5573\ : Odrv12
    port map (
            O => \N__24970\,
            I => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__24967\,
            I => \N__24956\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__24966\,
            I => \N__24951\
        );

    \I__5570\ : CascadeMux
    port map (
            O => \N__24965\,
            I => \N__24944\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__24964\,
            I => \N__24941\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__24963\,
            I => \N__24935\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__24962\,
            I => \N__24932\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__24961\,
            I => \N__24929\
        );

    \I__5565\ : CascadeMux
    port map (
            O => \N__24960\,
            I => \N__24926\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__24959\,
            I => \N__24923\
        );

    \I__5563\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24920\
        );

    \I__5562\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24917\
        );

    \I__5561\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24914\
        );

    \I__5560\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24904\
        );

    \I__5559\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24891\
        );

    \I__5558\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24891\
        );

    \I__5557\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24891\
        );

    \I__5556\ : InMux
    port map (
            O => \N__24947\,
            I => \N__24891\
        );

    \I__5555\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24891\
        );

    \I__5554\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24891\
        );

    \I__5553\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24880\
        );

    \I__5552\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24880\
        );

    \I__5551\ : InMux
    port map (
            O => \N__24938\,
            I => \N__24880\
        );

    \I__5550\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24880\
        );

    \I__5549\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24880\
        );

    \I__5548\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24877\
        );

    \I__5547\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24874\
        );

    \I__5546\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24871\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__24920\,
            I => \N__24857\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__24917\,
            I => \N__24857\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__24914\,
            I => \N__24857\
        );

    \I__5542\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24854\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__24912\,
            I => \N__24850\
        );

    \I__5540\ : CascadeMux
    port map (
            O => \N__24911\,
            I => \N__24847\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__24910\,
            I => \N__24844\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__24909\,
            I => \N__24837\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__24908\,
            I => \N__24834\
        );

    \I__5536\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24831\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24828\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__24891\,
            I => \N__24823\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__24880\,
            I => \N__24823\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24820\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__24874\,
            I => \N__24815\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__24871\,
            I => \N__24815\
        );

    \I__5529\ : CascadeMux
    port map (
            O => \N__24870\,
            I => \N__24812\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__24869\,
            I => \N__24809\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__24868\,
            I => \N__24806\
        );

    \I__5526\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24799\
        );

    \I__5525\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24799\
        );

    \I__5524\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24799\
        );

    \I__5523\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24794\
        );

    \I__5522\ : Span4Mux_v
    port map (
            O => \N__24857\,
            I => \N__24791\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__24854\,
            I => \N__24788\
        );

    \I__5520\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24779\
        );

    \I__5519\ : InMux
    port map (
            O => \N__24850\,
            I => \N__24779\
        );

    \I__5518\ : InMux
    port map (
            O => \N__24847\,
            I => \N__24779\
        );

    \I__5517\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24779\
        );

    \I__5516\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24770\
        );

    \I__5515\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24770\
        );

    \I__5514\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24770\
        );

    \I__5513\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24770\
        );

    \I__5512\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24767\
        );

    \I__5511\ : InMux
    port map (
            O => \N__24834\,
            I => \N__24764\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__24831\,
            I => \N__24761\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__24828\,
            I => \N__24754\
        );

    \I__5508\ : Span4Mux_v
    port map (
            O => \N__24823\,
            I => \N__24754\
        );

    \I__5507\ : Span4Mux_h
    port map (
            O => \N__24820\,
            I => \N__24754\
        );

    \I__5506\ : Span4Mux_v
    port map (
            O => \N__24815\,
            I => \N__24751\
        );

    \I__5505\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24744\
        );

    \I__5504\ : InMux
    port map (
            O => \N__24809\,
            I => \N__24744\
        );

    \I__5503\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24744\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__24799\,
            I => \N__24741\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__24798\,
            I => \N__24738\
        );

    \I__5500\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24735\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__24794\,
            I => \N__24732\
        );

    \I__5498\ : Span4Mux_h
    port map (
            O => \N__24791\,
            I => \N__24727\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__24788\,
            I => \N__24727\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24714\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24714\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__24767\,
            I => \N__24714\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__24764\,
            I => \N__24714\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__24761\,
            I => \N__24714\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__24754\,
            I => \N__24714\
        );

    \I__5490\ : Span4Mux_h
    port map (
            O => \N__24751\,
            I => \N__24707\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__24744\,
            I => \N__24707\
        );

    \I__5488\ : Span4Mux_h
    port map (
            O => \N__24741\,
            I => \N__24707\
        );

    \I__5487\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24704\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__24735\,
            I => \N__24701\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__24732\,
            I => \N__24696\
        );

    \I__5484\ : Span4Mux_v
    port map (
            O => \N__24727\,
            I => \N__24696\
        );

    \I__5483\ : Span4Mux_v
    port map (
            O => \N__24714\,
            I => \N__24693\
        );

    \I__5482\ : Span4Mux_v
    port map (
            O => \N__24707\,
            I => \N__24690\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__24704\,
            I => \N__24685\
        );

    \I__5480\ : Span4Mux_v
    port map (
            O => \N__24701\,
            I => \N__24685\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__24696\,
            I => pid_altitude_dv
        );

    \I__5478\ : Odrv4
    port map (
            O => \N__24693\,
            I => pid_altitude_dv
        );

    \I__5477\ : Odrv4
    port map (
            O => \N__24690\,
            I => pid_altitude_dv
        );

    \I__5476\ : Odrv4
    port map (
            O => \N__24685\,
            I => pid_altitude_dv
        );

    \I__5475\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24671\
        );

    \I__5474\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24668\
        );

    \I__5473\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24665\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24660\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__24668\,
            I => \N__24660\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__24665\,
            I => \N__24655\
        );

    \I__5469\ : Span4Mux_h
    port map (
            O => \N__24660\,
            I => \N__24655\
        );

    \I__5468\ : Odrv4
    port map (
            O => \N__24655\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__5467\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24648\
        );

    \I__5466\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24645\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24642\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__24645\,
            I => \N__24639\
        );

    \I__5463\ : Odrv4
    port map (
            O => \N__24642\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__5462\ : Odrv12
    port map (
            O => \N__24639\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__5461\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24628\
        );

    \I__5460\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24628\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__24628\,
            I => \frame_decoder_CH4data_7\
        );

    \I__5458\ : CEMux
    port map (
            O => \N__24625\,
            I => \N__24621\
        );

    \I__5457\ : CEMux
    port map (
            O => \N__24624\,
            I => \N__24618\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__24621\,
            I => \N__24614\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__24618\,
            I => \N__24611\
        );

    \I__5454\ : CEMux
    port map (
            O => \N__24617\,
            I => \N__24608\
        );

    \I__5453\ : Span4Mux_h
    port map (
            O => \N__24614\,
            I => \N__24605\
        );

    \I__5452\ : Span4Mux_v
    port map (
            O => \N__24611\,
            I => \N__24600\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24600\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__24605\,
            I => \N__24597\
        );

    \I__5449\ : Sp12to4
    port map (
            O => \N__24600\,
            I => \N__24594\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__24597\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\
        );

    \I__5447\ : Odrv12
    port map (
            O => \N__24594\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\
        );

    \I__5446\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24586\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__24586\,
            I => \N__24583\
        );

    \I__5444\ : Span4Mux_v
    port map (
            O => \N__24583\,
            I => \N__24580\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__24580\,
            I => \N__24577\
        );

    \I__5442\ : Span4Mux_h
    port map (
            O => \N__24577\,
            I => \N__24574\
        );

    \I__5441\ : Odrv4
    port map (
            O => \N__24574\,
            I => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\
        );

    \I__5440\ : InMux
    port map (
            O => \N__24571\,
            I => \ppm_encoder_1.un1_elevator_cry_6\
        );

    \I__5439\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24565\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__5437\ : Span4Mux_v
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__24559\,
            I => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\
        );

    \I__5435\ : InMux
    port map (
            O => \N__24556\,
            I => \ppm_encoder_1.un1_elevator_cry_7\
        );

    \I__5434\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24550\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__24550\,
            I => \N__24547\
        );

    \I__5432\ : Span4Mux_v
    port map (
            O => \N__24547\,
            I => \N__24544\
        );

    \I__5431\ : Span4Mux_h
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__24541\,
            I => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\
        );

    \I__5429\ : InMux
    port map (
            O => \N__24538\,
            I => \ppm_encoder_1.un1_elevator_cry_8\
        );

    \I__5428\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24532\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__24532\,
            I => \N__24529\
        );

    \I__5426\ : Odrv4
    port map (
            O => \N__24529\,
            I => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\
        );

    \I__5425\ : InMux
    port map (
            O => \N__24526\,
            I => \ppm_encoder_1.un1_elevator_cry_9\
        );

    \I__5424\ : InMux
    port map (
            O => \N__24523\,
            I => \ppm_encoder_1.un1_elevator_cry_10\
        );

    \I__5423\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24517\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__5421\ : Odrv4
    port map (
            O => \N__24514\,
            I => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\
        );

    \I__5420\ : InMux
    port map (
            O => \N__24511\,
            I => \ppm_encoder_1.un1_elevator_cry_11\
        );

    \I__5419\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__24505\,
            I => \N__24502\
        );

    \I__5417\ : Span4Mux_h
    port map (
            O => \N__24502\,
            I => \N__24499\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__24499\,
            I => \N__24495\
        );

    \I__5415\ : CascadeMux
    port map (
            O => \N__24498\,
            I => \N__24492\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__24495\,
            I => \N__24489\
        );

    \I__5413\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24486\
        );

    \I__5412\ : Odrv4
    port map (
            O => \N__24489\,
            I => scaler_3_data_4
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__24486\,
            I => scaler_3_data_4
        );

    \I__5410\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__5408\ : Span4Mux_h
    port map (
            O => \N__24475\,
            I => \N__24472\
        );

    \I__5407\ : Span4Mux_h
    port map (
            O => \N__24472\,
            I => \N__24469\
        );

    \I__5406\ : Span4Mux_v
    port map (
            O => \N__24469\,
            I => \N__24465\
        );

    \I__5405\ : CascadeMux
    port map (
            O => \N__24468\,
            I => \N__24462\
        );

    \I__5404\ : Span4Mux_v
    port map (
            O => \N__24465\,
            I => \N__24459\
        );

    \I__5403\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24456\
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__24459\,
            I => scaler_4_data_4
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__24456\,
            I => scaler_4_data_4
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__24451\,
            I => \Commands_frame_decoder.N_282_0_cascade_\
        );

    \I__5399\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24444\
        );

    \I__5398\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24441\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24436\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__24441\,
            I => \N__24436\
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__24436\,
            I => \Commands_frame_decoder.state_1_ns_0_a4_0_0Z0Z_1\
        );

    \I__5394\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24430\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24427\
        );

    \I__5392\ : Span4Mux_h
    port map (
            O => \N__24427\,
            I => \N__24424\
        );

    \I__5391\ : Span4Mux_h
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__24421\,
            I => \Commands_frame_decoder.source_CH1data8lto7Z0Z_1\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__24418\,
            I => \Commands_frame_decoder.N_319_cascade_\
        );

    \I__5388\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24412\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__24412\,
            I => \Commands_frame_decoder.N_318\
        );

    \I__5386\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24406\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__24406\,
            I => \Commands_frame_decoder.N_282_0\
        );

    \I__5384\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__24400\,
            I => \Commands_frame_decoder.state_1_RNO_1Z0Z_0\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__24397\,
            I => \Commands_frame_decoder.state_1_ns_i_0_0_cascade_\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__24394\,
            I => \N__24390\
        );

    \I__5380\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24385\
        );

    \I__5379\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24385\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__24385\,
            I => \Commands_frame_decoder.state_1Z0Z_0\
        );

    \I__5377\ : InMux
    port map (
            O => \N__24382\,
            I => \N__24376\
        );

    \I__5376\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24376\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24373\
        );

    \I__5374\ : Span4Mux_h
    port map (
            O => \N__24373\,
            I => \N__24370\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__24370\,
            I => \Commands_frame_decoder.N_323\
        );

    \I__5372\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24364\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__24364\,
            I => \Commands_frame_decoder.state_1_ns_0_a4_0_2_1\
        );

    \I__5370\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24358\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24355\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__24355\,
            I => \N__24350\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__24354\,
            I => \N__24347\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__24353\,
            I => \N__24344\
        );

    \I__5365\ : Span4Mux_h
    port map (
            O => \N__24350\,
            I => \N__24340\
        );

    \I__5364\ : InMux
    port map (
            O => \N__24347\,
            I => \N__24333\
        );

    \I__5363\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24333\
        );

    \I__5362\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24333\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__24340\,
            I => \Commands_frame_decoder.state_1Z0Z_1\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__24333\,
            I => \Commands_frame_decoder.state_1Z0Z_1\
        );

    \I__5359\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24324\
        );

    \I__5358\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24321\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__24324\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__24321\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__24316\,
            I => \N__24313\
        );

    \I__5354\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24310\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__24310\,
            I => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\
        );

    \I__5352\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24303\
        );

    \I__5351\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24300\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__24303\,
            I => \N__24297\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24294\
        );

    \I__5348\ : Span12Mux_s9_h
    port map (
            O => \N__24297\,
            I => \N__24291\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__24294\,
            I => \N__24288\
        );

    \I__5346\ : Odrv12
    port map (
            O => \N__24291\,
            I => scaler_2_data_13
        );

    \I__5345\ : Odrv4
    port map (
            O => \N__24288\,
            I => scaler_2_data_13
        );

    \I__5344\ : InMux
    port map (
            O => \N__24283\,
            I => \bfn_9_14_0_\
        );

    \I__5343\ : InMux
    port map (
            O => \N__24280\,
            I => \scaler_2.un2_source_data_0_cry_9\
        );

    \I__5342\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24274\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__24274\,
            I => \N__24271\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__24271\,
            I => \N__24268\
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__24268\,
            I => scaler_2_data_14
        );

    \I__5338\ : InMux
    port map (
            O => \N__24265\,
            I => \N__24262\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__24262\,
            I => \N__24259\
        );

    \I__5336\ : Sp12to4
    port map (
            O => \N__24259\,
            I => \N__24256\
        );

    \I__5335\ : Span12Mux_v
    port map (
            O => \N__24256\,
            I => \N__24253\
        );

    \I__5334\ : Odrv12
    port map (
            O => \N__24253\,
            I => scaler_2_data_5
        );

    \I__5333\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24247\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__24247\,
            I => \N__24244\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__24244\,
            I => \N__24241\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__24241\,
            I => \N__24238\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__24238\,
            I => \N__24235\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__24235\,
            I => scaler_3_data_5
        );

    \I__5327\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24229\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24226\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__24226\,
            I => \N__24223\
        );

    \I__5324\ : Span4Mux_v
    port map (
            O => \N__24223\,
            I => \N__24220\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__24220\,
            I => \N__24217\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__24217\,
            I => scaler_4_data_5
        );

    \I__5321\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24211\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__24211\,
            I => \uart_drone.data_Auxce_0_0_0\
        );

    \I__5319\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24205\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__24205\,
            I => \N__24202\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__24202\,
            I => \N__24199\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__24199\,
            I => \N__24195\
        );

    \I__5315\ : CascadeMux
    port map (
            O => \N__24198\,
            I => \N__24192\
        );

    \I__5314\ : Span4Mux_h
    port map (
            O => \N__24195\,
            I => \N__24189\
        );

    \I__5313\ : InMux
    port map (
            O => \N__24192\,
            I => \N__24186\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__24189\,
            I => scaler_2_data_4
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__24186\,
            I => scaler_2_data_4
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__24181\,
            I => \N__24178\
        );

    \I__5309\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24175\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__24175\,
            I => \frame_decoder_OFF2data_2\
        );

    \I__5307\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24169\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__24169\,
            I => \N__24166\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__24166\,
            I => \N__24163\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__24163\,
            I => \N__24159\
        );

    \I__5303\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24156\
        );

    \I__5302\ : Span4Mux_h
    port map (
            O => \N__24159\,
            I => \N__24151\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__24156\,
            I => \N__24151\
        );

    \I__5300\ : Sp12to4
    port map (
            O => \N__24151\,
            I => \N__24148\
        );

    \I__5299\ : Odrv12
    port map (
            O => \N__24148\,
            I => scaler_2_data_6
        );

    \I__5298\ : InMux
    port map (
            O => \N__24145\,
            I => \scaler_2.un2_source_data_0_cry_1\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__24142\,
            I => \N__24139\
        );

    \I__5296\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24133\
        );

    \I__5295\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24133\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__24133\,
            I => \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\
        );

    \I__5293\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24126\
        );

    \I__5292\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24123\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__24126\,
            I => \N__24120\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__24123\,
            I => \N__24117\
        );

    \I__5289\ : Span12Mux_s9_h
    port map (
            O => \N__24120\,
            I => \N__24114\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__24117\,
            I => \N__24111\
        );

    \I__5287\ : Odrv12
    port map (
            O => \N__24114\,
            I => scaler_2_data_7
        );

    \I__5286\ : Odrv4
    port map (
            O => \N__24111\,
            I => scaler_2_data_7
        );

    \I__5285\ : InMux
    port map (
            O => \N__24106\,
            I => \scaler_2.un2_source_data_0_cry_2\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__24103\,
            I => \N__24100\
        );

    \I__5283\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24094\
        );

    \I__5282\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24094\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__24094\,
            I => \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\
        );

    \I__5280\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24088\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__24088\,
            I => \N__24085\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__24085\,
            I => \N__24081\
        );

    \I__5277\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24078\
        );

    \I__5276\ : Span4Mux_h
    port map (
            O => \N__24081\,
            I => \N__24073\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24073\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__24073\,
            I => \N__24070\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__24070\,
            I => scaler_2_data_8
        );

    \I__5272\ : InMux
    port map (
            O => \N__24067\,
            I => \scaler_2.un2_source_data_0_cry_3\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__24064\,
            I => \N__24061\
        );

    \I__5270\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24055\
        );

    \I__5269\ : InMux
    port map (
            O => \N__24060\,
            I => \N__24055\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__24055\,
            I => \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\
        );

    \I__5267\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24049\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24045\
        );

    \I__5265\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24042\
        );

    \I__5264\ : Span4Mux_v
    port map (
            O => \N__24045\,
            I => \N__24039\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__24042\,
            I => \N__24036\
        );

    \I__5262\ : Span4Mux_v
    port map (
            O => \N__24039\,
            I => \N__24033\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__24036\,
            I => \N__24030\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__24033\,
            I => scaler_2_data_9
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__24030\,
            I => scaler_2_data_9
        );

    \I__5258\ : InMux
    port map (
            O => \N__24025\,
            I => \scaler_2.un2_source_data_0_cry_4\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__24022\,
            I => \N__24019\
        );

    \I__5256\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24013\
        );

    \I__5255\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24013\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__24013\,
            I => \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\
        );

    \I__5253\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24007\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__24007\,
            I => \N__24004\
        );

    \I__5251\ : Span4Mux_h
    port map (
            O => \N__24004\,
            I => \N__24000\
        );

    \I__5250\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23997\
        );

    \I__5249\ : Span4Mux_v
    port map (
            O => \N__24000\,
            I => \N__23994\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__23997\,
            I => \N__23991\
        );

    \I__5247\ : Span4Mux_v
    port map (
            O => \N__23994\,
            I => \N__23988\
        );

    \I__5246\ : Span4Mux_v
    port map (
            O => \N__23991\,
            I => \N__23985\
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__23988\,
            I => scaler_2_data_10
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__23985\,
            I => scaler_2_data_10
        );

    \I__5243\ : InMux
    port map (
            O => \N__23980\,
            I => \scaler_2.un2_source_data_0_cry_5\
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__23977\,
            I => \N__23974\
        );

    \I__5241\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23968\
        );

    \I__5240\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23968\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__23968\,
            I => \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\
        );

    \I__5238\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23962\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__23962\,
            I => \N__23959\
        );

    \I__5236\ : Span4Mux_v
    port map (
            O => \N__23959\,
            I => \N__23955\
        );

    \I__5235\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23952\
        );

    \I__5234\ : Sp12to4
    port map (
            O => \N__23955\,
            I => \N__23947\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__23952\,
            I => \N__23947\
        );

    \I__5232\ : Span12Mux_s9_h
    port map (
            O => \N__23947\,
            I => \N__23944\
        );

    \I__5231\ : Odrv12
    port map (
            O => \N__23944\,
            I => scaler_2_data_11
        );

    \I__5230\ : InMux
    port map (
            O => \N__23941\,
            I => \scaler_2.un2_source_data_0_cry_6\
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__23938\,
            I => \N__23935\
        );

    \I__5228\ : InMux
    port map (
            O => \N__23935\,
            I => \N__23929\
        );

    \I__5227\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23929\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__23929\,
            I => \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\
        );

    \I__5225\ : InMux
    port map (
            O => \N__23926\,
            I => \N__23923\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__23923\,
            I => \N__23920\
        );

    \I__5223\ : Span4Mux_v
    port map (
            O => \N__23920\,
            I => \N__23916\
        );

    \I__5222\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23913\
        );

    \I__5221\ : Sp12to4
    port map (
            O => \N__23916\,
            I => \N__23910\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__23913\,
            I => \N__23907\
        );

    \I__5219\ : Span12Mux_s9_h
    port map (
            O => \N__23910\,
            I => \N__23904\
        );

    \I__5218\ : Span4Mux_v
    port map (
            O => \N__23907\,
            I => \N__23901\
        );

    \I__5217\ : Odrv12
    port map (
            O => \N__23904\,
            I => scaler_2_data_12
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__23901\,
            I => scaler_2_data_12
        );

    \I__5215\ : InMux
    port map (
            O => \N__23896\,
            I => \scaler_2.un2_source_data_0_cry_7\
        );

    \I__5214\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__5212\ : Span4Mux_s3_v
    port map (
            O => \N__23887\,
            I => \N__23882\
        );

    \I__5211\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23877\
        );

    \I__5210\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23877\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__23882\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__23877\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__23872\,
            I => \N__23867\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__23871\,
            I => \N__23864\
        );

    \I__5205\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23857\
        );

    \I__5204\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23857\
        );

    \I__5203\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23857\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__23857\,
            I => \N__23854\
        );

    \I__5201\ : Span4Mux_s3_v
    port map (
            O => \N__23854\,
            I => \N__23851\
        );

    \I__5200\ : Span4Mux_v
    port map (
            O => \N__23851\,
            I => \N__23846\
        );

    \I__5199\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23843\
        );

    \I__5198\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23840\
        );

    \I__5197\ : Sp12to4
    port map (
            O => \N__23846\,
            I => \N__23835\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__23843\,
            I => \N__23835\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__23840\,
            I => \N__23832\
        );

    \I__5194\ : Odrv12
    port map (
            O => \N__23835\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_158_d\
        );

    \I__5193\ : Odrv12
    port map (
            O => \N__23832\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_158_d\
        );

    \I__5192\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23814\
        );

    \I__5191\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23814\
        );

    \I__5190\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23814\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__23824\,
            I => \N__23804\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__23823\,
            I => \N__23801\
        );

    \I__5187\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23789\
        );

    \I__5186\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23789\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__23814\,
            I => \N__23781\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__23813\,
            I => \N__23777\
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__23812\,
            I => \N__23774\
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__23811\,
            I => \N__23768\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__23810\,
            I => \N__23764\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__23809\,
            I => \N__23757\
        );

    \I__5179\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23750\
        );

    \I__5178\ : CascadeMux
    port map (
            O => \N__23807\,
            I => \N__23745\
        );

    \I__5177\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23737\
        );

    \I__5176\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23737\
        );

    \I__5175\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23737\
        );

    \I__5174\ : CascadeMux
    port map (
            O => \N__23799\,
            I => \N__23734\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__23798\,
            I => \N__23728\
        );

    \I__5172\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23725\
        );

    \I__5171\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23717\
        );

    \I__5170\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23717\
        );

    \I__5169\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23717\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__23789\,
            I => \N__23714\
        );

    \I__5167\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23703\
        );

    \I__5166\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23703\
        );

    \I__5165\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23703\
        );

    \I__5164\ : InMux
    port map (
            O => \N__23785\,
            I => \N__23703\
        );

    \I__5163\ : InMux
    port map (
            O => \N__23784\,
            I => \N__23703\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__23781\,
            I => \N__23699\
        );

    \I__5161\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23696\
        );

    \I__5160\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23687\
        );

    \I__5159\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23687\
        );

    \I__5158\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23687\
        );

    \I__5157\ : InMux
    port map (
            O => \N__23772\,
            I => \N__23687\
        );

    \I__5156\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23676\
        );

    \I__5155\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23676\
        );

    \I__5154\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23676\
        );

    \I__5153\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23676\
        );

    \I__5152\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23676\
        );

    \I__5151\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23669\
        );

    \I__5150\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23669\
        );

    \I__5149\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23669\
        );

    \I__5148\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23658\
        );

    \I__5147\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23658\
        );

    \I__5146\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23658\
        );

    \I__5145\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23658\
        );

    \I__5144\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23658\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__23750\,
            I => \N__23647\
        );

    \I__5142\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23638\
        );

    \I__5141\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23638\
        );

    \I__5140\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23638\
        );

    \I__5139\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23638\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__23737\,
            I => \N__23635\
        );

    \I__5137\ : InMux
    port map (
            O => \N__23734\,
            I => \N__23630\
        );

    \I__5136\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23630\
        );

    \I__5135\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23624\
        );

    \I__5134\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23624\
        );

    \I__5133\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23621\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__23725\,
            I => \N__23618\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__23724\,
            I => \N__23614\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__23717\,
            I => \N__23605\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__23714\,
            I => \N__23605\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__23703\,
            I => \N__23605\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__23702\,
            I => \N__23602\
        );

    \I__5126\ : Span4Mux_h
    port map (
            O => \N__23699\,
            I => \N__23588\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__23696\,
            I => \N__23588\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__23687\,
            I => \N__23588\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__23676\,
            I => \N__23588\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__23669\,
            I => \N__23588\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__23658\,
            I => \N__23588\
        );

    \I__5120\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23575\
        );

    \I__5119\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23575\
        );

    \I__5118\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23575\
        );

    \I__5117\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23575\
        );

    \I__5116\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23575\
        );

    \I__5115\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23575\
        );

    \I__5114\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23570\
        );

    \I__5113\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23570\
        );

    \I__5112\ : Span4Mux_v
    port map (
            O => \N__23647\,
            I => \N__23561\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23561\
        );

    \I__5110\ : Span4Mux_v
    port map (
            O => \N__23635\,
            I => \N__23561\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23561\
        );

    \I__5108\ : CascadeMux
    port map (
            O => \N__23629\,
            I => \N__23553\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__23624\,
            I => \N__23549\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__23621\,
            I => \N__23544\
        );

    \I__5105\ : Span12Mux_h
    port map (
            O => \N__23618\,
            I => \N__23544\
        );

    \I__5104\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23535\
        );

    \I__5103\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23535\
        );

    \I__5102\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23535\
        );

    \I__5101\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23535\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__23605\,
            I => \N__23532\
        );

    \I__5099\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23527\
        );

    \I__5098\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23527\
        );

    \I__5097\ : Span4Mux_v
    port map (
            O => \N__23588\,
            I => \N__23518\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__23575\,
            I => \N__23518\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23518\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__23561\,
            I => \N__23518\
        );

    \I__5093\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23509\
        );

    \I__5092\ : InMux
    port map (
            O => \N__23559\,
            I => \N__23509\
        );

    \I__5091\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23509\
        );

    \I__5090\ : InMux
    port map (
            O => \N__23557\,
            I => \N__23509\
        );

    \I__5089\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23502\
        );

    \I__5088\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23502\
        );

    \I__5087\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23502\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__23549\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5085\ : Odrv12
    port map (
            O => \N__23544\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__23535\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__23532\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__23527\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__23518\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__23509\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__23502\,
            I => \ppm_encoder_1.PPM_STATE_58_d\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__23485\,
            I => \N__23481\
        );

    \I__5077\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23478\
        );

    \I__5076\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23475\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__23478\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__23475\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__5073\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23465\
        );

    \I__5072\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23462\
        );

    \I__5071\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23459\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__23465\,
            I => \N__23456\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__23462\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__23459\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5067\ : Odrv4
    port map (
            O => \N__23456\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5066\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23444\
        );

    \I__5065\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23441\
        );

    \I__5064\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23438\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23435\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__23441\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__23438\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__23435\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5059\ : CascadeMux
    port map (
            O => \N__23428\,
            I => \N__23423\
        );

    \I__5058\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23420\
        );

    \I__5057\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23417\
        );

    \I__5056\ : InMux
    port map (
            O => \N__23423\,
            I => \N__23414\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__23420\,
            I => \N__23411\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__23417\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__23414\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__23411\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5051\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23399\
        );

    \I__5050\ : InMux
    port map (
            O => \N__23403\,
            I => \N__23396\
        );

    \I__5049\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23393\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__23399\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__23396\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__23393\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5045\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23382\
        );

    \I__5044\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23379\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__23382\,
            I => \N__23376\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__23379\,
            I => \N__23373\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__23376\,
            I => \N__23370\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__23373\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__23370\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\
        );

    \I__5038\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23362\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__23362\,
            I => uart_input_pc_c
        );

    \I__5036\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23356\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__23356\,
            I => \uart_pc_sync.aux_0__0__0_0\
        );

    \I__5034\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23350\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__23350\,
            I => \N__23347\
        );

    \I__5032\ : Odrv4
    port map (
            O => \N__23347\,
            I => \uart_pc_sync.aux_1__0__0_0\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__23344\,
            I => \N__23341\
        );

    \I__5030\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23335\
        );

    \I__5029\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23335\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__23335\,
            I => \frame_decoder_OFF2data_7\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__23332\,
            I => \N__23329\
        );

    \I__5026\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23326\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__23326\,
            I => \frame_decoder_OFF2data_1\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__23323\,
            I => \N__23320\
        );

    \I__5023\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23317\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__23317\,
            I => \frame_decoder_OFF2data_4\
        );

    \I__5021\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23309\
        );

    \I__5020\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23306\
        );

    \I__5019\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23303\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__23309\,
            I => \N__23300\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__23306\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__23303\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__23300\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5014\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23290\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__23290\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\
        );

    \I__5012\ : CascadeMux
    port map (
            O => \N__23287\,
            I => \N__23283\
        );

    \I__5011\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23279\
        );

    \I__5010\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23276\
        );

    \I__5009\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23273\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__23279\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__23276\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__23273\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__23266\,
            I => \N__23263\
        );

    \I__5004\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23260\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__23260\,
            I => \N__23257\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__23257\,
            I => \ppm_encoder_1.pulses2countZ0Z_7\
        );

    \I__5001\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23249\
        );

    \I__5000\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23246\
        );

    \I__4999\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23243\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__23249\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__23246\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__23243\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__4995\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23233\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__23233\,
            I => \N__23230\
        );

    \I__4993\ : Odrv12
    port map (
            O => \N__23230\,
            I => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\
        );

    \I__4992\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23224\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__23224\,
            I => \N__23221\
        );

    \I__4990\ : Span4Mux_v
    port map (
            O => \N__23221\,
            I => \N__23218\
        );

    \I__4989\ : Span4Mux_h
    port map (
            O => \N__23218\,
            I => \N__23215\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__23215\,
            I => \N__23212\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__23212\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\
        );

    \I__4986\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23206\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__23206\,
            I => \N__23203\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__23203\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\
        );

    \I__4983\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23197\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__23197\,
            I => \ppm_encoder_1.pulses2countZ0Z_6\
        );

    \I__4981\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23191\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23188\
        );

    \I__4979\ : Span4Mux_s2_v
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__4978\ : Span4Mux_v
    port map (
            O => \N__23185\,
            I => \N__23182\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__23182\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\
        );

    \I__4976\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23176\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23173\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__23173\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__23170\,
            I => \N__23167\
        );

    \I__4972\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23164\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__23164\,
            I => \N__23161\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__23161\,
            I => \ppm_encoder_1.pulses2countZ0Z_13\
        );

    \I__4969\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23155\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__23152\
        );

    \I__4967\ : Span4Mux_v
    port map (
            O => \N__23152\,
            I => \N__23149\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__23149\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\
        );

    \I__4965\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23143\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23140\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__23140\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\
        );

    \I__4962\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23128\
        );

    \I__4961\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23128\
        );

    \I__4960\ : InMux
    port map (
            O => \N__23135\,
            I => \N__23128\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23120\
        );

    \I__4958\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23117\
        );

    \I__4957\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23108\
        );

    \I__4956\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23108\
        );

    \I__4955\ : InMux
    port map (
            O => \N__23124\,
            I => \N__23108\
        );

    \I__4954\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23108\
        );

    \I__4953\ : Span4Mux_s3_v
    port map (
            O => \N__23120\,
            I => \N__23101\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23101\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__23108\,
            I => \N__23098\
        );

    \I__4950\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23088\
        );

    \I__4949\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23088\
        );

    \I__4948\ : Span4Mux_h
    port map (
            O => \N__23101\,
            I => \N__23083\
        );

    \I__4947\ : Span4Mux_s3_v
    port map (
            O => \N__23098\,
            I => \N__23083\
        );

    \I__4946\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23072\
        );

    \I__4945\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23072\
        );

    \I__4944\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23072\
        );

    \I__4943\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23072\
        );

    \I__4942\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23072\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__23088\,
            I => \N__23069\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__23083\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__23072\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__4938\ : Odrv12
    port map (
            O => \N__23069\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__4937\ : CEMux
    port map (
            O => \N__23062\,
            I => \N__23057\
        );

    \I__4936\ : CEMux
    port map (
            O => \N__23061\,
            I => \N__23053\
        );

    \I__4935\ : CEMux
    port map (
            O => \N__23060\,
            I => \N__23049\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23046\
        );

    \I__4933\ : CEMux
    port map (
            O => \N__23056\,
            I => \N__23043\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__23053\,
            I => \N__23040\
        );

    \I__4931\ : CEMux
    port map (
            O => \N__23052\,
            I => \N__23037\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__23049\,
            I => \N__23034\
        );

    \I__4929\ : Span4Mux_h
    port map (
            O => \N__23046\,
            I => \N__23029\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__23043\,
            I => \N__23029\
        );

    \I__4927\ : Span4Mux_s3_v
    port map (
            O => \N__23040\,
            I => \N__23026\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__23037\,
            I => \N__23023\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__23034\,
            I => \N__23020\
        );

    \I__4924\ : Span4Mux_s3_v
    port map (
            O => \N__23029\,
            I => \N__23015\
        );

    \I__4923\ : Span4Mux_h
    port map (
            O => \N__23026\,
            I => \N__23015\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__23023\,
            I => \N__23010\
        );

    \I__4921\ : Span4Mux_s2_v
    port map (
            O => \N__23020\,
            I => \N__23010\
        );

    \I__4920\ : Span4Mux_h
    port map (
            O => \N__23015\,
            I => \N__23007\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__23010\,
            I => \ppm_encoder_1.N_590_0\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__23007\,
            I => \ppm_encoder_1.N_590_0\
        );

    \I__4917\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22999\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__22999\,
            I => \ppm_encoder_1.pulses2countZ0Z_14\
        );

    \I__4915\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22991\
        );

    \I__4914\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22988\
        );

    \I__4913\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22985\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__22991\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__22988\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__22985\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__4909\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22975\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__22975\,
            I => \N__22972\
        );

    \I__4907\ : Odrv12
    port map (
            O => \N__22972\,
            I => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\
        );

    \I__4906\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22965\
        );

    \I__4905\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22962\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22959\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__22962\,
            I => \N__22956\
        );

    \I__4902\ : Span12Mux_h
    port map (
            O => \N__22959\,
            I => \N__22952\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__22956\,
            I => \N__22949\
        );

    \I__4900\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22946\
        );

    \I__4899\ : Odrv12
    port map (
            O => \N__22952\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__22949\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__22946\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__4896\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22935\
        );

    \I__4895\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22932\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__22935\,
            I => \N__22929\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__22932\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__4892\ : Odrv12
    port map (
            O => \N__22929\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__4891\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__22921\,
            I => \N__22918\
        );

    \I__4889\ : Span4Mux_s2_v
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__4888\ : Span4Mux_h
    port map (
            O => \N__22915\,
            I => \N__22910\
        );

    \I__4887\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22907\
        );

    \I__4886\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22904\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__22910\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__22907\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__22904\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__22897\,
            I => \N__22893\
        );

    \I__4881\ : CascadeMux
    port map (
            O => \N__22896\,
            I => \N__22890\
        );

    \I__4880\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22887\
        );

    \I__4879\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22884\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22881\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__22884\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__22881\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__4875\ : InMux
    port map (
            O => \N__22876\,
            I => \N__22869\
        );

    \I__4874\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22869\
        );

    \I__4873\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22866\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22863\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__22866\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__4870\ : Odrv12
    port map (
            O => \N__22863\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__4869\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22852\
        );

    \I__4868\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22843\
        );

    \I__4867\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22838\
        );

    \I__4866\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22838\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__22852\,
            I => \N__22835\
        );

    \I__4864\ : InMux
    port map (
            O => \N__22851\,
            I => \N__22832\
        );

    \I__4863\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22829\
        );

    \I__4862\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22823\
        );

    \I__4861\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22823\
        );

    \I__4860\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22820\
        );

    \I__4859\ : CascadeMux
    port map (
            O => \N__22846\,
            I => \N__22817\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__22843\,
            I => \N__22810\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__22838\,
            I => \N__22810\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__22835\,
            I => \N__22803\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__22832\,
            I => \N__22803\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__22829\,
            I => \N__22803\
        );

    \I__4853\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22800\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__22823\,
            I => \N__22795\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22792\
        );

    \I__4850\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22785\
        );

    \I__4849\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22785\
        );

    \I__4848\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22785\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__22810\,
            I => \N__22782\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__22803\,
            I => \N__22779\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__22800\,
            I => \N__22776\
        );

    \I__4844\ : InMux
    port map (
            O => \N__22799\,
            I => \N__22773\
        );

    \I__4843\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22769\
        );

    \I__4842\ : Span4Mux_v
    port map (
            O => \N__22795\,
            I => \N__22764\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__22792\,
            I => \N__22764\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__22785\,
            I => \N__22758\
        );

    \I__4839\ : Span4Mux_v
    port map (
            O => \N__22782\,
            I => \N__22749\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__22779\,
            I => \N__22749\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__22776\,
            I => \N__22749\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__22773\,
            I => \N__22749\
        );

    \I__4835\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22746\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22741\
        );

    \I__4833\ : Span4Mux_h
    port map (
            O => \N__22764\,
            I => \N__22741\
        );

    \I__4832\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22738\
        );

    \I__4831\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22733\
        );

    \I__4830\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22733\
        );

    \I__4829\ : Span4Mux_h
    port map (
            O => \N__22758\,
            I => \N__22730\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__22749\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__22746\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__22741\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__22738\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__22733\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__22730\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__4822\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22714\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__22714\,
            I => \N__22709\
        );

    \I__4820\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22706\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__22712\,
            I => \N__22703\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__22709\,
            I => \N__22700\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__22706\,
            I => \N__22697\
        );

    \I__4816\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22694\
        );

    \I__4815\ : Span4Mux_h
    port map (
            O => \N__22700\,
            I => \N__22689\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__22697\,
            I => \N__22689\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__22694\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__22689\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4811\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22680\
        );

    \I__4810\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22677\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22673\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__22677\,
            I => \N__22670\
        );

    \I__4807\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22667\
        );

    \I__4806\ : Span4Mux_v
    port map (
            O => \N__22673\,
            I => \N__22662\
        );

    \I__4805\ : Span4Mux_h
    port map (
            O => \N__22670\,
            I => \N__22662\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__22667\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__4803\ : Odrv4
    port map (
            O => \N__22662\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__4802\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__22654\,
            I => \ppm_encoder_1.N_301\
        );

    \I__4800\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22648\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__22648\,
            I => \N__22645\
        );

    \I__4798\ : Span4Mux_v
    port map (
            O => \N__22645\,
            I => \N__22642\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__22642\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\
        );

    \I__4796\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22636\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__22636\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\
        );

    \I__4794\ : InMux
    port map (
            O => \N__22633\,
            I => \N__22628\
        );

    \I__4793\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22625\
        );

    \I__4792\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22622\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__22628\,
            I => \N__22619\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__22625\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__22622\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__22619\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__4787\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22607\
        );

    \I__4786\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22604\
        );

    \I__4785\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22601\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__22607\,
            I => \N__22598\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__22604\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__22601\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__22598\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__4780\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22586\
        );

    \I__4779\ : InMux
    port map (
            O => \N__22590\,
            I => \N__22583\
        );

    \I__4778\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22580\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22577\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__22583\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__22580\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__4774\ : Odrv12
    port map (
            O => \N__22577\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__4773\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22565\
        );

    \I__4772\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22562\
        );

    \I__4771\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22559\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22556\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__22562\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__22559\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__4767\ : Odrv4
    port map (
            O => \N__22556\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__22549\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\
        );

    \I__4765\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22543\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22540\
        );

    \I__4763\ : Span4Mux_s2_v
    port map (
            O => \N__22540\,
            I => \N__22537\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__22537\,
            I => \ppm_encoder_1.N_144_17\
        );

    \I__4761\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__22528\,
            I => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\
        );

    \I__4758\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__22519\,
            I => \N__22516\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__22516\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\
        );

    \I__4754\ : CascadeMux
    port map (
            O => \N__22513\,
            I => \ppm_encoder_1.N_144_17_cascade_\
        );

    \I__4753\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22507\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__22507\,
            I => \N__22504\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__4750\ : Span4Mux_v
    port map (
            O => \N__22501\,
            I => \N__22498\
        );

    \I__4749\ : Odrv4
    port map (
            O => \N__22498\,
            I => \ppm_encoder_1.N_144\
        );

    \I__4748\ : InMux
    port map (
            O => \N__22495\,
            I => \N__22492\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__22492\,
            I => \N__22489\
        );

    \I__4746\ : Span4Mux_h
    port map (
            O => \N__22489\,
            I => \N__22486\
        );

    \I__4745\ : Span4Mux_v
    port map (
            O => \N__22486\,
            I => \N__22483\
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__22483\,
            I => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\
        );

    \I__4743\ : InMux
    port map (
            O => \N__22480\,
            I => \ppm_encoder_1.un1_aileron_cry_6\
        );

    \I__4742\ : InMux
    port map (
            O => \N__22477\,
            I => \N__22474\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__22474\,
            I => \N__22471\
        );

    \I__4740\ : Span12Mux_s8_h
    port map (
            O => \N__22471\,
            I => \N__22468\
        );

    \I__4739\ : Odrv12
    port map (
            O => \N__22468\,
            I => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\
        );

    \I__4738\ : InMux
    port map (
            O => \N__22465\,
            I => \ppm_encoder_1.un1_aileron_cry_7\
        );

    \I__4737\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22459\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__22459\,
            I => \N__22456\
        );

    \I__4735\ : Odrv4
    port map (
            O => \N__22456\,
            I => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\
        );

    \I__4734\ : InMux
    port map (
            O => \N__22453\,
            I => \ppm_encoder_1.un1_aileron_cry_8\
        );

    \I__4733\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22447\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__22447\,
            I => \N__22444\
        );

    \I__4731\ : Span4Mux_h
    port map (
            O => \N__22444\,
            I => \N__22441\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__22441\,
            I => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\
        );

    \I__4729\ : InMux
    port map (
            O => \N__22438\,
            I => \ppm_encoder_1.un1_aileron_cry_9\
        );

    \I__4728\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__22429\,
            I => \N__22426\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__22426\,
            I => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\
        );

    \I__4724\ : InMux
    port map (
            O => \N__22423\,
            I => \ppm_encoder_1.un1_aileron_cry_10\
        );

    \I__4723\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22417\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22414\
        );

    \I__4721\ : Span4Mux_h
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__22411\,
            I => \N__22408\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__22408\,
            I => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\
        );

    \I__4718\ : InMux
    port map (
            O => \N__22405\,
            I => \ppm_encoder_1.un1_aileron_cry_11\
        );

    \I__4717\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22399\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__22399\,
            I => \N__22396\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__22396\,
            I => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\
        );

    \I__4714\ : InMux
    port map (
            O => \N__22393\,
            I => \ppm_encoder_1.un1_aileron_cry_12\
        );

    \I__4713\ : InMux
    port map (
            O => \N__22390\,
            I => \bfn_8_20_0_\
        );

    \I__4712\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22383\
        );

    \I__4711\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22380\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22377\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__22380\,
            I => \N__22374\
        );

    \I__4708\ : Span4Mux_h
    port map (
            O => \N__22377\,
            I => \N__22371\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__22374\,
            I => \N__22368\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__22371\,
            I => \N__22365\
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__22368\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__22365\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__4703\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22357\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__4701\ : Span4Mux_h
    port map (
            O => \N__22354\,
            I => \N__22351\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__22351\,
            I => \Commands_frame_decoder.state_1_RNO_4Z0Z_0\
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__22348\,
            I => \N__22345\
        );

    \I__4698\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22342\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__4696\ : Span4Mux_h
    port map (
            O => \N__22339\,
            I => \N__22334\
        );

    \I__4695\ : InMux
    port map (
            O => \N__22338\,
            I => \N__22331\
        );

    \I__4694\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22327\
        );

    \I__4693\ : Span4Mux_h
    port map (
            O => \N__22334\,
            I => \N__22324\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22321\
        );

    \I__4691\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22318\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__22327\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__22324\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__22321\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__22318\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4686\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22306\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__22306\,
            I => \N__22302\
        );

    \I__4684\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22299\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__22302\,
            I => \N__22295\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__22299\,
            I => \N__22292\
        );

    \I__4681\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22289\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__22295\,
            I => \Commands_frame_decoder.WDT8lt14_0\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__22292\,
            I => \Commands_frame_decoder.WDT8lt14_0\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__22289\,
            I => \Commands_frame_decoder.WDT8lt14_0\
        );

    \I__4677\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22279\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22276\
        );

    \I__4675\ : Odrv12
    port map (
            O => \N__22276\,
            I => \uart_pc.un1_state_2_0_a3_0\
        );

    \I__4674\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22268\
        );

    \I__4673\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22265\
        );

    \I__4672\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22262\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__22268\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__22265\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__22262\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__4668\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22252\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__22252\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_2\
        );

    \I__4666\ : InMux
    port map (
            O => \N__22249\,
            I => \uart_pc.un4_timer_Count_1_cry_1\
        );

    \I__4665\ : InMux
    port map (
            O => \N__22246\,
            I => \uart_pc.un4_timer_Count_1_cry_2\
        );

    \I__4664\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22232\
        );

    \I__4663\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22232\
        );

    \I__4662\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22227\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__22240\,
            I => \N__22224\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__22239\,
            I => \N__22221\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__22238\,
            I => \N__22218\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__22237\,
            I => \N__22215\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__22232\,
            I => \N__22212\
        );

    \I__4656\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22207\
        );

    \I__4655\ : InMux
    port map (
            O => \N__22230\,
            I => \N__22207\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22204\
        );

    \I__4653\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22199\
        );

    \I__4652\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22199\
        );

    \I__4651\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22194\
        );

    \I__4650\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22194\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__22212\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__22207\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__22204\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__22199\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__22194\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__4644\ : InMux
    port map (
            O => \N__22183\,
            I => \uart_pc.un4_timer_Count_1_cry_3\
        );

    \I__4643\ : InMux
    port map (
            O => \N__22180\,
            I => \N__22177\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__22177\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_4\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__22174\,
            I => \N__22170\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__22173\,
            I => \N__22166\
        );

    \I__4639\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22162\
        );

    \I__4638\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22155\
        );

    \I__4637\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22155\
        );

    \I__4636\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22155\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__22162\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__22155\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__4633\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22144\
        );

    \I__4632\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22144\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__22141\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__4628\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__22129\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_1\
        );

    \I__4625\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22123\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__22123\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_3\
        );

    \I__4623\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22113\
        );

    \I__4622\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22110\
        );

    \I__4621\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22107\
        );

    \I__4620\ : InMux
    port map (
            O => \N__22117\,
            I => \N__22102\
        );

    \I__4619\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22102\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__22113\,
            I => \uart_pc.N_143\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__22110\,
            I => \uart_pc.N_143\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__22107\,
            I => \uart_pc.N_143\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__22102\,
            I => \uart_pc.N_143\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__22093\,
            I => \N__22088\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__22092\,
            I => \N__22085\
        );

    \I__4612\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22080\
        );

    \I__4611\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22077\
        );

    \I__4610\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22074\
        );

    \I__4609\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22069\
        );

    \I__4608\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22069\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__22080\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__22077\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__22074\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__22069\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4603\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__22047\
        );

    \I__4601\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22044\
        );

    \I__4600\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22035\
        );

    \I__4599\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22035\
        );

    \I__4598\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22035\
        );

    \I__4597\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22035\
        );

    \I__4596\ : InMux
    port map (
            O => \N__22051\,
            I => \N__22030\
        );

    \I__4595\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22030\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__22047\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__22044\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__22035\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__22030\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22021\,
            I => \N__22016\
        );

    \I__4589\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22011\
        );

    \I__4588\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22008\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__22005\
        );

    \I__4586\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22000\
        );

    \I__4585\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22000\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__22011\,
            I => \N__21995\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__22008\,
            I => \N__21992\
        );

    \I__4582\ : Span4Mux_v
    port map (
            O => \N__22005\,
            I => \N__21986\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__22000\,
            I => \N__21986\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__21999\,
            I => \N__21982\
        );

    \I__4579\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21979\
        );

    \I__4578\ : Span4Mux_h
    port map (
            O => \N__21995\,
            I => \N__21976\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__21992\,
            I => \N__21973\
        );

    \I__4576\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21970\
        );

    \I__4575\ : Span4Mux_h
    port map (
            O => \N__21986\,
            I => \N__21967\
        );

    \I__4574\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21962\
        );

    \I__4573\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21962\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__21979\,
            I => \N__21959\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__21976\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__21973\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__21970\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__21967\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__21962\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__4566\ : Odrv12
    port map (
            O => \N__21959\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__4565\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21938\
        );

    \I__4564\ : InMux
    port map (
            O => \N__21945\,
            I => \N__21938\
        );

    \I__4563\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21935\
        );

    \I__4562\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21932\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__21938\,
            I => \N__21928\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__21935\,
            I => \N__21923\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__21932\,
            I => \N__21923\
        );

    \I__4558\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21919\
        );

    \I__4557\ : Span4Mux_h
    port map (
            O => \N__21928\,
            I => \N__21914\
        );

    \I__4556\ : Span4Mux_h
    port map (
            O => \N__21923\,
            I => \N__21911\
        );

    \I__4555\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21908\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21905\
        );

    \I__4553\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21900\
        );

    \I__4552\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21900\
        );

    \I__4551\ : Odrv4
    port map (
            O => \N__21914\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__4550\ : Odrv4
    port map (
            O => \N__21911\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__21908\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__4548\ : Odrv12
    port map (
            O => \N__21905\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__21900\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__4546\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21882\
        );

    \I__4545\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21882\
        );

    \I__4544\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21877\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21873\
        );

    \I__4542\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21870\
        );

    \I__4541\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21867\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__21877\,
            I => \N__21864\
        );

    \I__4539\ : InMux
    port map (
            O => \N__21876\,
            I => \N__21861\
        );

    \I__4538\ : Span4Mux_h
    port map (
            O => \N__21873\,
            I => \N__21858\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__21870\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__21867\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__21864\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__21861\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__4533\ : Odrv4
    port map (
            O => \N__21858\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__4532\ : InMux
    port map (
            O => \N__21847\,
            I => \N__21844\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__21844\,
            I => \uart_drone.data_Auxce_0_0_2\
        );

    \I__4530\ : InMux
    port map (
            O => \N__21841\,
            I => \N__21837\
        );

    \I__4529\ : CascadeMux
    port map (
            O => \N__21840\,
            I => \N__21834\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__21837\,
            I => \N__21831\
        );

    \I__4527\ : InMux
    port map (
            O => \N__21834\,
            I => \N__21828\
        );

    \I__4526\ : Odrv12
    port map (
            O => \N__21831\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__21828\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__4524\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__4522\ : Odrv12
    port map (
            O => \N__21817\,
            I => \uart_drone.data_Auxce_0_3\
        );

    \I__4521\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21810\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__21813\,
            I => \N__21807\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__21810\,
            I => \N__21804\
        );

    \I__4518\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21801\
        );

    \I__4517\ : Odrv12
    port map (
            O => \N__21804\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__21801\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__4515\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21781\
        );

    \I__4514\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21781\
        );

    \I__4513\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21781\
        );

    \I__4512\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21781\
        );

    \I__4511\ : InMux
    port map (
            O => \N__21792\,
            I => \N__21781\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__21781\,
            I => \N__21778\
        );

    \I__4509\ : Span4Mux_h
    port map (
            O => \N__21778\,
            I => \N__21772\
        );

    \I__4508\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21765\
        );

    \I__4507\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21765\
        );

    \I__4506\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21765\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__21772\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__21765\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__4503\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21757\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__21757\,
            I => \N__21751\
        );

    \I__4501\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21743\
        );

    \I__4500\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21733\
        );

    \I__4499\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21733\
        );

    \I__4498\ : Span4Mux_v
    port map (
            O => \N__21751\,
            I => \N__21730\
        );

    \I__4497\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21727\
        );

    \I__4496\ : IoInMux
    port map (
            O => \N__21749\,
            I => \N__21724\
        );

    \I__4495\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21721\
        );

    \I__4494\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21716\
        );

    \I__4493\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21716\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__21743\,
            I => \N__21713\
        );

    \I__4491\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21706\
        );

    \I__4490\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21706\
        );

    \I__4489\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21706\
        );

    \I__4488\ : InMux
    port map (
            O => \N__21739\,
            I => \N__21701\
        );

    \I__4487\ : InMux
    port map (
            O => \N__21738\,
            I => \N__21701\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__21733\,
            I => \N__21694\
        );

    \I__4485\ : Span4Mux_h
    port map (
            O => \N__21730\,
            I => \N__21694\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21694\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__21724\,
            I => \N__21691\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__21721\,
            I => \N__21686\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21686\
        );

    \I__4480\ : Span4Mux_h
    port map (
            O => \N__21713\,
            I => \N__21683\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__21706\,
            I => \N__21676\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21676\
        );

    \I__4477\ : Sp12to4
    port map (
            O => \N__21694\,
            I => \N__21676\
        );

    \I__4476\ : Span4Mux_s1_v
    port map (
            O => \N__21691\,
            I => \N__21673\
        );

    \I__4475\ : Span12Mux_v
    port map (
            O => \N__21686\,
            I => \N__21668\
        );

    \I__4474\ : Sp12to4
    port map (
            O => \N__21683\,
            I => \N__21668\
        );

    \I__4473\ : Span12Mux_v
    port map (
            O => \N__21676\,
            I => \N__21665\
        );

    \I__4472\ : Sp12to4
    port map (
            O => \N__21673\,
            I => \N__21660\
        );

    \I__4471\ : Span12Mux_v
    port map (
            O => \N__21668\,
            I => \N__21660\
        );

    \I__4470\ : Odrv12
    port map (
            O => \N__21665\,
            I => uart_drone_input_debug_c
        );

    \I__4469\ : Odrv12
    port map (
            O => \N__21660\,
            I => uart_drone_input_debug_c
        );

    \I__4468\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21651\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__21654\,
            I => \N__21648\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__21651\,
            I => \N__21645\
        );

    \I__4465\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21642\
        );

    \I__4464\ : Odrv12
    port map (
            O => \N__21645\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__21642\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__4462\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__21634\,
            I => \uart_drone.data_Auxce_0_0_4\
        );

    \I__4460\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21626\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__21630\,
            I => \N__21623\
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__21629\,
            I => \N__21620\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__21626\,
            I => \N__21616\
        );

    \I__4456\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21611\
        );

    \I__4455\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21611\
        );

    \I__4454\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21608\
        );

    \I__4453\ : Span4Mux_h
    port map (
            O => \N__21616\,
            I => \N__21603\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__21611\,
            I => \N__21603\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__21608\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__21603\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__4448\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21592\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__21589\,
            I => \uart_drone.N_145\
        );

    \I__4445\ : SRMux
    port map (
            O => \N__21586\,
            I => \N__21583\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__21583\,
            I => \N__21580\
        );

    \I__4443\ : Span4Mux_h
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__21577\,
            I => \N__21573\
        );

    \I__4441\ : SRMux
    port map (
            O => \N__21576\,
            I => \N__21570\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__21573\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__21570\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__4438\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21561\
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__21564\,
            I => \N__21558\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21554\
        );

    \I__4435\ : InMux
    port map (
            O => \N__21558\,
            I => \N__21547\
        );

    \I__4434\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21547\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__21554\,
            I => \N__21544\
        );

    \I__4432\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21539\
        );

    \I__4431\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21539\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__21547\,
            I => \uart_drone.N_143\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__21544\,
            I => \uart_drone.N_143\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__21539\,
            I => \uart_drone.N_143\
        );

    \I__4427\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21526\
        );

    \I__4426\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21526\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__21526\,
            I => \N__21523\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__21523\,
            I => \uart_drone.N_144_1\
        );

    \I__4423\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21517\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__21517\,
            I => \N__21514\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__21514\,
            I => \scaler_2.N_521_i_l_ofxZ0\
        );

    \I__4420\ : InMux
    port map (
            O => \N__21511\,
            I => \bfn_8_14_0_\
        );

    \I__4419\ : InMux
    port map (
            O => \N__21508\,
            I => \scaler_2.un3_source_data_0_cry_8\
        );

    \I__4418\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21501\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__21504\,
            I => \N__21498\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21495\
        );

    \I__4415\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21492\
        );

    \I__4414\ : Odrv12
    port map (
            O => \N__21495\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__21492\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__4412\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21484\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__21484\,
            I => \N__21480\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__21483\,
            I => \N__21477\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__21480\,
            I => \N__21474\
        );

    \I__4408\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21471\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__21474\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__21471\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__4405\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21463\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__21463\,
            I => \N__21460\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__21460\,
            I => \frame_decoder_CH2data_1\
        );

    \I__4402\ : InMux
    port map (
            O => \N__21457\,
            I => \scaler_2.un3_source_data_0_cry_0\
        );

    \I__4401\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21451\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__21451\,
            I => \frame_decoder_CH2data_2\
        );

    \I__4399\ : InMux
    port map (
            O => \N__21448\,
            I => \scaler_2.un3_source_data_0_cry_1\
        );

    \I__4398\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21442\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__21442\,
            I => \frame_decoder_CH2data_3\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__21439\,
            I => \N__21436\
        );

    \I__4395\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21433\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__21433\,
            I => \frame_decoder_OFF2data_3\
        );

    \I__4393\ : InMux
    port map (
            O => \N__21430\,
            I => \scaler_2.un3_source_data_0_cry_2\
        );

    \I__4392\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21424\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21421\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__21421\,
            I => \frame_decoder_CH2data_4\
        );

    \I__4389\ : InMux
    port map (
            O => \N__21418\,
            I => \scaler_2.un3_source_data_0_cry_3\
        );

    \I__4388\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21412\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__21412\,
            I => \frame_decoder_CH2data_5\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__21409\,
            I => \N__21406\
        );

    \I__4385\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21403\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__21403\,
            I => \frame_decoder_OFF2data_5\
        );

    \I__4383\ : InMux
    port map (
            O => \N__21400\,
            I => \scaler_2.un3_source_data_0_cry_4\
        );

    \I__4382\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21394\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__21394\,
            I => \frame_decoder_CH2data_6\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__21391\,
            I => \N__21388\
        );

    \I__4379\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21385\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__21385\,
            I => \N__21382\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__21382\,
            I => \frame_decoder_OFF2data_6\
        );

    \I__4376\ : InMux
    port map (
            O => \N__21379\,
            I => \scaler_2.un3_source_data_0_cry_5\
        );

    \I__4375\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21373\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__21373\,
            I => \N__21370\
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__21370\,
            I => \scaler_2.un3_source_data_0_axb_7\
        );

    \I__4372\ : InMux
    port map (
            O => \N__21367\,
            I => \scaler_2.un3_source_data_0_cry_6\
        );

    \I__4371\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21361\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__21361\,
            I => \uart_drone_sync.aux_0__0_Z0Z_0\
        );

    \I__4369\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21355\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__21355\,
            I => \uart_drone_sync.aux_1__0_Z0Z_0\
        );

    \I__4367\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21349\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__21349\,
            I => \uart_drone_sync.aux_2__0_Z0Z_0\
        );

    \I__4365\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21343\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__21343\,
            I => \uart_drone_sync.aux_3__0_Z0Z_0\
        );

    \I__4363\ : CEMux
    port map (
            O => \N__21340\,
            I => \N__21335\
        );

    \I__4362\ : CEMux
    port map (
            O => \N__21339\,
            I => \N__21332\
        );

    \I__4361\ : CEMux
    port map (
            O => \N__21338\,
            I => \N__21329\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21326\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21321\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N__21321\
        );

    \I__4357\ : Span4Mux_h
    port map (
            O => \N__21326\,
            I => \N__21318\
        );

    \I__4356\ : Span4Mux_v
    port map (
            O => \N__21321\,
            I => \N__21315\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__21318\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__21315\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__4353\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21304\
        );

    \I__4352\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21304\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__21304\,
            I => \frame_decoder_CH2data_7\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__21301\,
            I => \N__21298\
        );

    \I__4349\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21291\
        );

    \I__4348\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21291\
        );

    \I__4347\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21288\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__21291\,
            I => \N__21285\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__21288\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__4344\ : Odrv12
    port map (
            O => \N__21285\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__4343\ : InMux
    port map (
            O => \N__21280\,
            I => \ppm_encoder_1.un1_counter_13_cry_10\
        );

    \I__4342\ : InMux
    port map (
            O => \N__21277\,
            I => \ppm_encoder_1.un1_counter_13_cry_11\
        );

    \I__4341\ : InMux
    port map (
            O => \N__21274\,
            I => \ppm_encoder_1.un1_counter_13_cry_12\
        );

    \I__4340\ : InMux
    port map (
            O => \N__21271\,
            I => \ppm_encoder_1.un1_counter_13_cry_13\
        );

    \I__4339\ : InMux
    port map (
            O => \N__21268\,
            I => \ppm_encoder_1.un1_counter_13_cry_14\
        );

    \I__4338\ : InMux
    port map (
            O => \N__21265\,
            I => \bfn_7_30_0_\
        );

    \I__4337\ : InMux
    port map (
            O => \N__21262\,
            I => \ppm_encoder_1.un1_counter_13_cry_16\
        );

    \I__4336\ : InMux
    port map (
            O => \N__21259\,
            I => \ppm_encoder_1.un1_counter_13_cry_17\
        );

    \I__4335\ : SRMux
    port map (
            O => \N__21256\,
            I => \N__21247\
        );

    \I__4334\ : SRMux
    port map (
            O => \N__21255\,
            I => \N__21247\
        );

    \I__4333\ : SRMux
    port map (
            O => \N__21254\,
            I => \N__21247\
        );

    \I__4332\ : GlobalMux
    port map (
            O => \N__21247\,
            I => \N__21244\
        );

    \I__4331\ : gio2CtrlBuf
    port map (
            O => \N__21244\,
            I => \ppm_encoder_1.N_168_g\
        );

    \I__4330\ : InMux
    port map (
            O => \N__21241\,
            I => \N__21238\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__21238\,
            I => uart_input_drone_c
        );

    \I__4328\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__4326\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21221\
        );

    \I__4325\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21221\
        );

    \I__4324\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21218\
        );

    \I__4323\ : Span4Mux_h
    port map (
            O => \N__21226\,
            I => \N__21215\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21212\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__21218\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__21215\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__21212\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4318\ : InMux
    port map (
            O => \N__21205\,
            I => \ppm_encoder_1.un1_counter_13_cry_1\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__21202\,
            I => \N__21199\
        );

    \I__4316\ : InMux
    port map (
            O => \N__21199\,
            I => \N__21195\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__21198\,
            I => \N__21192\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__21195\,
            I => \N__21187\
        );

    \I__4313\ : InMux
    port map (
            O => \N__21192\,
            I => \N__21182\
        );

    \I__4312\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21182\
        );

    \I__4311\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21179\
        );

    \I__4310\ : Span4Mux_h
    port map (
            O => \N__21187\,
            I => \N__21176\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__21182\,
            I => \N__21173\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__21179\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__21176\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__21173\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4305\ : InMux
    port map (
            O => \N__21166\,
            I => \ppm_encoder_1.un1_counter_13_cry_2\
        );

    \I__4304\ : InMux
    port map (
            O => \N__21163\,
            I => \ppm_encoder_1.un1_counter_13_cry_3\
        );

    \I__4303\ : InMux
    port map (
            O => \N__21160\,
            I => \ppm_encoder_1.un1_counter_13_cry_4\
        );

    \I__4302\ : InMux
    port map (
            O => \N__21157\,
            I => \ppm_encoder_1.un1_counter_13_cry_5\
        );

    \I__4301\ : InMux
    port map (
            O => \N__21154\,
            I => \ppm_encoder_1.un1_counter_13_cry_6\
        );

    \I__4300\ : InMux
    port map (
            O => \N__21151\,
            I => \bfn_7_29_0_\
        );

    \I__4299\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21143\
        );

    \I__4298\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21140\
        );

    \I__4297\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21137\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__21143\,
            I => \N__21132\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21132\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__21137\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__4293\ : Odrv12
    port map (
            O => \N__21132\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__4292\ : InMux
    port map (
            O => \N__21127\,
            I => \ppm_encoder_1.un1_counter_13_cry_8\
        );

    \I__4291\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21117\
        );

    \I__4290\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21117\
        );

    \I__4289\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21114\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__21117\,
            I => \N__21111\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__21114\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__21111\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__4285\ : InMux
    port map (
            O => \N__21106\,
            I => \ppm_encoder_1.un1_counter_13_cry_9\
        );

    \I__4284\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21099\
        );

    \I__4283\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21096\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21093\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__21096\,
            I => \N__21090\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__21093\,
            I => \N__21084\
        );

    \I__4279\ : Span4Mux_v
    port map (
            O => \N__21090\,
            I => \N__21084\
        );

    \I__4278\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21081\
        );

    \I__4277\ : Odrv4
    port map (
            O => \N__21084\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__21081\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__21076\,
            I => \N__21073\
        );

    \I__4274\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21069\
        );

    \I__4273\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21066\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__21069\,
            I => \N__21062\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21059\
        );

    \I__4270\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21056\
        );

    \I__4269\ : Span4Mux_h
    port map (
            O => \N__21062\,
            I => \N__21053\
        );

    \I__4268\ : Span4Mux_h
    port map (
            O => \N__21059\,
            I => \N__21050\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__21056\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__21053\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4265\ : Odrv4
    port map (
            O => \N__21050\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4264\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21039\
        );

    \I__4263\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21036\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__21039\,
            I => \N__21033\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__21036\,
            I => \N__21029\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__21033\,
            I => \N__21026\
        );

    \I__4259\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21023\
        );

    \I__4258\ : Odrv12
    port map (
            O => \N__21029\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__21026\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__21023\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4255\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21011\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__21015\,
            I => \N__21008\
        );

    \I__4253\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21005\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__21002\
        );

    \I__4251\ : InMux
    port map (
            O => \N__21008\,
            I => \N__20999\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__20996\
        );

    \I__4249\ : Span4Mux_s3_h
    port map (
            O => \N__21002\,
            I => \N__20993\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20990\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__20996\,
            I => \N__20985\
        );

    \I__4246\ : Span4Mux_h
    port map (
            O => \N__20993\,
            I => \N__20985\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__20990\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__20985\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__20980\,
            I => \N__20976\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__20979\,
            I => \N__20973\
        );

    \I__4241\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20969\
        );

    \I__4240\ : InMux
    port map (
            O => \N__20973\,
            I => \N__20966\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__20972\,
            I => \N__20963\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__20969\,
            I => \N__20952\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__20966\,
            I => \N__20952\
        );

    \I__4236\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20949\
        );

    \I__4235\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20944\
        );

    \I__4234\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20939\
        );

    \I__4233\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20939\
        );

    \I__4232\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20935\
        );

    \I__4231\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20928\
        );

    \I__4230\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20925\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__20952\,
            I => \N__20915\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20915\
        );

    \I__4227\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20912\
        );

    \I__4226\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20909\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__20944\,
            I => \N__20904\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__20939\,
            I => \N__20904\
        );

    \I__4223\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20901\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__20935\,
            I => \N__20898\
        );

    \I__4221\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20895\
        );

    \I__4220\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20892\
        );

    \I__4219\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20889\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__20931\,
            I => \N__20886\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__20928\,
            I => \N__20882\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20879\
        );

    \I__4215\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20872\
        );

    \I__4214\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20872\
        );

    \I__4213\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20872\
        );

    \I__4212\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20869\
        );

    \I__4211\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20866\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__20915\,
            I => \N__20861\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__20912\,
            I => \N__20861\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20856\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__20904\,
            I => \N__20856\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__20901\,
            I => \N__20849\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__20898\,
            I => \N__20849\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__20895\,
            I => \N__20849\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__20892\,
            I => \N__20844\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20844\
        );

    \I__4201\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20839\
        );

    \I__4200\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20839\
        );

    \I__4199\ : Span12Mux_v
    port map (
            O => \N__20882\,
            I => \N__20828\
        );

    \I__4198\ : Span12Mux_s3_v
    port map (
            O => \N__20879\,
            I => \N__20828\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__20872\,
            I => \N__20828\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__20869\,
            I => \N__20828\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20828\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__20861\,
            I => \N__20825\
        );

    \I__4193\ : Span4Mux_h
    port map (
            O => \N__20856\,
            I => \N__20820\
        );

    \I__4192\ : Span4Mux_v
    port map (
            O => \N__20849\,
            I => \N__20820\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__20844\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__20839\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__4189\ : Odrv12
    port map (
            O => \N__20828\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__20825\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__20820\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__20809\,
            I => \N__20803\
        );

    \I__4185\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20800\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__20807\,
            I => \N__20794\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__20806\,
            I => \N__20787\
        );

    \I__4182\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20770\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__20800\,
            I => \N__20767\
        );

    \I__4180\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20760\
        );

    \I__4179\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20760\
        );

    \I__4178\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20760\
        );

    \I__4177\ : InMux
    port map (
            O => \N__20794\,
            I => \N__20756\
        );

    \I__4176\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20747\
        );

    \I__4175\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20747\
        );

    \I__4174\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20747\
        );

    \I__4173\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20747\
        );

    \I__4172\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20738\
        );

    \I__4171\ : InMux
    port map (
            O => \N__20786\,
            I => \N__20738\
        );

    \I__4170\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20738\
        );

    \I__4169\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20738\
        );

    \I__4168\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20731\
        );

    \I__4167\ : InMux
    port map (
            O => \N__20782\,
            I => \N__20731\
        );

    \I__4166\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20731\
        );

    \I__4165\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20722\
        );

    \I__4164\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20722\
        );

    \I__4163\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20722\
        );

    \I__4162\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20722\
        );

    \I__4161\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20715\
        );

    \I__4160\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20715\
        );

    \I__4159\ : InMux
    port map (
            O => \N__20774\,
            I => \N__20715\
        );

    \I__4158\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20710\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__20770\,
            I => \N__20703\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__20767\,
            I => \N__20703\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__20760\,
            I => \N__20703\
        );

    \I__4154\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20699\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20694\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__20747\,
            I => \N__20694\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20682\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20679\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20676\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__20715\,
            I => \N__20673\
        );

    \I__4147\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20668\
        );

    \I__4146\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20668\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__20710\,
            I => \N__20663\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__20703\,
            I => \N__20660\
        );

    \I__4143\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20657\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__20699\,
            I => \N__20652\
        );

    \I__4141\ : Span4Mux_s2_v
    port map (
            O => \N__20694\,
            I => \N__20652\
        );

    \I__4140\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20641\
        );

    \I__4139\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20641\
        );

    \I__4138\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20641\
        );

    \I__4137\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20641\
        );

    \I__4136\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20641\
        );

    \I__4135\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20638\
        );

    \I__4134\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20635\
        );

    \I__4133\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20630\
        );

    \I__4132\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20630\
        );

    \I__4131\ : Span4Mux_v
    port map (
            O => \N__20682\,
            I => \N__20619\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__20679\,
            I => \N__20619\
        );

    \I__4129\ : Span4Mux_h
    port map (
            O => \N__20676\,
            I => \N__20619\
        );

    \I__4128\ : Span4Mux_v
    port map (
            O => \N__20673\,
            I => \N__20619\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__20668\,
            I => \N__20619\
        );

    \I__4126\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20614\
        );

    \I__4125\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20614\
        );

    \I__4124\ : Odrv12
    port map (
            O => \N__20663\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__20660\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__20657\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__20652\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__20641\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__20638\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__20635\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__20630\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4116\ : Odrv4
    port map (
            O => \N__20619\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__20614\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__20593\,
            I => \N__20590\
        );

    \I__4113\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20587\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__20587\,
            I => \N__20584\
        );

    \I__4111\ : Span4Mux_s3_h
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__4110\ : Span4Mux_h
    port map (
            O => \N__20581\,
            I => \N__20578\
        );

    \I__4109\ : Odrv4
    port map (
            O => \N__20578\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__4108\ : CascadeMux
    port map (
            O => \N__20575\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__20572\,
            I => \N__20565\
        );

    \I__4106\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20560\
        );

    \I__4105\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20560\
        );

    \I__4104\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20556\
        );

    \I__4103\ : InMux
    port map (
            O => \N__20568\,
            I => \N__20546\
        );

    \I__4102\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20546\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__20560\,
            I => \N__20541\
        );

    \I__4100\ : InMux
    port map (
            O => \N__20559\,
            I => \N__20538\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__20556\,
            I => \N__20534\
        );

    \I__4098\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20531\
        );

    \I__4097\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20528\
        );

    \I__4096\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20521\
        );

    \I__4095\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20521\
        );

    \I__4094\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20521\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__20546\,
            I => \N__20518\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__20545\,
            I => \N__20510\
        );

    \I__4091\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20507\
        );

    \I__4090\ : Span4Mux_s2_v
    port map (
            O => \N__20541\,
            I => \N__20504\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__20538\,
            I => \N__20501\
        );

    \I__4088\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20498\
        );

    \I__4087\ : Span4Mux_v
    port map (
            O => \N__20534\,
            I => \N__20491\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__20531\,
            I => \N__20491\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20491\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__20521\,
            I => \N__20486\
        );

    \I__4083\ : Span4Mux_h
    port map (
            O => \N__20518\,
            I => \N__20486\
        );

    \I__4082\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20483\
        );

    \I__4081\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20478\
        );

    \I__4080\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20478\
        );

    \I__4079\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20475\
        );

    \I__4078\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20470\
        );

    \I__4077\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20470\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__20507\,
            I => \N__20467\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__20504\,
            I => \N__20462\
        );

    \I__4074\ : Span4Mux_h
    port map (
            O => \N__20501\,
            I => \N__20462\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__20498\,
            I => \N__20455\
        );

    \I__4072\ : Span4Mux_h
    port map (
            O => \N__20491\,
            I => \N__20455\
        );

    \I__4071\ : Span4Mux_v
    port map (
            O => \N__20486\,
            I => \N__20455\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__20483\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__20478\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__20475\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__20470\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__4066\ : Odrv12
    port map (
            O => \N__20467\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__20462\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__20455\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__4063\ : InMux
    port map (
            O => \N__20440\,
            I => \N__20435\
        );

    \I__4062\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20430\
        );

    \I__4061\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20430\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__20435\,
            I => \N__20427\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__20430\,
            I => \N__20424\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__20427\,
            I => \N__20419\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__20424\,
            I => \N__20419\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__20419\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__4055\ : CascadeMux
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__4054\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20409\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__20412\,
            I => \N__20405\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20402\
        );

    \I__4051\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20399\
        );

    \I__4050\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20396\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__20402\,
            I => \N__20393\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__20399\,
            I => \N__20390\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__20396\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__20393\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__4045\ : Odrv12
    port map (
            O => \N__20390\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__20383\,
            I => \N__20376\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__20382\,
            I => \N__20373\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__20381\,
            I => \N__20370\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__20380\,
            I => \N__20366\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__20379\,
            I => \N__20362\
        );

    \I__4039\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20355\
        );

    \I__4038\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20355\
        );

    \I__4037\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20352\
        );

    \I__4036\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20346\
        );

    \I__4035\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20346\
        );

    \I__4034\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20340\
        );

    \I__4033\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20340\
        );

    \I__4032\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20337\
        );

    \I__4031\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20334\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20331\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__20352\,
            I => \N__20328\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__20351\,
            I => \N__20324\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__20346\,
            I => \N__20318\
        );

    \I__4026\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20315\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__20340\,
            I => \N__20312\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__20337\,
            I => \N__20309\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__20334\,
            I => \N__20302\
        );

    \I__4022\ : Span4Mux_s3_v
    port map (
            O => \N__20331\,
            I => \N__20302\
        );

    \I__4021\ : Span4Mux_s2_h
    port map (
            O => \N__20328\,
            I => \N__20302\
        );

    \I__4020\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20293\
        );

    \I__4019\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20293\
        );

    \I__4018\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20293\
        );

    \I__4017\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20293\
        );

    \I__4016\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20290\
        );

    \I__4015\ : Span4Mux_v
    port map (
            O => \N__20318\,
            I => \N__20285\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__20315\,
            I => \N__20285\
        );

    \I__4013\ : Span4Mux_h
    port map (
            O => \N__20312\,
            I => \N__20282\
        );

    \I__4012\ : Span4Mux_h
    port map (
            O => \N__20309\,
            I => \N__20277\
        );

    \I__4011\ : Span4Mux_h
    port map (
            O => \N__20302\,
            I => \N__20277\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__20293\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__20290\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__20285\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__20282\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__20277\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__4005\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20262\
        );

    \I__4004\ : CascadeMux
    port map (
            O => \N__20265\,
            I => \N__20259\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__20262\,
            I => \N__20256\
        );

    \I__4002\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20253\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__20256\,
            I => \ppm_encoder_1.N_590_i\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__20253\,
            I => \ppm_encoder_1.N_590_i\
        );

    \I__3999\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20245\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__20245\,
            I => \N__20240\
        );

    \I__3997\ : InMux
    port map (
            O => \N__20244\,
            I => \N__20237\
        );

    \I__3996\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20234\
        );

    \I__3995\ : Span4Mux_s2_v
    port map (
            O => \N__20240\,
            I => \N__20229\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20229\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__20234\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__20229\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__3991\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20221\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__20221\,
            I => \N__20215\
        );

    \I__3989\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20210\
        );

    \I__3988\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20210\
        );

    \I__3987\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20207\
        );

    \I__3986\ : Span4Mux_h
    port map (
            O => \N__20215\,
            I => \N__20204\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__20210\,
            I => \N__20201\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__20207\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__20204\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__20201\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__3981\ : InMux
    port map (
            O => \N__20194\,
            I => \ppm_encoder_1.un1_counter_13_cry_0\
        );

    \I__3980\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20188\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__20185\,
            I => \N__20181\
        );

    \I__3977\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20178\
        );

    \I__3976\ : Span4Mux_h
    port map (
            O => \N__20181\,
            I => \N__20173\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20173\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__20173\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__20170\,
            I => \ppm_encoder_1.N_305_cascade_\
        );

    \I__3972\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20164\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20161\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__20161\,
            I => \N__20158\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__20158\,
            I => \ppm_encoder_1.N_298\
        );

    \I__3968\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20152\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__20152\,
            I => \N__20147\
        );

    \I__3966\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20142\
        );

    \I__3965\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20142\
        );

    \I__3964\ : Odrv12
    port map (
            O => \N__20147\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__20142\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__3962\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20133\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__20136\,
            I => \N__20130\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__20133\,
            I => \N__20126\
        );

    \I__3959\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20123\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__20129\,
            I => \N__20120\
        );

    \I__3957\ : Span4Mux_v
    port map (
            O => \N__20126\,
            I => \N__20117\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__20123\,
            I => \N__20114\
        );

    \I__3955\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20111\
        );

    \I__3954\ : Span4Mux_h
    port map (
            O => \N__20117\,
            I => \N__20108\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__20114\,
            I => \N__20105\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__20111\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__20108\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__20105\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__20098\,
            I => \ppm_encoder_1.N_304_cascade_\
        );

    \I__3948\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20092\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__20092\,
            I => \N__20088\
        );

    \I__3946\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20084\
        );

    \I__3945\ : Span4Mux_s3_h
    port map (
            O => \N__20088\,
            I => \N__20081\
        );

    \I__3944\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20078\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__20084\,
            I => \N__20073\
        );

    \I__3942\ : Span4Mux_h
    port map (
            O => \N__20081\,
            I => \N__20073\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__20078\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__20073\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__3939\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20063\
        );

    \I__3938\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20058\
        );

    \I__3937\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20058\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__20063\,
            I => \N__20055\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__20058\,
            I => \N__20052\
        );

    \I__3934\ : Span4Mux_h
    port map (
            O => \N__20055\,
            I => \N__20049\
        );

    \I__3933\ : Span4Mux_h
    port map (
            O => \N__20052\,
            I => \N__20046\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__20049\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__3931\ : Odrv4
    port map (
            O => \N__20046\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__3930\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20036\
        );

    \I__3929\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20033\
        );

    \I__3928\ : InMux
    port map (
            O => \N__20039\,
            I => \N__20030\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__20036\,
            I => \N__20027\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__20033\,
            I => \N__20024\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__20030\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__20027\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__3923\ : Odrv12
    port map (
            O => \N__20024\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__3921\ : InMux
    port map (
            O => \N__20014\,
            I => \N__20011\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__20011\,
            I => \N__20006\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__20010\,
            I => \N__20001\
        );

    \I__3918\ : InMux
    port map (
            O => \N__20009\,
            I => \N__19998\
        );

    \I__3917\ : Span4Mux_h
    port map (
            O => \N__20006\,
            I => \N__19995\
        );

    \I__3916\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19988\
        );

    \I__3915\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19988\
        );

    \I__3914\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19988\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__19998\,
            I => \N__19985\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__19995\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__19988\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__19985\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__19978\,
            I => \ppm_encoder_1.N_319_cascade_\
        );

    \I__3908\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19972\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19969\
        );

    \I__3906\ : Span4Mux_v
    port map (
            O => \N__19969\,
            I => \N__19966\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__19966\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__19963\,
            I => \N__19959\
        );

    \I__3903\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19956\
        );

    \I__3902\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19953\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__19956\,
            I => \N__19949\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__19953\,
            I => \N__19946\
        );

    \I__3899\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19943\
        );

    \I__3898\ : Span4Mux_v
    port map (
            O => \N__19949\,
            I => \N__19938\
        );

    \I__3897\ : Span4Mux_h
    port map (
            O => \N__19946\,
            I => \N__19938\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__19943\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__19938\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__3894\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19930\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__19930\,
            I => \N__19927\
        );

    \I__3892\ : Span4Mux_s3_v
    port map (
            O => \N__19927\,
            I => \N__19924\
        );

    \I__3891\ : Span4Mux_h
    port map (
            O => \N__19924\,
            I => \N__19921\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__19921\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\
        );

    \I__3889\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19915\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19910\
        );

    \I__3887\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19905\
        );

    \I__3886\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19905\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__19910\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__19905\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__3883\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19897\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19893\
        );

    \I__3881\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19890\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__19893\,
            I => \N__19887\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__19890\,
            I => \N__19884\
        );

    \I__3878\ : Span4Mux_h
    port map (
            O => \N__19887\,
            I => \N__19881\
        );

    \I__3877\ : Odrv12
    port map (
            O => \N__19884\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__19881\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__3875\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19871\
        );

    \I__3874\ : InMux
    port map (
            O => \N__19875\,
            I => \N__19868\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__19874\,
            I => \N__19865\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__19871\,
            I => \N__19862\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__19868\,
            I => \N__19859\
        );

    \I__3870\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19856\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__19862\,
            I => \N__19853\
        );

    \I__3868\ : Span4Mux_h
    port map (
            O => \N__19859\,
            I => \N__19850\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__19856\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__3866\ : Odrv4
    port map (
            O => \N__19853\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__19850\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__3864\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19840\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__19840\,
            I => \N__19837\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__19837\,
            I => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\
        );

    \I__3861\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19831\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__19831\,
            I => \N__19827\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__19830\,
            I => \N__19824\
        );

    \I__3858\ : Span4Mux_s3_v
    port map (
            O => \N__19827\,
            I => \N__19821\
        );

    \I__3857\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19818\
        );

    \I__3856\ : Span4Mux_v
    port map (
            O => \N__19821\,
            I => \N__19812\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__19818\,
            I => \N__19812\
        );

    \I__3854\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19809\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__19812\,
            I => \N__19806\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__19809\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__19806\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3850\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19798\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__19798\,
            I => \N__19793\
        );

    \I__3848\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19790\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__19796\,
            I => \N__19787\
        );

    \I__3846\ : Span4Mux_s3_h
    port map (
            O => \N__19793\,
            I => \N__19784\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19781\
        );

    \I__3844\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19778\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__19784\,
            I => \N__19775\
        );

    \I__3842\ : Span4Mux_h
    port map (
            O => \N__19781\,
            I => \N__19772\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__19778\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3840\ : Odrv4
    port map (
            O => \N__19775\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__19772\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3838\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19762\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__19762\,
            I => \N__19759\
        );

    \I__3836\ : Odrv12
    port map (
            O => \N__19759\,
            I => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\
        );

    \I__3835\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19753\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__19753\,
            I => \N__19750\
        );

    \I__3833\ : Span4Mux_s3_v
    port map (
            O => \N__19750\,
            I => \N__19745\
        );

    \I__3832\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19742\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__19748\,
            I => \N__19739\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__19745\,
            I => \N__19736\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19733\
        );

    \I__3828\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19730\
        );

    \I__3827\ : Span4Mux_v
    port map (
            O => \N__19736\,
            I => \N__19725\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__19733\,
            I => \N__19725\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__19730\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__19725\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__3823\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19717\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19714\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__19714\,
            I => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\
        );

    \I__3820\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19704\
        );

    \I__3819\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19704\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__19709\,
            I => \N__19701\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__19704\,
            I => \N__19698\
        );

    \I__3816\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19695\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__19698\,
            I => \N__19692\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__19695\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__19692\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__3812\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19684\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19681\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__19681\,
            I => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\
        );

    \I__3809\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19675\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19672\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__19672\,
            I => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\
        );

    \I__3806\ : InMux
    port map (
            O => \N__19669\,
            I => \ppm_encoder_1.un1_rudder_cry_7\
        );

    \I__3805\ : InMux
    port map (
            O => \N__19666\,
            I => \ppm_encoder_1.un1_rudder_cry_8\
        );

    \I__3804\ : InMux
    port map (
            O => \N__19663\,
            I => \ppm_encoder_1.un1_rudder_cry_9\
        );

    \I__3803\ : InMux
    port map (
            O => \N__19660\,
            I => \ppm_encoder_1.un1_rudder_cry_10\
        );

    \I__3802\ : InMux
    port map (
            O => \N__19657\,
            I => \ppm_encoder_1.un1_rudder_cry_11\
        );

    \I__3801\ : InMux
    port map (
            O => \N__19654\,
            I => \ppm_encoder_1.un1_rudder_cry_12\
        );

    \I__3800\ : InMux
    port map (
            O => \N__19651\,
            I => \bfn_7_20_0_\
        );

    \I__3799\ : InMux
    port map (
            O => \N__19648\,
            I => \N__19645\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__19645\,
            I => \N__19642\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__19642\,
            I => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\
        );

    \I__3796\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19632\
        );

    \I__3795\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19632\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \N__19629\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19626\
        );

    \I__3792\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19623\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__19626\,
            I => \N__19620\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__19623\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__19620\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__3788\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19610\
        );

    \I__3787\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19607\
        );

    \I__3786\ : CascadeMux
    port map (
            O => \N__19613\,
            I => \N__19604\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19599\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__19607\,
            I => \N__19599\
        );

    \I__3783\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19596\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__19599\,
            I => \N__19593\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__19596\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__19593\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__19588\,
            I => \uart_pc.N_143_cascade_\
        );

    \I__3778\ : SRMux
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__19582\,
            I => \N__19578\
        );

    \I__3776\ : SRMux
    port map (
            O => \N__19581\,
            I => \N__19575\
        );

    \I__3775\ : Span4Mux_h
    port map (
            O => \N__19578\,
            I => \N__19572\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__19575\,
            I => \N__19569\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__19572\,
            I => \N__19566\
        );

    \I__3772\ : Span12Mux_s7_h
    port map (
            O => \N__19569\,
            I => \N__19563\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__19566\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__3770\ : Odrv12
    port map (
            O => \N__19563\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__3769\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19552\
        );

    \I__3768\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19547\
        );

    \I__3767\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19547\
        );

    \I__3766\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19544\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__19552\,
            I => \N__19541\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__19547\,
            I => \N__19536\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19536\
        );

    \I__3762\ : Span4Mux_h
    port map (
            O => \N__19541\,
            I => \N__19531\
        );

    \I__3761\ : Span4Mux_v
    port map (
            O => \N__19536\,
            I => \N__19531\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__19531\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__3759\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__19525\,
            I => \N__19521\
        );

    \I__3757\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19518\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__19521\,
            I => \uart_pc.N_126_li\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__19518\,
            I => \uart_pc.N_126_li\
        );

    \I__3754\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19505\
        );

    \I__3753\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19496\
        );

    \I__3752\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19496\
        );

    \I__3751\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19496\
        );

    \I__3750\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19496\
        );

    \I__3749\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19493\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__19505\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__19496\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__19493\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__3745\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19479\
        );

    \I__3743\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19476\
        );

    \I__3742\ : Span4Mux_v
    port map (
            O => \N__19479\,
            I => \N__19466\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19466\
        );

    \I__3740\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19458\
        );

    \I__3739\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19458\
        );

    \I__3738\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19458\
        );

    \I__3737\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19453\
        );

    \I__3736\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19453\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__19466\,
            I => \N__19450\
        );

    \I__3734\ : InMux
    port map (
            O => \N__19465\,
            I => \N__19447\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__19458\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__19453\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__19450\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__19447\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__19438\,
            I => \uart_pc.N_126_li_cascade_\
        );

    \I__3728\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19425\
        );

    \I__3727\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19410\
        );

    \I__3726\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19410\
        );

    \I__3725\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19410\
        );

    \I__3724\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19410\
        );

    \I__3723\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19410\
        );

    \I__3722\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19410\
        );

    \I__3721\ : InMux
    port map (
            O => \N__19428\,
            I => \N__19410\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__19425\,
            I => \N__19407\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__19410\,
            I => \N__19404\
        );

    \I__3718\ : Span4Mux_h
    port map (
            O => \N__19407\,
            I => \N__19401\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__19404\,
            I => \N__19398\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__19401\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__19398\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__3714\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19390\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__19390\,
            I => \N__19387\
        );

    \I__3712\ : Span4Mux_v
    port map (
            O => \N__19387\,
            I => \N__19384\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__19384\,
            I => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\
        );

    \I__3710\ : InMux
    port map (
            O => \N__19381\,
            I => \ppm_encoder_1.un1_rudder_cry_6\
        );

    \I__3709\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19374\
        );

    \I__3708\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19371\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__19374\,
            I => \N__19367\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__19371\,
            I => \N__19364\
        );

    \I__3705\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19361\
        );

    \I__3704\ : Span4Mux_v
    port map (
            O => \N__19367\,
            I => \N__19358\
        );

    \I__3703\ : Span4Mux_h
    port map (
            O => \N__19364\,
            I => \N__19355\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__19361\,
            I => \uart_pc.N_152\
        );

    \I__3701\ : Odrv4
    port map (
            O => \N__19358\,
            I => \uart_pc.N_152\
        );

    \I__3700\ : Odrv4
    port map (
            O => \N__19355\,
            I => \uart_pc.N_152\
        );

    \I__3699\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19345\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__19345\,
            I => \uart_pc.N_144_1\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__19342\,
            I => \uart_pc.N_144_1_cascade_\
        );

    \I__3696\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19335\
        );

    \I__3695\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19332\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__19335\,
            I => \N__19329\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__19332\,
            I => \N__19324\
        );

    \I__3692\ : Span4Mux_h
    port map (
            O => \N__19329\,
            I => \N__19321\
        );

    \I__3691\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19316\
        );

    \I__3690\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19316\
        );

    \I__3689\ : Span4Mux_h
    port map (
            O => \N__19324\,
            I => \N__19313\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__19321\,
            I => \N__19310\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19307\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__19313\,
            I => \uart_pc.state_1_sqmuxa\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__19310\,
            I => \uart_pc.state_1_sqmuxa\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__19307\,
            I => \uart_pc.state_1_sqmuxa\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__19300\,
            I => \N__19297\
        );

    \I__3682\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19294\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__19294\,
            I => \uart_pc.N_145\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__19291\,
            I => \N__19286\
        );

    \I__3679\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19279\
        );

    \I__3678\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19279\
        );

    \I__3677\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19279\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__19279\,
            I => \N__19275\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__19278\,
            I => \N__19271\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__19275\,
            I => \N__19268\
        );

    \I__3673\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19263\
        );

    \I__3672\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19263\
        );

    \I__3671\ : Sp12to4
    port map (
            O => \N__19268\,
            I => \N__19260\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__19263\,
            I => \N__19257\
        );

    \I__3669\ : Odrv12
    port map (
            O => \N__19260\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__19257\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__19252\,
            I => \N__19246\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__19251\,
            I => \N__19243\
        );

    \I__3665\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19240\
        );

    \I__3664\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19233\
        );

    \I__3663\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19233\
        );

    \I__3662\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19233\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__19240\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__19233\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__3659\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19225\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__19225\,
            I => \N__19222\
        );

    \I__3657\ : Span4Mux_h
    port map (
            O => \N__19222\,
            I => \N__19219\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__19219\,
            I => \uart_drone.data_Auxce_0_6\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__19216\,
            I => \uart_pc.state_srsts_0_0_0_cascade_\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__19213\,
            I => \N__19210\
        );

    \I__3653\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19206\
        );

    \I__3652\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19203\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__19206\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__19203\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__3649\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19195\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__19195\,
            I => \N__19192\
        );

    \I__3647\ : Span4Mux_h
    port map (
            O => \N__19192\,
            I => \N__19188\
        );

    \I__3646\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19185\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__19188\,
            I => \uart_drone.N_126_li\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__19185\,
            I => \uart_drone.N_126_li\
        );

    \I__3643\ : CascadeMux
    port map (
            O => \N__19180\,
            I => \uart_drone.state_srsts_0_0_0_cascade_\
        );

    \I__3642\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19173\
        );

    \I__3641\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19170\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__19173\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__19170\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__3638\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19162\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__19162\,
            I => \N__19159\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__19159\,
            I => \uart_drone.data_Auxce_0_5\
        );

    \I__3635\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19148\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__19155\,
            I => \N__19145\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__19154\,
            I => \N__19142\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__19153\,
            I => \N__19138\
        );

    \I__3631\ : CascadeMux
    port map (
            O => \N__19152\,
            I => \N__19134\
        );

    \I__3630\ : IoInMux
    port map (
            O => \N__19151\,
            I => \N__19129\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19126\
        );

    \I__3628\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19111\
        );

    \I__3627\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19111\
        );

    \I__3626\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19111\
        );

    \I__3625\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19111\
        );

    \I__3624\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19111\
        );

    \I__3623\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19111\
        );

    \I__3622\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19111\
        );

    \I__3621\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19108\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__19129\,
            I => \N__19105\
        );

    \I__3619\ : Span4Mux_v
    port map (
            O => \N__19126\,
            I => \N__19101\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__19111\,
            I => \N__19098\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19095\
        );

    \I__3616\ : IoSpan4Mux
    port map (
            O => \N__19105\,
            I => \N__19089\
        );

    \I__3615\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19086\
        );

    \I__3614\ : Sp12to4
    port map (
            O => \N__19101\,
            I => \N__19083\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__19098\,
            I => \N__19080\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__19095\,
            I => \N__19077\
        );

    \I__3611\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19072\
        );

    \I__3610\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19072\
        );

    \I__3609\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19069\
        );

    \I__3608\ : Span4Mux_s1_v
    port map (
            O => \N__19089\,
            I => \N__19066\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__19086\,
            I => \N__19055\
        );

    \I__3606\ : Span12Mux_h
    port map (
            O => \N__19083\,
            I => \N__19055\
        );

    \I__3605\ : Sp12to4
    port map (
            O => \N__19080\,
            I => \N__19055\
        );

    \I__3604\ : Sp12to4
    port map (
            O => \N__19077\,
            I => \N__19055\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__19072\,
            I => \N__19055\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__19069\,
            I => \N__19052\
        );

    \I__3601\ : Span4Mux_h
    port map (
            O => \N__19066\,
            I => \N__19049\
        );

    \I__3600\ : Span12Mux_v
    port map (
            O => \N__19055\,
            I => \N__19044\
        );

    \I__3599\ : Span12Mux_s7_h
    port map (
            O => \N__19052\,
            I => \N__19044\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__19049\,
            I => uart_commands_input_debug_c
        );

    \I__3597\ : Odrv12
    port map (
            O => \N__19044\,
            I => uart_commands_input_debug_c
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__19039\,
            I => \N__19034\
        );

    \I__3595\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19031\
        );

    \I__3594\ : InMux
    port map (
            O => \N__19037\,
            I => \N__19026\
        );

    \I__3593\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19026\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__19031\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__19026\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__19021\,
            I => \uart_pc.state_srsts_i_0_2_cascade_\
        );

    \I__3589\ : InMux
    port map (
            O => \N__19018\,
            I => \N__19015\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__19015\,
            I => \N__19012\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__19012\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__3586\ : InMux
    port map (
            O => \N__19009\,
            I => \N__19006\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__19006\,
            I => \N__19003\
        );

    \I__3584\ : Span4Mux_h
    port map (
            O => \N__19003\,
            I => \N__19000\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__19000\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__18997\,
            I => \uart_drone.state_srsts_i_0_2_cascade_\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__18994\,
            I => \N__18989\
        );

    \I__3580\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18986\
        );

    \I__3579\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18981\
        );

    \I__3578\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18981\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__18986\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__18981\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__3575\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__18973\,
            I => \N__18970\
        );

    \I__3573\ : Span4Mux_v
    port map (
            O => \N__18970\,
            I => \N__18965\
        );

    \I__3572\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18962\
        );

    \I__3571\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18959\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__18965\,
            I => \N__18955\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__18962\,
            I => \N__18950\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__18959\,
            I => \N__18950\
        );

    \I__3567\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18947\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__18955\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__3565\ : Odrv12
    port map (
            O => \N__18950\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__18947\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__18940\,
            I => \ppm_encoder_1.N_237_cascade_\
        );

    \I__3562\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18932\
        );

    \I__3561\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18929\
        );

    \I__3560\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18925\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18922\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__18929\,
            I => \N__18919\
        );

    \I__3557\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18916\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__18925\,
            I => \N__18913\
        );

    \I__3555\ : Span4Mux_v
    port map (
            O => \N__18922\,
            I => \N__18910\
        );

    \I__3554\ : Span4Mux_s2_v
    port map (
            O => \N__18919\,
            I => \N__18905\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__18916\,
            I => \N__18905\
        );

    \I__3552\ : Span4Mux_v
    port map (
            O => \N__18913\,
            I => \N__18895\
        );

    \I__3551\ : Span4Mux_h
    port map (
            O => \N__18910\,
            I => \N__18895\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__18905\,
            I => \N__18895\
        );

    \I__3549\ : InMux
    port map (
            O => \N__18904\,
            I => \N__18888\
        );

    \I__3548\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18888\
        );

    \I__3547\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18888\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__18895\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__18888\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__3544\ : IoInMux
    port map (
            O => \N__18883\,
            I => \N__18880\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18877\
        );

    \I__3542\ : Span4Mux_s1_v
    port map (
            O => \N__18877\,
            I => \N__18874\
        );

    \I__3541\ : Span4Mux_h
    port map (
            O => \N__18874\,
            I => \N__18871\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__18871\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\
        );

    \I__3539\ : InMux
    port map (
            O => \N__18868\,
            I => \N__18864\
        );

    \I__3538\ : InMux
    port map (
            O => \N__18867\,
            I => \N__18861\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__18864\,
            I => \N__18858\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__18861\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__3535\ : Odrv12
    port map (
            O => \N__18858\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__3534\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18850\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__18850\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\
        );

    \I__3532\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__18844\,
            I => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\
        );

    \I__3530\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18838\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__18838\,
            I => \uart_pc_sync.aux_2__0__0_0\
        );

    \I__3528\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18832\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__18832\,
            I => \uart_pc_sync.aux_3__0__0_0\
        );

    \I__3526\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18826\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__18826\,
            I => \N__18823\
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__18823\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\
        );

    \I__3523\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18817\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__18817\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__18814\,
            I => \N__18811\
        );

    \I__3520\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18808\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__18808\,
            I => \ppm_encoder_1.pulses2countZ0Z_3\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__18805\,
            I => \N__18802\
        );

    \I__3517\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18799\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__18799\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\
        );

    \I__3515\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18793\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__18793\,
            I => \N__18790\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__18790\,
            I => \N__18787\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__18787\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\
        );

    \I__3511\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18781\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__18781\,
            I => \ppm_encoder_1.pulses2countZ0Z_0\
        );

    \I__3509\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__18775\,
            I => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\
        );

    \I__3507\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18769\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__18769\,
            I => \N__18766\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__18766\,
            I => \N__18763\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__18763\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\
        );

    \I__3503\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18757\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__18757\,
            I => \N__18754\
        );

    \I__3501\ : Span4Mux_v
    port map (
            O => \N__18754\,
            I => \N__18751\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__18751\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__18748\,
            I => \N__18745\
        );

    \I__3498\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18742\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__18742\,
            I => \ppm_encoder_1.pulses2countZ0Z_1\
        );

    \I__3496\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18736\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__18736\,
            I => \ppm_encoder_1.pulses2countZ0Z_10\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__18733\,
            I => \N__18730\
        );

    \I__3493\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18727\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__18727\,
            I => \ppm_encoder_1.pulses2countZ0Z_11\
        );

    \I__3491\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18721\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__18721\,
            I => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\
        );

    \I__3489\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18715\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__18715\,
            I => \ppm_encoder_1.pulses2countZ0Z_12\
        );

    \I__3487\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18709\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__18709\,
            I => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\
        );

    \I__3485\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__18703\,
            I => \N__18700\
        );

    \I__3483\ : Odrv12
    port map (
            O => \N__18700\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__18697\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_\
        );

    \I__3481\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18688\
        );

    \I__3480\ : InMux
    port map (
            O => \N__18693\,
            I => \N__18688\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__18688\,
            I => \N__18685\
        );

    \I__3478\ : Span4Mux_h
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__3477\ : Span4Mux_v
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__18679\,
            I => \ppm_encoder_1.N_237\
        );

    \I__3475\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18670\
        );

    \I__3474\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18670\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__18670\,
            I => \N__18667\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__18667\,
            I => \N__18663\
        );

    \I__3471\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18660\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__18663\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__18660\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__3468\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18651\
        );

    \I__3467\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18648\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__18651\,
            I => \N__18643\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__18648\,
            I => \N__18643\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__18640\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__3462\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__18634\,
            I => \N__18631\
        );

    \I__3460\ : Span4Mux_v
    port map (
            O => \N__18631\,
            I => \N__18626\
        );

    \I__3459\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18621\
        );

    \I__3458\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18621\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__18626\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__18621\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__3455\ : InMux
    port map (
            O => \N__18616\,
            I => \N__18613\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__18613\,
            I => \N__18609\
        );

    \I__3453\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18606\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__18609\,
            I => \N__18600\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18600\
        );

    \I__3450\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18597\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__18600\,
            I => \N__18594\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__18597\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__18594\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__3446\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18586\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__18586\,
            I => \N__18583\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__18583\,
            I => \N__18579\
        );

    \I__3443\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18576\
        );

    \I__3442\ : Odrv4
    port map (
            O => \N__18579\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__18576\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__3440\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18567\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__18570\,
            I => \N__18564\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__18567\,
            I => \N__18558\
        );

    \I__3437\ : InMux
    port map (
            O => \N__18564\,
            I => \N__18555\
        );

    \I__3436\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18552\
        );

    \I__3435\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18547\
        );

    \I__3434\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18547\
        );

    \I__3433\ : Span4Mux_h
    port map (
            O => \N__18558\,
            I => \N__18542\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__18555\,
            I => \N__18542\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__18552\,
            I => \N__18539\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18532\
        );

    \I__3429\ : Span4Mux_v
    port map (
            O => \N__18542\,
            I => \N__18532\
        );

    \I__3428\ : Span4Mux_h
    port map (
            O => \N__18539\,
            I => \N__18529\
        );

    \I__3427\ : InMux
    port map (
            O => \N__18538\,
            I => \N__18524\
        );

    \I__3426\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18524\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__18532\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__18529\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__18524\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__18517\,
            I => \ppm_encoder_1.N_296_cascade_\
        );

    \I__3421\ : InMux
    port map (
            O => \N__18514\,
            I => \N__18511\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__18511\,
            I => \N__18508\
        );

    \I__3419\ : Span4Mux_v
    port map (
            O => \N__18508\,
            I => \N__18504\
        );

    \I__3418\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18501\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__18504\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__18501\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__3415\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18493\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__18493\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\
        );

    \I__3413\ : InMux
    port map (
            O => \N__18490\,
            I => \N__18487\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__18487\,
            I => \N__18481\
        );

    \I__3411\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18474\
        );

    \I__3410\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18474\
        );

    \I__3409\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18474\
        );

    \I__3408\ : Odrv12
    port map (
            O => \N__18481\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__18474\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__3406\ : InMux
    port map (
            O => \N__18469\,
            I => \N__18466\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__18466\,
            I => \N__18463\
        );

    \I__3404\ : Span4Mux_h
    port map (
            O => \N__18463\,
            I => \N__18457\
        );

    \I__3403\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18450\
        );

    \I__3402\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18450\
        );

    \I__3401\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18450\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__18457\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__18450\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__3398\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18442\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__18442\,
            I => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\
        );

    \I__3396\ : InMux
    port map (
            O => \N__18439\,
            I => \N__18436\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__18436\,
            I => \N__18433\
        );

    \I__3394\ : Span4Mux_h
    port map (
            O => \N__18433\,
            I => \N__18430\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__18430\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\
        );

    \I__3392\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18424\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18421\
        );

    \I__3390\ : Span4Mux_s3_v
    port map (
            O => \N__18421\,
            I => \N__18418\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__18418\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\
        );

    \I__3388\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18412\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__18412\,
            I => \ppm_encoder_1.pulses2countZ0Z_2\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__18409\,
            I => \N__18406\
        );

    \I__3385\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18397\
        );

    \I__3384\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18397\
        );

    \I__3383\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18397\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__18397\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__3381\ : InMux
    port map (
            O => \N__18394\,
            I => \N__18391\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__18391\,
            I => \N__18388\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__18388\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\
        );

    \I__3378\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18382\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__18382\,
            I => \N__18379\
        );

    \I__3376\ : Span4Mux_h
    port map (
            O => \N__18379\,
            I => \N__18376\
        );

    \I__3375\ : Span4Mux_h
    port map (
            O => \N__18376\,
            I => \N__18373\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__18373\,
            I => \ppm_encoder_1.un1_init_pulses_11_6\
        );

    \I__3373\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18367\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__18367\,
            I => \N__18364\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__18364\,
            I => \ppm_encoder_1.un1_init_pulses_10_6\
        );

    \I__3370\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18358\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__18358\,
            I => \N__18354\
        );

    \I__3368\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18351\
        );

    \I__3367\ : Span4Mux_h
    port map (
            O => \N__18354\,
            I => \N__18348\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__18351\,
            I => \N__18345\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__18348\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__18345\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__3363\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18337\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__18337\,
            I => \N__18334\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__18334\,
            I => \N__18331\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__18331\,
            I => \ppm_encoder_1.un1_init_pulses_11_7\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__18328\,
            I => \N__18325\
        );

    \I__3358\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18322\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__18322\,
            I => \N__18319\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__18319\,
            I => \ppm_encoder_1.un1_init_pulses_10_7\
        );

    \I__3355\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18313\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__18313\,
            I => \N__18310\
        );

    \I__3353\ : Span4Mux_h
    port map (
            O => \N__18310\,
            I => \N__18307\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__18307\,
            I => \ppm_encoder_1.un1_init_pulses_11_14\
        );

    \I__3351\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18301\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__18301\,
            I => \N__18298\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__18298\,
            I => \ppm_encoder_1.un1_init_pulses_10_14\
        );

    \I__3348\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18291\
        );

    \I__3347\ : InMux
    port map (
            O => \N__18294\,
            I => \N__18288\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__18291\,
            I => \N__18285\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__18288\,
            I => \N__18282\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__18285\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__18282\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__3342\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18274\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__18274\,
            I => \N__18271\
        );

    \I__3340\ : Span4Mux_h
    port map (
            O => \N__18271\,
            I => \N__18268\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__18268\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__18265\,
            I => \N__18262\
        );

    \I__3337\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18259\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__18259\,
            I => \N__18256\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__18256\,
            I => \N__18253\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__18253\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_16\
        );

    \I__3333\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18245\
        );

    \I__3332\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18238\
        );

    \I__3331\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18238\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__18245\,
            I => \N__18235\
        );

    \I__3329\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18232\
        );

    \I__3328\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18228\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__18238\,
            I => \N__18224\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__18235\,
            I => \N__18221\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__18232\,
            I => \N__18218\
        );

    \I__3324\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18215\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__18228\,
            I => \N__18212\
        );

    \I__3322\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18206\
        );

    \I__3321\ : Span4Mux_v
    port map (
            O => \N__18224\,
            I => \N__18195\
        );

    \I__3320\ : Span4Mux_h
    port map (
            O => \N__18221\,
            I => \N__18192\
        );

    \I__3319\ : Span4Mux_h
    port map (
            O => \N__18218\,
            I => \N__18187\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__18215\,
            I => \N__18187\
        );

    \I__3317\ : Span4Mux_h
    port map (
            O => \N__18212\,
            I => \N__18184\
        );

    \I__3316\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18177\
        );

    \I__3315\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18177\
        );

    \I__3314\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18177\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__18206\,
            I => \N__18174\
        );

    \I__3312\ : InMux
    port map (
            O => \N__18205\,
            I => \N__18171\
        );

    \I__3311\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18166\
        );

    \I__3310\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18166\
        );

    \I__3309\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18161\
        );

    \I__3308\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18161\
        );

    \I__3307\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18158\
        );

    \I__3306\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18153\
        );

    \I__3305\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18153\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__18195\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__18192\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__18187\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__18184\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__18177\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3299\ : Odrv12
    port map (
            O => \N__18174\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__18171\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__18166\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__18161\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__18158\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__18153\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3293\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18127\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__18127\,
            I => \N__18124\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__18124\,
            I => \N__18121\
        );

    \I__3290\ : Span4Mux_s2_h
    port map (
            O => \N__18121\,
            I => \N__18118\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__18118\,
            I => \ppm_encoder_1.un1_init_pulses_11_4\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__18115\,
            I => \N__18104\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__18114\,
            I => \N__18101\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__18113\,
            I => \N__18098\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__18112\,
            I => \N__18095\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__18111\,
            I => \N__18091\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__18110\,
            I => \N__18087\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__18109\,
            I => \N__18084\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__18108\,
            I => \N__18081\
        );

    \I__3280\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18072\
        );

    \I__3279\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18072\
        );

    \I__3278\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18072\
        );

    \I__3277\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18067\
        );

    \I__3276\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18067\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__18094\,
            I => \N__18064\
        );

    \I__3274\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18055\
        );

    \I__3273\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18055\
        );

    \I__3272\ : InMux
    port map (
            O => \N__18087\,
            I => \N__18055\
        );

    \I__3271\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18050\
        );

    \I__3270\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18050\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__18080\,
            I => \N__18046\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__18079\,
            I => \N__18042\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__18072\,
            I => \N__18039\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__18067\,
            I => \N__18036\
        );

    \I__3265\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18033\
        );

    \I__3264\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18030\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__18062\,
            I => \N__18027\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__18055\,
            I => \N__18023\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__18050\,
            I => \N__18020\
        );

    \I__3260\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18011\
        );

    \I__3259\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18011\
        );

    \I__3258\ : InMux
    port map (
            O => \N__18045\,
            I => \N__18011\
        );

    \I__3257\ : InMux
    port map (
            O => \N__18042\,
            I => \N__18011\
        );

    \I__3256\ : Span4Mux_v
    port map (
            O => \N__18039\,
            I => \N__18001\
        );

    \I__3255\ : Span4Mux_s2_v
    port map (
            O => \N__18036\,
            I => \N__18001\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__18033\,
            I => \N__18001\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__18030\,
            I => \N__18001\
        );

    \I__3252\ : InMux
    port map (
            O => \N__18027\,
            I => \N__17998\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__18026\,
            I => \N__17995\
        );

    \I__3250\ : Span4Mux_v
    port map (
            O => \N__18023\,
            I => \N__17988\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__18020\,
            I => \N__17988\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__18011\,
            I => \N__17988\
        );

    \I__3247\ : InMux
    port map (
            O => \N__18010\,
            I => \N__17985\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__18001\,
            I => \N__17980\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__17998\,
            I => \N__17980\
        );

    \I__3244\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17977\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__17988\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__17985\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__17980\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__17977\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__3239\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__17965\,
            I => \N__17962\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__17962\,
            I => \N__17959\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__17959\,
            I => \ppm_encoder_1.un1_init_pulses_10_4\
        );

    \I__3235\ : InMux
    port map (
            O => \N__17956\,
            I => \N__17953\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__17953\,
            I => \N__17948\
        );

    \I__3233\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17945\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__17951\,
            I => \N__17942\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__17948\,
            I => \N__17938\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__17945\,
            I => \N__17935\
        );

    \I__3229\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17930\
        );

    \I__3228\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17930\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__17938\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__3226\ : Odrv12
    port map (
            O => \N__17935\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__17930\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__3224\ : InMux
    port map (
            O => \N__17923\,
            I => \N__17920\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__17920\,
            I => \N__17915\
        );

    \I__3222\ : InMux
    port map (
            O => \N__17919\,
            I => \N__17912\
        );

    \I__3221\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17909\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__17915\,
            I => \N__17904\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17904\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__17909\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__17904\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__17899\,
            I => \N__17895\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__17898\,
            I => \N__17891\
        );

    \I__3214\ : InMux
    port map (
            O => \N__17895\,
            I => \N__17888\
        );

    \I__3213\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17885\
        );

    \I__3212\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17882\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__17888\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__17885\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__17882\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__17875\,
            I => \ppm_encoder_1.N_302_cascade_\
        );

    \I__3207\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17869\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__17869\,
            I => \N__17866\
        );

    \I__3205\ : Span4Mux_s3_v
    port map (
            O => \N__17866\,
            I => \N__17863\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__17863\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\
        );

    \I__3203\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17852\
        );

    \I__3202\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17852\
        );

    \I__3201\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17847\
        );

    \I__3200\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17847\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__17852\,
            I => \N__17844\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17839\
        );

    \I__3197\ : Span4Mux_h
    port map (
            O => \N__17844\,
            I => \N__17836\
        );

    \I__3196\ : InMux
    port map (
            O => \N__17843\,
            I => \N__17831\
        );

    \I__3195\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17831\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__17839\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__17836\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__17831\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__17824\,
            I => \N__17820\
        );

    \I__3190\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17815\
        );

    \I__3189\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17810\
        );

    \I__3188\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17810\
        );

    \I__3187\ : InMux
    port map (
            O => \N__17818\,
            I => \N__17805\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__17815\,
            I => \N__17802\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__17810\,
            I => \N__17798\
        );

    \I__3184\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17793\
        );

    \I__3183\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17793\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__17805\,
            I => \N__17788\
        );

    \I__3181\ : Span4Mux_v
    port map (
            O => \N__17802\,
            I => \N__17788\
        );

    \I__3180\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17785\
        );

    \I__3179\ : Span4Mux_h
    port map (
            O => \N__17798\,
            I => \N__17780\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__17793\,
            I => \N__17780\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__17788\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__17785\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__17780\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3174\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17770\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__17770\,
            I => \N__17767\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__17767\,
            I => \N__17764\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__17764\,
            I => \ppm_encoder_1.un1_init_pulses_11_5\
        );

    \I__3170\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17758\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17755\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__17755\,
            I => \ppm_encoder_1.un1_init_pulses_10_5\
        );

    \I__3167\ : InMux
    port map (
            O => \N__17752\,
            I => \N__17749\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__17749\,
            I => \N__17746\
        );

    \I__3165\ : Span4Mux_v
    port map (
            O => \N__17746\,
            I => \N__17742\
        );

    \I__3164\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17739\
        );

    \I__3163\ : Sp12to4
    port map (
            O => \N__17742\,
            I => \N__17734\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__17739\,
            I => \N__17734\
        );

    \I__3161\ : Odrv12
    port map (
            O => \N__17734\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__3160\ : InMux
    port map (
            O => \N__17731\,
            I => \N__17728\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17725\
        );

    \I__3158\ : Span4Mux_h
    port map (
            O => \N__17725\,
            I => \N__17722\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__17722\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_5\
        );

    \I__3156\ : InMux
    port map (
            O => \N__17719\,
            I => \N__17716\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__17716\,
            I => \N__17712\
        );

    \I__3154\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17709\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__17712\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__17709\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__3151\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17701\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__17701\,
            I => \uart_pc.data_Auxce_0_3\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__17698\,
            I => \N__17695\
        );

    \I__3148\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17692\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17689\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__17689\,
            I => \N__17685\
        );

    \I__3145\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17682\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__17685\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__17682\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__3142\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17674\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__17674\,
            I => \uart_pc.data_Auxce_0_0_4\
        );

    \I__3140\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17667\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__17670\,
            I => \N__17664\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__17667\,
            I => \N__17661\
        );

    \I__3137\ : InMux
    port map (
            O => \N__17664\,
            I => \N__17658\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__17661\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__17658\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__3134\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17650\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__17650\,
            I => \uart_pc.data_Auxce_0_5\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__17647\,
            I => \N__17644\
        );

    \I__3131\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17641\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__17641\,
            I => \N__17638\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__17638\,
            I => \N__17634\
        );

    \I__3128\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17631\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__17634\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__17631\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__17626\,
            I => \N__17623\
        );

    \I__3124\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17620\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__3122\ : Span4Mux_h
    port map (
            O => \N__17617\,
            I => \N__17613\
        );

    \I__3121\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17610\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__17613\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__17610\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__3118\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17602\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__17602\,
            I => \N__17599\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__17599\,
            I => \N__17596\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__17596\,
            I => \uart_pc.data_Auxce_0_6\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__17593\,
            I => \N__17590\
        );

    \I__3113\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17587\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__17587\,
            I => \N__17583\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__17586\,
            I => \N__17580\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__17583\,
            I => \N__17577\
        );

    \I__3109\ : InMux
    port map (
            O => \N__17580\,
            I => \N__17574\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__17577\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__17574\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__17569\,
            I => \N__17566\
        );

    \I__3105\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17562\
        );

    \I__3104\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17559\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__17562\,
            I => \N__17556\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__17559\,
            I => \N__17553\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__17556\,
            I => \N__17549\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__17553\,
            I => \N__17546\
        );

    \I__3099\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17543\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__17549\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__17546\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__17543\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__3095\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17532\
        );

    \I__3094\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17529\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__17532\,
            I => \N__17526\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__17529\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__17526\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__17521\,
            I => \N__17517\
        );

    \I__3089\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17510\
        );

    \I__3088\ : InMux
    port map (
            O => \N__17517\,
            I => \N__17510\
        );

    \I__3087\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17505\
        );

    \I__3086\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17505\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17502\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__17505\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__17502\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__17497\,
            I => \N__17494\
        );

    \I__3081\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17491\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__17491\,
            I => \N__17488\
        );

    \I__3079\ : Odrv4
    port map (
            O => \N__17488\,
            I => \uart_drone.un1_state_2_0_a3_0\
        );

    \I__3078\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17480\
        );

    \I__3077\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17475\
        );

    \I__3076\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17475\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__17480\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__17475\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__3073\ : InMux
    port map (
            O => \N__17470\,
            I => \N__17467\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__17467\,
            I => \uart_drone.timer_Count_RNO_0_0_2\
        );

    \I__3071\ : InMux
    port map (
            O => \N__17464\,
            I => \uart_drone.un4_timer_Count_1_cry_1\
        );

    \I__3070\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17458\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__17458\,
            I => \uart_drone.timer_Count_RNO_0_0_3\
        );

    \I__3068\ : InMux
    port map (
            O => \N__17455\,
            I => \uart_drone.un4_timer_Count_1_cry_2\
        );

    \I__3067\ : InMux
    port map (
            O => \N__17452\,
            I => \uart_drone.un4_timer_Count_1_cry_3\
        );

    \I__3066\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17446\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__17446\,
            I => \uart_drone.timer_Count_RNO_0_0_4\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__17443\,
            I => \N__17440\
        );

    \I__3063\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17433\
        );

    \I__3062\ : InMux
    port map (
            O => \N__17439\,
            I => \N__17433\
        );

    \I__3061\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17429\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__17433\,
            I => \N__17426\
        );

    \I__3059\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17423\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__17429\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__17426\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__17423\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__3055\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17412\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__17415\,
            I => \N__17409\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__17412\,
            I => \N__17406\
        );

    \I__3052\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17403\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__17406\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__17403\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__3049\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17394\
        );

    \I__3048\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17391\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__17394\,
            I => \N__17381\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__17391\,
            I => \N__17381\
        );

    \I__3045\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17372\
        );

    \I__3044\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17372\
        );

    \I__3043\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17372\
        );

    \I__3042\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17372\
        );

    \I__3041\ : InMux
    port map (
            O => \N__17386\,
            I => \N__17367\
        );

    \I__3040\ : Span4Mux_v
    port map (
            O => \N__17381\,
            I => \N__17362\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17362\
        );

    \I__3038\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17357\
        );

    \I__3037\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17357\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__17367\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__17362\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__17357\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__3033\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17345\
        );

    \I__3032\ : InMux
    port map (
            O => \N__17349\,
            I => \N__17342\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__17348\,
            I => \N__17336\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__17345\,
            I => \N__17333\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__17342\,
            I => \N__17330\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__17341\,
            I => \N__17327\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__17340\,
            I => \N__17323\
        );

    \I__3026\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17315\
        );

    \I__3025\ : InMux
    port map (
            O => \N__17336\,
            I => \N__17315\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__17333\,
            I => \N__17312\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__17330\,
            I => \N__17309\
        );

    \I__3022\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17300\
        );

    \I__3021\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17300\
        );

    \I__3020\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17300\
        );

    \I__3019\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17300\
        );

    \I__3018\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17295\
        );

    \I__3017\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17295\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__17315\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__17312\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__17309\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__17300\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__17295\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__3011\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17274\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__17283\,
            I => \N__17270\
        );

    \I__3009\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17265\
        );

    \I__3008\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17265\
        );

    \I__3007\ : InMux
    port map (
            O => \N__17280\,
            I => \N__17256\
        );

    \I__3006\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17256\
        );

    \I__3005\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17256\
        );

    \I__3004\ : InMux
    port map (
            O => \N__17277\,
            I => \N__17256\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__17274\,
            I => \N__17253\
        );

    \I__3002\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17250\
        );

    \I__3001\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17245\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__17265\,
            I => \N__17240\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__17256\,
            I => \N__17240\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__17253\,
            I => \N__17235\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__17250\,
            I => \N__17235\
        );

    \I__2996\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17230\
        );

    \I__2995\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17230\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__17245\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__17240\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__17235\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__17230\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__2990\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17218\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__17218\,
            I => \N__17215\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__17215\,
            I => \uart_pc.data_Auxce_0_0_0\
        );

    \I__2987\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17208\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__17211\,
            I => \N__17205\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__17208\,
            I => \N__17202\
        );

    \I__2984\ : InMux
    port map (
            O => \N__17205\,
            I => \N__17199\
        );

    \I__2983\ : Odrv12
    port map (
            O => \N__17202\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__17199\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__2981\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17191\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__17191\,
            I => \uart_pc.data_Auxce_0_1\
        );

    \I__2979\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17185\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__17185\,
            I => \N__17182\
        );

    \I__2977\ : Span4Mux_h
    port map (
            O => \N__17182\,
            I => \N__17178\
        );

    \I__2976\ : InMux
    port map (
            O => \N__17181\,
            I => \N__17175\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__17178\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__17175\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__2973\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17167\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__17167\,
            I => \N__17164\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__17164\,
            I => \N__17161\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__17161\,
            I => \uart_pc.data_Auxce_0_0_2\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__17158\,
            I => \N__17155\
        );

    \I__2968\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17151\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__17154\,
            I => \N__17148\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__17151\,
            I => \N__17145\
        );

    \I__2965\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17142\
        );

    \I__2964\ : Odrv12
    port map (
            O => \N__17145\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__17142\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__2962\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17132\
        );

    \I__2961\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17127\
        );

    \I__2960\ : InMux
    port map (
            O => \N__17135\,
            I => \N__17127\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__17132\,
            I => \N__17124\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__17127\,
            I => \N__17121\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__17124\,
            I => \uart_drone.state_1_sqmuxa\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__17121\,
            I => \uart_drone.state_1_sqmuxa\
        );

    \I__2955\ : SRMux
    port map (
            O => \N__17116\,
            I => \N__17113\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__17113\,
            I => \N__17109\
        );

    \I__2953\ : SRMux
    port map (
            O => \N__17112\,
            I => \N__17106\
        );

    \I__2952\ : Sp12to4
    port map (
            O => \N__17109\,
            I => \N__17103\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__2950\ : Odrv12
    port map (
            O => \N__17103\,
            I => \Commands_frame_decoder.un1_state49_iZ0\
        );

    \I__2949\ : Odrv12
    port map (
            O => \N__17100\,
            I => \Commands_frame_decoder.un1_state49_iZ0\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__17095\,
            I => \uart_drone.N_126_li_cascade_\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__17092\,
            I => \uart_drone.N_143_cascade_\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__17089\,
            I => \N__17085\
        );

    \I__2945\ : InMux
    port map (
            O => \N__17088\,
            I => \N__17082\
        );

    \I__2944\ : InMux
    port map (
            O => \N__17085\,
            I => \N__17079\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__17082\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__17079\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__17074\,
            I => \N__17070\
        );

    \I__2940\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17067\
        );

    \I__2939\ : InMux
    port map (
            O => \N__17070\,
            I => \N__17064\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__17067\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__17064\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__17059\,
            I => \N__17055\
        );

    \I__2935\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17052\
        );

    \I__2934\ : InMux
    port map (
            O => \N__17055\,
            I => \N__17049\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__17052\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__17049\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__17044\,
            I => \uart_drone.timer_Count_RNO_0_0_1_cascade_\
        );

    \I__2930\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17038\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__17038\,
            I => \N__17033\
        );

    \I__2928\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17030\
        );

    \I__2927\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17027\
        );

    \I__2926\ : Span4Mux_h
    port map (
            O => \N__17033\,
            I => \N__17019\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__17030\,
            I => \N__17019\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__17027\,
            I => \N__17016\
        );

    \I__2923\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17011\
        );

    \I__2922\ : InMux
    port map (
            O => \N__17025\,
            I => \N__17011\
        );

    \I__2921\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17008\
        );

    \I__2920\ : Odrv4
    port map (
            O => \N__17019\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__17016\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__17011\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__17008\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__2916\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16996\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16988\
        );

    \I__2914\ : InMux
    port map (
            O => \N__16995\,
            I => \N__16982\
        );

    \I__2913\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16982\
        );

    \I__2912\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16975\
        );

    \I__2911\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16975\
        );

    \I__2910\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16975\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__16988\,
            I => \N__16972\
        );

    \I__2908\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16968\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__16982\,
            I => \N__16963\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__16975\,
            I => \N__16963\
        );

    \I__2905\ : Span4Mux_h
    port map (
            O => \N__16972\,
            I => \N__16960\
        );

    \I__2904\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16957\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__16968\,
            I => \N__16952\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__16963\,
            I => \N__16952\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__16960\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__16957\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__16952\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__2898\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__2897\ : InMux
    port map (
            O => \N__16944\,
            I => \N__16939\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__16939\,
            I => \Commands_frame_decoder.state_1Z0Z_5\
        );

    \I__2895\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16933\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__16933\,
            I => \N__16930\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__16930\,
            I => \Commands_frame_decoder.state_1_ns_i_a2_3_1Z0Z_0\
        );

    \I__2892\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16924\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__16924\,
            I => \Commands_frame_decoder.state_1_ns_0_a4_0_3_2\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__16921\,
            I => \Commands_frame_decoder.N_323_cascade_\
        );

    \I__2889\ : CEMux
    port map (
            O => \N__16918\,
            I => \N__16915\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__16915\,
            I => \N__16912\
        );

    \I__2887\ : Span4Mux_h
    port map (
            O => \N__16912\,
            I => \N__16909\
        );

    \I__2886\ : Odrv4
    port map (
            O => \N__16909\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\
        );

    \I__2885\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16902\
        );

    \I__2884\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16899\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__16902\,
            I => \Commands_frame_decoder.state_1Z0Z_2\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__16899\,
            I => \Commands_frame_decoder.state_1Z0Z_2\
        );

    \I__2881\ : InMux
    port map (
            O => \N__16894\,
            I => \N__16882\
        );

    \I__2880\ : InMux
    port map (
            O => \N__16893\,
            I => \N__16882\
        );

    \I__2879\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16882\
        );

    \I__2878\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16882\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__16882\,
            I => \N__16879\
        );

    \I__2876\ : Span4Mux_h
    port map (
            O => \N__16879\,
            I => \N__16875\
        );

    \I__2875\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16872\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__16875\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__16872\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__16867\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\
        );

    \I__2871\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16858\
        );

    \I__2870\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16858\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__16858\,
            I => \Commands_frame_decoder.state_1Z0Z_3\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__16855\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_\
        );

    \I__2867\ : InMux
    port map (
            O => \N__16852\,
            I => \N__16848\
        );

    \I__2866\ : InMux
    port map (
            O => \N__16851\,
            I => \N__16845\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__16848\,
            I => \N__16842\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__16845\,
            I => \Commands_frame_decoder.state_1Z0Z_4\
        );

    \I__2863\ : Odrv12
    port map (
            O => \N__16842\,
            I => \Commands_frame_decoder.state_1Z0Z_4\
        );

    \I__2862\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16833\
        );

    \I__2861\ : InMux
    port map (
            O => \N__16836\,
            I => \N__16830\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__16833\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__16830\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__2858\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16821\
        );

    \I__2857\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16818\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__16821\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__16818\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__16813\,
            I => \N__16810\
        );

    \I__2853\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16806\
        );

    \I__2852\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16803\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__16806\,
            I => \N__16800\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__16803\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__16800\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__2848\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16791\
        );

    \I__2847\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16788\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__16791\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__16788\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__16783\,
            I => \N__16778\
        );

    \I__2843\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16774\
        );

    \I__2842\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16771\
        );

    \I__2841\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16766\
        );

    \I__2840\ : InMux
    port map (
            O => \N__16777\,
            I => \N__16766\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__16774\,
            I => \N__16761\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__16771\,
            I => \N__16761\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__16766\,
            I => \reset_module_System.reset6_15\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__16761\,
            I => \reset_module_System.reset6_15\
        );

    \I__2835\ : InMux
    port map (
            O => \N__16756\,
            I => \N__16753\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__16753\,
            I => \N__16749\
        );

    \I__2833\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16746\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__16749\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__16746\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__2830\ : InMux
    port map (
            O => \N__16741\,
            I => \N__16737\
        );

    \I__2829\ : InMux
    port map (
            O => \N__16740\,
            I => \N__16734\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__16737\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__16734\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__16729\,
            I => \N__16726\
        );

    \I__2825\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16722\
        );

    \I__2824\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16719\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__16722\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__16719\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__2821\ : InMux
    port map (
            O => \N__16714\,
            I => \N__16710\
        );

    \I__2820\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16707\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__16710\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__16707\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__2817\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16696\
        );

    \I__2816\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16691\
        );

    \I__2815\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16691\
        );

    \I__2814\ : InMux
    port map (
            O => \N__16699\,
            I => \N__16688\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__16696\,
            I => \N__16681\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__16691\,
            I => \N__16681\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__16688\,
            I => \N__16681\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__16681\,
            I => \reset_module_System.reset6_14\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__16678\,
            I => \N__16673\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__16677\,
            I => \N__16669\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__16676\,
            I => \N__16666\
        );

    \I__2806\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16654\
        );

    \I__2805\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16654\
        );

    \I__2804\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16654\
        );

    \I__2803\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16654\
        );

    \I__2802\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16651\
        );

    \I__2801\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16646\
        );

    \I__2800\ : InMux
    port map (
            O => \N__16663\,
            I => \N__16646\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__16654\,
            I => \N__16639\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__16651\,
            I => \N__16639\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__16646\,
            I => \N__16639\
        );

    \I__2796\ : Span4Mux_v
    port map (
            O => \N__16639\,
            I => \N__16636\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__16636\,
            I => \Commands_frame_decoder.state_1_RNIVM1OZ0Z_6\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__16633\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\
        );

    \I__2793\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16627\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__16627\,
            I => \N__16624\
        );

    \I__2791\ : Span4Mux_v
    port map (
            O => \N__16624\,
            I => \N__16620\
        );

    \I__2790\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16617\
        );

    \I__2789\ : Span4Mux_h
    port map (
            O => \N__16620\,
            I => \N__16614\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__16617\,
            I => alt_kp_4
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__16614\,
            I => alt_kp_4
        );

    \I__2786\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16606\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__16606\,
            I => \N__16603\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__16603\,
            I => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\
        );

    \I__2783\ : InMux
    port map (
            O => \N__16600\,
            I => \ppm_encoder_1.counter24_0_N_2\
        );

    \I__2782\ : InMux
    port map (
            O => \N__16597\,
            I => \N__16592\
        );

    \I__2781\ : InMux
    port map (
            O => \N__16596\,
            I => \N__16589\
        );

    \I__2780\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16586\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__16592\,
            I => \reset_module_System.reset6_19\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__16589\,
            I => \reset_module_System.reset6_19\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__16586\,
            I => \reset_module_System.reset6_19\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__16579\,
            I => \N__16576\
        );

    \I__2775\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16573\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__16573\,
            I => \N__16570\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__16570\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\
        );

    \I__2772\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16564\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__16564\,
            I => \N__16561\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__16561\,
            I => \N__16558\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__16558\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\
        );

    \I__2768\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16552\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__16552\,
            I => \ppm_encoder_1.pulses2countZ0Z_4\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__16549\,
            I => \N__16546\
        );

    \I__2765\ : InMux
    port map (
            O => \N__16546\,
            I => \N__16543\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__16543\,
            I => \ppm_encoder_1.pulses2countZ0Z_5\
        );

    \I__2763\ : InMux
    port map (
            O => \N__16540\,
            I => \N__16537\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__16537\,
            I => \N__16534\
        );

    \I__2761\ : Odrv12
    port map (
            O => \N__16534\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\
        );

    \I__2760\ : InMux
    port map (
            O => \N__16531\,
            I => \N__16528\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__16528\,
            I => \N__16525\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__16525\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\
        );

    \I__2757\ : InMux
    port map (
            O => \N__16522\,
            I => \N__16519\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__16519\,
            I => \N__16516\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__16516\,
            I => \N__16513\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__16513\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\
        );

    \I__2753\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16507\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__16507\,
            I => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\
        );

    \I__2751\ : InMux
    port map (
            O => \N__16504\,
            I => \N__16501\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__16501\,
            I => \N__16498\
        );

    \I__2749\ : Span4Mux_v
    port map (
            O => \N__16498\,
            I => \N__16495\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__16495\,
            I => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__16492\,
            I => \N__16489\
        );

    \I__2746\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16486\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16483\
        );

    \I__2744\ : Span4Mux_h
    port map (
            O => \N__16483\,
            I => \N__16480\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__16480\,
            I => \ppm_encoder_1.un1_init_pulses_11_15\
        );

    \I__2742\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16474\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__16474\,
            I => \ppm_encoder_1.un1_init_pulses_10_15\
        );

    \I__2740\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16468\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__16468\,
            I => \N__16465\
        );

    \I__2738\ : Span4Mux_s3_v
    port map (
            O => \N__16465\,
            I => \N__16462\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__16462\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_15\
        );

    \I__2736\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16452\
        );

    \I__2735\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16452\
        );

    \I__2734\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16449\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__16452\,
            I => \N__16444\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__16449\,
            I => \N__16437\
        );

    \I__2731\ : InMux
    port map (
            O => \N__16448\,
            I => \N__16432\
        );

    \I__2730\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16432\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__16444\,
            I => \N__16429\
        );

    \I__2728\ : InMux
    port map (
            O => \N__16443\,
            I => \N__16426\
        );

    \I__2727\ : InMux
    port map (
            O => \N__16442\,
            I => \N__16419\
        );

    \I__2726\ : InMux
    port map (
            O => \N__16441\,
            I => \N__16419\
        );

    \I__2725\ : InMux
    port map (
            O => \N__16440\,
            I => \N__16419\
        );

    \I__2724\ : Span4Mux_s3_v
    port map (
            O => \N__16437\,
            I => \N__16414\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__16432\,
            I => \N__16414\
        );

    \I__2722\ : Odrv4
    port map (
            O => \N__16429\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__16426\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__16419\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__16414\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__2718\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16402\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__16402\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_18\
        );

    \I__2716\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16396\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__16396\,
            I => \N__16393\
        );

    \I__2714\ : Span4Mux_h
    port map (
            O => \N__16393\,
            I => \N__16390\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__16390\,
            I => \ppm_encoder_1.un1_init_pulses_11_18\
        );

    \I__2712\ : InMux
    port map (
            O => \N__16387\,
            I => \N__16384\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__16384\,
            I => \ppm_encoder_1.un1_init_pulses_10_18\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__16381\,
            I => \N__16378\
        );

    \I__2709\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16375\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__16375\,
            I => \N__16372\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__16372\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\
        );

    \I__2706\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16366\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__16366\,
            I => \N__16363\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__16363\,
            I => \N__16360\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__16360\,
            I => \ppm_encoder_1.un1_init_pulses_11_13\
        );

    \I__2702\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16354\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__16354\,
            I => \ppm_encoder_1.un1_init_pulses_10_13\
        );

    \I__2700\ : InMux
    port map (
            O => \N__16351\,
            I => \N__16348\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__16348\,
            I => \N__16345\
        );

    \I__2698\ : Span4Mux_h
    port map (
            O => \N__16345\,
            I => \N__16341\
        );

    \I__2697\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16338\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__16341\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__16338\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__16333\,
            I => \N__16330\
        );

    \I__2693\ : InMux
    port map (
            O => \N__16330\,
            I => \N__16327\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__16327\,
            I => \N__16323\
        );

    \I__2691\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16320\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__16323\,
            I => \N__16314\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__16320\,
            I => \N__16314\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__16319\,
            I => \N__16308\
        );

    \I__2687\ : Span4Mux_h
    port map (
            O => \N__16314\,
            I => \N__16305\
        );

    \I__2686\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16302\
        );

    \I__2685\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16295\
        );

    \I__2684\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16295\
        );

    \I__2683\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16295\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__16305\,
            I => \ppm_encoder_1.N_226\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__16302\,
            I => \ppm_encoder_1.N_226\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__16295\,
            I => \ppm_encoder_1.N_226\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__16288\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\
        );

    \I__2678\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16282\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__16282\,
            I => \ppm_encoder_1.un1_init_pulses_10_1\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__16279\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_\
        );

    \I__2675\ : InMux
    port map (
            O => \N__16276\,
            I => \N__16273\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__16273\,
            I => \N__16270\
        );

    \I__2673\ : Span4Mux_h
    port map (
            O => \N__16270\,
            I => \N__16267\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__16267\,
            I => \ppm_encoder_1.un1_init_pulses_11_1\
        );

    \I__2671\ : InMux
    port map (
            O => \N__16264\,
            I => \N__16261\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__16261\,
            I => \N__16257\
        );

    \I__2669\ : InMux
    port map (
            O => \N__16260\,
            I => \N__16254\
        );

    \I__2668\ : Span4Mux_v
    port map (
            O => \N__16257\,
            I => \N__16251\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__16251\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__16248\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__2664\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16240\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__16240\,
            I => \N__16235\
        );

    \I__2662\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16230\
        );

    \I__2661\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16230\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__16235\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__16230\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__2658\ : InMux
    port map (
            O => \N__16225\,
            I => \N__16222\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__16222\,
            I => \N__16219\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__16216\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_1\
        );

    \I__2654\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16207\
        );

    \I__2652\ : Span4Mux_h
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__16204\,
            I => \ppm_encoder_1.un1_init_pulses_11_10\
        );

    \I__2650\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16198\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__16198\,
            I => \ppm_encoder_1.un1_init_pulses_10_10\
        );

    \I__2648\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16188\
        );

    \I__2647\ : InMux
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__16193\,
            I => \N__16185\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__16188\,
            I => \N__16182\
        );

    \I__2644\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16179\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__16182\,
            I => \N__16176\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__16179\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__16176\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__16171\,
            I => \N__16168\
        );

    \I__2639\ : InMux
    port map (
            O => \N__16168\,
            I => \N__16165\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__16165\,
            I => \N__16162\
        );

    \I__2637\ : Span4Mux_h
    port map (
            O => \N__16162\,
            I => \N__16159\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__16159\,
            I => \ppm_encoder_1.un1_init_pulses_11_11\
        );

    \I__2635\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16153\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__16153\,
            I => \ppm_encoder_1.un1_init_pulses_10_11\
        );

    \I__2633\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16145\
        );

    \I__2632\ : InMux
    port map (
            O => \N__16149\,
            I => \N__16142\
        );

    \I__2631\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16139\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__16145\,
            I => \N__16136\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__16142\,
            I => \N__16133\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__16139\,
            I => \N__16128\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__16136\,
            I => \N__16128\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__16133\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__16128\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__2624\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16120\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16120\,
            I => \N__16117\
        );

    \I__2622\ : Span4Mux_v
    port map (
            O => \N__16117\,
            I => \N__16114\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__16114\,
            I => \ppm_encoder_1.un1_init_pulses_11_12\
        );

    \I__2620\ : InMux
    port map (
            O => \N__16111\,
            I => \N__16108\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__16108\,
            I => \ppm_encoder_1.un1_init_pulses_10_12\
        );

    \I__2618\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16101\
        );

    \I__2617\ : InMux
    port map (
            O => \N__16104\,
            I => \N__16098\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__16101\,
            I => \N__16095\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16092\
        );

    \I__2614\ : Span4Mux_v
    port map (
            O => \N__16095\,
            I => \N__16089\
        );

    \I__2613\ : Span4Mux_h
    port map (
            O => \N__16092\,
            I => \N__16086\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__16089\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__16086\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__16081\,
            I => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__16078\,
            I => \N__16075\
        );

    \I__2608\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16072\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__16072\,
            I => \N__16069\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__16069\,
            I => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__16066\,
            I => \N__16062\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__16065\,
            I => \N__16057\
        );

    \I__2603\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16047\
        );

    \I__2602\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16047\
        );

    \I__2601\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16047\
        );

    \I__2600\ : InMux
    port map (
            O => \N__16057\,
            I => \N__16044\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__16056\,
            I => \N__16038\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__16055\,
            I => \N__16035\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \N__16032\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__16047\,
            I => \N__16028\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__16044\,
            I => \N__16025\
        );

    \I__2594\ : InMux
    port map (
            O => \N__16043\,
            I => \N__16020\
        );

    \I__2593\ : InMux
    port map (
            O => \N__16042\,
            I => \N__16020\
        );

    \I__2592\ : InMux
    port map (
            O => \N__16041\,
            I => \N__16015\
        );

    \I__2591\ : InMux
    port map (
            O => \N__16038\,
            I => \N__16015\
        );

    \I__2590\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16012\
        );

    \I__2589\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16007\
        );

    \I__2588\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16007\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__16028\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__16025\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__16020\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__16015\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__16012\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__16007\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__2581\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15981\
        );

    \I__2580\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15981\
        );

    \I__2579\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15981\
        );

    \I__2578\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15978\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__15990\,
            I => \N__15974\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__15989\,
            I => \N__15971\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__15988\,
            I => \N__15966\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__15981\,
            I => \N__15961\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__15978\,
            I => \N__15958\
        );

    \I__2572\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15955\
        );

    \I__2571\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15950\
        );

    \I__2570\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15950\
        );

    \I__2569\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15947\
        );

    \I__2568\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15942\
        );

    \I__2567\ : InMux
    port map (
            O => \N__15966\,
            I => \N__15942\
        );

    \I__2566\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15937\
        );

    \I__2565\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15937\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__15961\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__15958\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__15955\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__15950\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__15947\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__15942\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__15937\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__2557\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15919\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__15919\,
            I => \ppm_encoder_1.un2_throttle_iv_1_11\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__15916\,
            I => \N__15913\
        );

    \I__2554\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15910\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__15910\,
            I => \N__15906\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__15909\,
            I => \N__15903\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__15906\,
            I => \N__15898\
        );

    \I__2550\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15895\
        );

    \I__2549\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15890\
        );

    \I__2548\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15890\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__15898\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__15895\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__15890\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__15883\,
            I => \N__15878\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__15882\,
            I => \N__15875\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__15881\,
            I => \N__15872\
        );

    \I__2541\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15869\
        );

    \I__2540\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15866\
        );

    \I__2539\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15859\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__15869\,
            I => \N__15856\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15853\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__15865\,
            I => \N__15841\
        );

    \I__2535\ : InMux
    port map (
            O => \N__15864\,
            I => \N__15838\
        );

    \I__2534\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15833\
        );

    \I__2533\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15833\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__15859\,
            I => \N__15830\
        );

    \I__2531\ : Span4Mux_h
    port map (
            O => \N__15856\,
            I => \N__15825\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__15853\,
            I => \N__15825\
        );

    \I__2529\ : InMux
    port map (
            O => \N__15852\,
            I => \N__15818\
        );

    \I__2528\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15818\
        );

    \I__2527\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15818\
        );

    \I__2526\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15815\
        );

    \I__2525\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15812\
        );

    \I__2524\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15809\
        );

    \I__2523\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15806\
        );

    \I__2522\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15801\
        );

    \I__2521\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15801\
        );

    \I__2520\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15798\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__15838\,
            I => \N__15793\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__15833\,
            I => \N__15793\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__15830\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__15825\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__15818\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__15815\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__15812\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__15809\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__15806\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__15801\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__15798\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__15793\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__15772\,
            I => \N__15766\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__15771\,
            I => \N__15762\
        );

    \I__2505\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15758\
        );

    \I__2504\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15754\
        );

    \I__2503\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15747\
        );

    \I__2502\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15747\
        );

    \I__2501\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15747\
        );

    \I__2500\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15742\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__15758\,
            I => \N__15739\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__15757\,
            I => \N__15736\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__15754\,
            I => \N__15733\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__15747\,
            I => \N__15730\
        );

    \I__2495\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15727\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__15745\,
            I => \N__15723\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__15742\,
            I => \N__15720\
        );

    \I__2492\ : Span4Mux_h
    port map (
            O => \N__15739\,
            I => \N__15717\
        );

    \I__2491\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15714\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__15733\,
            I => \N__15709\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__15730\,
            I => \N__15709\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__15727\,
            I => \N__15706\
        );

    \I__2487\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15701\
        );

    \I__2486\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15701\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__15720\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__15717\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__15714\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__15709\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__15706\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__15701\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__2479\ : InMux
    port map (
            O => \N__15688\,
            I => \N__15684\
        );

    \I__2478\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15681\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__15684\,
            I => \N__15676\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__15681\,
            I => \N__15676\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__15676\,
            I => \N__15673\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__15673\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__15670\,
            I => \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\
        );

    \I__2472\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15664\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__15664\,
            I => \ppm_encoder_1.un2_throttle_iv_1_10\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__15661\,
            I => \N__15658\
        );

    \I__2469\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15655\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__15655\,
            I => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\
        );

    \I__2467\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15649\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__15649\,
            I => \ppm_encoder_1.N_318\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__15646\,
            I => \ppm_encoder_1.N_300_cascade_\
        );

    \I__2464\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15640\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__15640\,
            I => \N__15637\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__15637\,
            I => \N__15634\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__15634\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\
        );

    \I__2460\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15628\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__15628\,
            I => \ppm_encoder_1.N_139_0\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__15625\,
            I => \N__15622\
        );

    \I__2457\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15619\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__15619\,
            I => \ppm_encoder_1.un2_throttle_iv_0_14\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__15616\,
            I => \N__15613\
        );

    \I__2454\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15610\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__15610\,
            I => \N__15607\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__15607\,
            I => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\
        );

    \I__2451\ : InMux
    port map (
            O => \N__15604\,
            I => \N__15601\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__15601\,
            I => \ppm_encoder_1.un2_throttle_iv_1_14\
        );

    \I__2449\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15593\
        );

    \I__2448\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15588\
        );

    \I__2447\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15588\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__15593\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__15588\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__2444\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15579\
        );

    \I__2443\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15576\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__15579\,
            I => \N__15573\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__15576\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__15573\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__2439\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15563\
        );

    \I__2438\ : InMux
    port map (
            O => \N__15567\,
            I => \N__15558\
        );

    \I__2437\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15558\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__15563\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__15558\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__2434\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15549\
        );

    \I__2433\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15546\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__15549\,
            I => \N__15543\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__15546\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__15543\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__2429\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15535\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__15535\,
            I => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__15532\,
            I => \Commands_frame_decoder.WDT8lto13_1_cascade_\
        );

    \I__2426\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15526\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__15526\,
            I => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\
        );

    \I__2424\ : IoInMux
    port map (
            O => \N__15523\,
            I => \N__15520\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__15520\,
            I => \N__15517\
        );

    \I__2422\ : Span4Mux_s2_v
    port map (
            O => \N__15517\,
            I => \N__15514\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__15514\,
            I => \N__15511\
        );

    \I__2420\ : Sp12to4
    port map (
            O => \N__15511\,
            I => \N__15508\
        );

    \I__2419\ : Span12Mux_h
    port map (
            O => \N__15508\,
            I => \N__15504\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__15507\,
            I => \N__15501\
        );

    \I__2417\ : Span12Mux_v
    port map (
            O => \N__15504\,
            I => \N__15498\
        );

    \I__2416\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15495\
        );

    \I__2415\ : Odrv12
    port map (
            O => \N__15498\,
            I => ppm_output_c
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__15495\,
            I => ppm_output_c
        );

    \I__2413\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15487\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15484\
        );

    \I__2411\ : Span4Mux_s1_v
    port map (
            O => \N__15484\,
            I => \N__15480\
        );

    \I__2410\ : InMux
    port map (
            O => \N__15483\,
            I => \N__15476\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__15480\,
            I => \N__15473\
        );

    \I__2408\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15470\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__15476\,
            I => \N__15465\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__15473\,
            I => \N__15465\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__15470\,
            I => \N__15462\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__15465\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__15462\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__2402\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15452\
        );

    \I__2401\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15449\
        );

    \I__2400\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15446\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__15452\,
            I => \N__15443\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__15449\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__15446\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__15443\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__2395\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15432\
        );

    \I__2394\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15429\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__15432\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__15429\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__2391\ : InMux
    port map (
            O => \N__15424\,
            I => \bfn_4_19_0_\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__15421\,
            I => \N__15417\
        );

    \I__2389\ : InMux
    port map (
            O => \N__15420\,
            I => \N__15414\
        );

    \I__2388\ : InMux
    port map (
            O => \N__15417\,
            I => \N__15411\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__15414\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__15411\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__2385\ : InMux
    port map (
            O => \N__15406\,
            I => \Commands_frame_decoder.un1_WDT_cry_8\
        );

    \I__2384\ : InMux
    port map (
            O => \N__15403\,
            I => \Commands_frame_decoder.un1_WDT_cry_9\
        );

    \I__2383\ : InMux
    port map (
            O => \N__15400\,
            I => \Commands_frame_decoder.un1_WDT_cry_10\
        );

    \I__2382\ : InMux
    port map (
            O => \N__15397\,
            I => \Commands_frame_decoder.un1_WDT_cry_11\
        );

    \I__2381\ : InMux
    port map (
            O => \N__15394\,
            I => \Commands_frame_decoder.un1_WDT_cry_12\
        );

    \I__2380\ : InMux
    port map (
            O => \N__15391\,
            I => \Commands_frame_decoder.un1_WDT_cry_13\
        );

    \I__2379\ : InMux
    port map (
            O => \N__15388\,
            I => \Commands_frame_decoder.un1_WDT_cry_14\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__15385\,
            I => \N__15381\
        );

    \I__2377\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15378\
        );

    \I__2376\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15375\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__15378\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__15375\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__2373\ : InMux
    port map (
            O => \N__15370\,
            I => \N__15366\
        );

    \I__2372\ : InMux
    port map (
            O => \N__15369\,
            I => \N__15363\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__15366\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__15363\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__2369\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15355\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__15355\,
            I => \Commands_frame_decoder.WDTZ0Z_0\
        );

    \I__2367\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15349\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__15349\,
            I => \Commands_frame_decoder.WDTZ0Z_1\
        );

    \I__2365\ : InMux
    port map (
            O => \N__15346\,
            I => \Commands_frame_decoder.un1_WDT_cry_0\
        );

    \I__2364\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15340\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__15340\,
            I => \Commands_frame_decoder.WDTZ0Z_2\
        );

    \I__2362\ : InMux
    port map (
            O => \N__15337\,
            I => \Commands_frame_decoder.un1_WDT_cry_1\
        );

    \I__2361\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15331\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__15331\,
            I => \Commands_frame_decoder.WDTZ0Z_3\
        );

    \I__2359\ : InMux
    port map (
            O => \N__15328\,
            I => \Commands_frame_decoder.un1_WDT_cry_2\
        );

    \I__2358\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15321\
        );

    \I__2357\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15318\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__15321\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__15318\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__2354\ : InMux
    port map (
            O => \N__15313\,
            I => \Commands_frame_decoder.un1_WDT_cry_3\
        );

    \I__2353\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15306\
        );

    \I__2352\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15303\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__15306\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__15303\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__2349\ : InMux
    port map (
            O => \N__15298\,
            I => \Commands_frame_decoder.un1_WDT_cry_4\
        );

    \I__2348\ : InMux
    port map (
            O => \N__15295\,
            I => \Commands_frame_decoder.un1_WDT_cry_5\
        );

    \I__2347\ : InMux
    port map (
            O => \N__15292\,
            I => \Commands_frame_decoder.un1_WDT_cry_6\
        );

    \I__2346\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15284\
        );

    \I__2345\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15278\
        );

    \I__2344\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15278\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__15284\,
            I => \N__15275\
        );

    \I__2342\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15272\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__15278\,
            I => \N__15269\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__15275\,
            I => \N__15264\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__15272\,
            I => \N__15264\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__15269\,
            I => \N__15261\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__15264\,
            I => uart_drone_data_2
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__15261\,
            I => uart_drone_data_2
        );

    \I__2335\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15249\
        );

    \I__2334\ : InMux
    port map (
            O => \N__15255\,
            I => \N__15244\
        );

    \I__2333\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15244\
        );

    \I__2332\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15241\
        );

    \I__2331\ : InMux
    port map (
            O => \N__15252\,
            I => \N__15238\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__15249\,
            I => \N__15235\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__15244\,
            I => \N__15230\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__15241\,
            I => \N__15225\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__15238\,
            I => \N__15225\
        );

    \I__2326\ : Span4Mux_h
    port map (
            O => \N__15235\,
            I => \N__15222\
        );

    \I__2325\ : InMux
    port map (
            O => \N__15234\,
            I => \N__15219\
        );

    \I__2324\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15216\
        );

    \I__2323\ : Span4Mux_h
    port map (
            O => \N__15230\,
            I => \N__15213\
        );

    \I__2322\ : Span4Mux_h
    port map (
            O => \N__15225\,
            I => \N__15210\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__15222\,
            I => uart_drone_data_3
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__15219\,
            I => uart_drone_data_3
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__15216\,
            I => uart_drone_data_3
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__15213\,
            I => uart_drone_data_3
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__15210\,
            I => uart_drone_data_3
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__15199\,
            I => \N__15196\
        );

    \I__2315\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15193\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__15193\,
            I => \N__15186\
        );

    \I__2313\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15183\
        );

    \I__2312\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15180\
        );

    \I__2311\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15175\
        );

    \I__2310\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15175\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__15186\,
            I => \N__15170\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__15183\,
            I => \N__15170\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__15180\,
            I => \N__15166\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__15175\,
            I => \N__15162\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__15170\,
            I => \N__15159\
        );

    \I__2304\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15156\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__15166\,
            I => \N__15153\
        );

    \I__2302\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15150\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__15162\,
            I => \N__15147\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__15159\,
            I => uart_drone_data_4
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__15156\,
            I => uart_drone_data_4
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__15153\,
            I => uart_drone_data_4
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__15150\,
            I => uart_drone_data_4
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__15147\,
            I => uart_drone_data_4
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__15136\,
            I => \N__15133\
        );

    \I__2294\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15129\
        );

    \I__2293\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15126\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__15129\,
            I => \N__15122\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__15126\,
            I => \N__15119\
        );

    \I__2290\ : InMux
    port map (
            O => \N__15125\,
            I => \N__15116\
        );

    \I__2289\ : Span4Mux_h
    port map (
            O => \N__15122\,
            I => \N__15113\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__15119\,
            I => \N__15108\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__15116\,
            I => \N__15108\
        );

    \I__2286\ : Span4Mux_h
    port map (
            O => \N__15113\,
            I => \N__15104\
        );

    \I__2285\ : Span4Mux_h
    port map (
            O => \N__15108\,
            I => \N__15101\
        );

    \I__2284\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15098\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__15104\,
            I => uart_drone_data_5
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__15101\,
            I => uart_drone_data_5
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__15098\,
            I => uart_drone_data_5
        );

    \I__2280\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15079\
        );

    \I__2279\ : InMux
    port map (
            O => \N__15090\,
            I => \N__15070\
        );

    \I__2278\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15070\
        );

    \I__2277\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15070\
        );

    \I__2276\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15070\
        );

    \I__2275\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15067\
        );

    \I__2274\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15062\
        );

    \I__2273\ : InMux
    port map (
            O => \N__15084\,
            I => \N__15062\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15057\
        );

    \I__2271\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15057\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15079\,
            I => \N__15054\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__15070\,
            I => \N__15051\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__15067\,
            I => \N__15044\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__15062\,
            I => \N__15044\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__15057\,
            I => \N__15041\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__15054\,
            I => \N__15036\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__15051\,
            I => \N__15036\
        );

    \I__2263\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15033\
        );

    \I__2262\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15030\
        );

    \I__2261\ : Span4Mux_h
    port map (
            O => \N__15044\,
            I => \N__15025\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__15041\,
            I => \N__15025\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__15036\,
            I => uart_drone_data_6
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__15033\,
            I => uart_drone_data_6
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__15030\,
            I => uart_drone_data_6
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__15025\,
            I => uart_drone_data_6
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__15016\,
            I => \N__15008\
        );

    \I__2254\ : InMux
    port map (
            O => \N__15015\,
            I => \N__15003\
        );

    \I__2253\ : InMux
    port map (
            O => \N__15014\,
            I => \N__15000\
        );

    \I__2252\ : InMux
    port map (
            O => \N__15013\,
            I => \N__14993\
        );

    \I__2251\ : InMux
    port map (
            O => \N__15012\,
            I => \N__14993\
        );

    \I__2250\ : InMux
    port map (
            O => \N__15011\,
            I => \N__14993\
        );

    \I__2249\ : InMux
    port map (
            O => \N__15008\,
            I => \N__14990\
        );

    \I__2248\ : InMux
    port map (
            O => \N__15007\,
            I => \N__14985\
        );

    \I__2247\ : InMux
    port map (
            O => \N__15006\,
            I => \N__14985\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__15003\,
            I => \N__14980\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__15000\,
            I => \N__14980\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__14993\,
            I => \N__14977\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__14990\,
            I => \N__14972\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__14985\,
            I => \N__14972\
        );

    \I__2241\ : Span4Mux_v
    port map (
            O => \N__14980\,
            I => \N__14968\
        );

    \I__2240\ : Span4Mux_h
    port map (
            O => \N__14977\,
            I => \N__14965\
        );

    \I__2239\ : Span4Mux_h
    port map (
            O => \N__14972\,
            I => \N__14962\
        );

    \I__2238\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14959\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__14968\,
            I => uart_drone_data_7
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__14965\,
            I => uart_drone_data_7
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__14962\,
            I => uart_drone_data_7
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__14959\,
            I => uart_drone_data_7
        );

    \I__2233\ : CEMux
    port map (
            O => \N__14950\,
            I => \N__14947\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__14947\,
            I => \uart_drone.state_1_sqmuxa_0\
        );

    \I__2231\ : SRMux
    port map (
            O => \N__14944\,
            I => \N__14941\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__14941\,
            I => \N__14938\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__14938\,
            I => \N__14935\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__14935\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__14932\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_\
        );

    \I__2226\ : InMux
    port map (
            O => \N__14929\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__2225\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14920\
        );

    \I__2224\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14920\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__14920\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__2222\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14913\
        );

    \I__2221\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14910\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__14913\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__14910\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__14905\,
            I => \N__14901\
        );

    \I__2217\ : InMux
    port map (
            O => \N__14904\,
            I => \N__14896\
        );

    \I__2216\ : InMux
    port map (
            O => \N__14901\,
            I => \N__14896\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__14896\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__2214\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14889\
        );

    \I__2213\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14886\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__14889\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__14886\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__2210\ : InMux
    port map (
            O => \N__14881\,
            I => \N__14878\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14875\
        );

    \I__2208\ : Odrv12
    port map (
            O => \N__14875\,
            I => \reset_module_System.reset6_11\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__14872\,
            I => \N__14869\
        );

    \I__2206\ : InMux
    port map (
            O => \N__14869\,
            I => \N__14866\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__14866\,
            I => \N__14863\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__14863\,
            I => \dron_frame_decoder_1.state_ns_i_a2_0_3_0\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__14860\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__14857\,
            I => \N__14854\
        );

    \I__2201\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14851\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__14851\,
            I => \Commands_frame_decoder.state_1_ns_0_a4_0_0_2\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__14848\,
            I => \N__14844\
        );

    \I__2198\ : InMux
    port map (
            O => \N__14847\,
            I => \N__14841\
        );

    \I__2197\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14838\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__14841\,
            I => \N__14835\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__14838\,
            I => \N__14832\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__14835\,
            I => \N__14828\
        );

    \I__2193\ : Span4Mux_v
    port map (
            O => \N__14832\,
            I => \N__14825\
        );

    \I__2192\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14822\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__14828\,
            I => uart_drone_data_0
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__14825\,
            I => uart_drone_data_0
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__14822\,
            I => uart_drone_data_0
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__14815\,
            I => \N__14811\
        );

    \I__2187\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14805\
        );

    \I__2186\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14800\
        );

    \I__2185\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14800\
        );

    \I__2184\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14794\
        );

    \I__2183\ : InMux
    port map (
            O => \N__14808\,
            I => \N__14794\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__14805\,
            I => \N__14790\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__14800\,
            I => \N__14787\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__14799\,
            I => \N__14784\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14781\
        );

    \I__2178\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14778\
        );

    \I__2177\ : Span4Mux_v
    port map (
            O => \N__14790\,
            I => \N__14773\
        );

    \I__2176\ : Span4Mux_v
    port map (
            O => \N__14787\,
            I => \N__14773\
        );

    \I__2175\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14770\
        );

    \I__2174\ : Span4Mux_v
    port map (
            O => \N__14781\,
            I => \N__14765\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__14778\,
            I => \N__14765\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__14773\,
            I => uart_drone_data_1
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__14770\,
            I => uart_drone_data_1
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__14765\,
            I => uart_drone_data_1
        );

    \I__2169\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14755\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__14755\,
            I => \N__14751\
        );

    \I__2167\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14748\
        );

    \I__2166\ : Odrv12
    port map (
            O => \N__14751\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__14748\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__2164\ : InMux
    port map (
            O => \N__14743\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__2163\ : InMux
    port map (
            O => \N__14740\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__2162\ : InMux
    port map (
            O => \N__14737\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__2161\ : InMux
    port map (
            O => \N__14734\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__2160\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14727\
        );

    \I__2159\ : InMux
    port map (
            O => \N__14730\,
            I => \N__14724\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__14727\,
            I => \N__14721\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__14724\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__14721\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__2155\ : InMux
    port map (
            O => \N__14716\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__2154\ : InMux
    port map (
            O => \N__14713\,
            I => \bfn_4_14_0_\
        );

    \I__2153\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14706\
        );

    \I__2152\ : InMux
    port map (
            O => \N__14709\,
            I => \N__14703\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__14706\,
            I => \N__14700\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__14703\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__14700\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__2148\ : InMux
    port map (
            O => \N__14695\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__2147\ : InMux
    port map (
            O => \N__14692\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__2146\ : InMux
    port map (
            O => \N__14689\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__2145\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14682\
        );

    \I__2144\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14679\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__14682\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__14679\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__2141\ : InMux
    port map (
            O => \N__14674\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__2140\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14667\
        );

    \I__2139\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14664\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__14667\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__14664\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__2136\ : InMux
    port map (
            O => \N__14659\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__2135\ : InMux
    port map (
            O => \N__14656\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__2134\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14649\
        );

    \I__2133\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14646\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__14649\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__14646\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__2130\ : InMux
    port map (
            O => \N__14641\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__2129\ : InMux
    port map (
            O => \N__14638\,
            I => \N__14634\
        );

    \I__2128\ : InMux
    port map (
            O => \N__14637\,
            I => \N__14631\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__14634\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__14631\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__2125\ : InMux
    port map (
            O => \N__14626\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__14623\,
            I => \N__14620\
        );

    \I__2123\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14616\
        );

    \I__2122\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14613\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__14616\,
            I => \N__14610\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__14613\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__14610\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__2118\ : InMux
    port map (
            O => \N__14605\,
            I => \bfn_4_13_0_\
        );

    \I__2117\ : InMux
    port map (
            O => \N__14602\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__2116\ : InMux
    port map (
            O => \N__14599\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__14596\,
            I => \reset_module_System.reset6_13_cascade_\
        );

    \I__2114\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14590\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__14590\,
            I => \reset_module_System.reset6_3\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__14587\,
            I => \reset_module_System.reset6_17_cascade_\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__14584\,
            I => \reset_module_System.reset6_19_cascade_\
        );

    \I__2110\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14577\
        );

    \I__2109\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14573\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__14577\,
            I => \N__14570\
        );

    \I__2107\ : InMux
    port map (
            O => \N__14576\,
            I => \N__14567\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__14573\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__14570\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__14567\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__14560\,
            I => \N__14554\
        );

    \I__2102\ : InMux
    port map (
            O => \N__14559\,
            I => \N__14551\
        );

    \I__2101\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14546\
        );

    \I__2100\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14546\
        );

    \I__2099\ : InMux
    port map (
            O => \N__14554\,
            I => \N__14543\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__14551\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__14546\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__14543\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__2095\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14533\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__14533\,
            I => \reset_module_System.count_1_2\
        );

    \I__2093\ : InMux
    port map (
            O => \N__14530\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__2092\ : InMux
    port map (
            O => \N__14527\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__2091\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__14521\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_16\
        );

    \I__2089\ : InMux
    port map (
            O => \N__14518\,
            I => \N__14515\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__14515\,
            I => \N__14512\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__14512\,
            I => \N__14509\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__14509\,
            I => \ppm_encoder_1.un1_init_pulses_11_16\
        );

    \I__2085\ : InMux
    port map (
            O => \N__14506\,
            I => \N__14503\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__14503\,
            I => \ppm_encoder_1.un1_init_pulses_10_16\
        );

    \I__2083\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14497\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__14497\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\
        );

    \I__2081\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14491\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__14491\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\
        );

    \I__2079\ : InMux
    port map (
            O => \N__14488\,
            I => \N__14485\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__14485\,
            I => \ppm_encoder_1.pulses2countZ0Z_8\
        );

    \I__2077\ : InMux
    port map (
            O => \N__14482\,
            I => \N__14479\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__14479\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__14476\,
            I => \N__14473\
        );

    \I__2074\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14470\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__14470\,
            I => \ppm_encoder_1.pulses2countZ0Z_9\
        );

    \I__2072\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14463\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__14466\,
            I => \N__14459\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__14463\,
            I => \N__14456\
        );

    \I__2069\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14453\
        );

    \I__2068\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14450\
        );

    \I__2067\ : Span12Mux_h
    port map (
            O => \N__14456\,
            I => \N__14445\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__14453\,
            I => \N__14445\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__14450\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__14445\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__2063\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14437\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14434\
        );

    \I__2061\ : Odrv12
    port map (
            O => \N__14434\,
            I => \ppm_encoder_1.N_295\
        );

    \I__2060\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14428\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__14428\,
            I => \N__14424\
        );

    \I__2058\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14421\
        );

    \I__2057\ : Odrv12
    port map (
            O => \N__14424\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__14421\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__14416\,
            I => \reset_module_System.count_1_1_cascade_\
        );

    \I__2054\ : InMux
    port map (
            O => \N__14413\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_12\
        );

    \I__2053\ : InMux
    port map (
            O => \N__14410\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_13\
        );

    \I__2052\ : InMux
    port map (
            O => \N__14407\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_14\
        );

    \I__2051\ : InMux
    port map (
            O => \N__14404\,
            I => \bfn_3_27_0_\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__14401\,
            I => \N__14398\
        );

    \I__2049\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14395\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__14395\,
            I => \ppm_encoder_1.un1_init_pulses_10_17\
        );

    \I__2047\ : InMux
    port map (
            O => \N__14392\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_16\
        );

    \I__2046\ : InMux
    port map (
            O => \N__14389\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_17\
        );

    \I__2045\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14383\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__14383\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_17\
        );

    \I__2043\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14375\
        );

    \I__2042\ : InMux
    port map (
            O => \N__14379\,
            I => \N__14370\
        );

    \I__2041\ : InMux
    port map (
            O => \N__14378\,
            I => \N__14370\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__14375\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__14370\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__14365\,
            I => \N__14362\
        );

    \I__2037\ : InMux
    port map (
            O => \N__14362\,
            I => \N__14359\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__14359\,
            I => \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\
        );

    \I__2035\ : InMux
    port map (
            O => \N__14356\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_4\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__14353\,
            I => \N__14350\
        );

    \I__2033\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14347\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__14347\,
            I => \N__14344\
        );

    \I__2031\ : Span4Mux_v
    port map (
            O => \N__14344\,
            I => \N__14341\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__14341\,
            I => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\
        );

    \I__2029\ : InMux
    port map (
            O => \N__14338\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_5\
        );

    \I__2028\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14331\
        );

    \I__2027\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14328\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__14331\,
            I => \N__14325\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__14328\,
            I => \N__14322\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__14325\,
            I => \N__14319\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__14322\,
            I => \N__14316\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__14319\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__14316\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__14311\,
            I => \N__14308\
        );

    \I__2019\ : InMux
    port map (
            O => \N__14308\,
            I => \N__14305\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__14305\,
            I => \N__14302\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__14302\,
            I => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\
        );

    \I__2016\ : InMux
    port map (
            O => \N__14299\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_6\
        );

    \I__2015\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14293\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__14293\,
            I => \N__14289\
        );

    \I__2013\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14286\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__14289\,
            I => \N__14281\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__14286\,
            I => \N__14281\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__14281\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__14278\,
            I => \N__14275\
        );

    \I__2008\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14272\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__14272\,
            I => \N__14269\
        );

    \I__2006\ : Odrv12
    port map (
            O => \N__14269\,
            I => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\
        );

    \I__2005\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14263\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14260\
        );

    \I__2003\ : Span4Mux_s2_v
    port map (
            O => \N__14260\,
            I => \N__14257\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__14257\,
            I => \ppm_encoder_1.un1_init_pulses_10_8\
        );

    \I__2001\ : InMux
    port map (
            O => \N__14254\,
            I => \bfn_3_26_0_\
        );

    \I__2000\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14248\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__14248\,
            I => \N__14244\
        );

    \I__1998\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14241\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__14244\,
            I => \N__14236\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14236\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__14236\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__14233\,
            I => \N__14230\
        );

    \I__1993\ : InMux
    port map (
            O => \N__14230\,
            I => \N__14227\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__14227\,
            I => \N__14224\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__14224\,
            I => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\
        );

    \I__1990\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14218\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__14218\,
            I => \N__14215\
        );

    \I__1988\ : Span4Mux_s3_v
    port map (
            O => \N__14215\,
            I => \N__14212\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__14212\,
            I => \ppm_encoder_1.un1_init_pulses_10_9\
        );

    \I__1986\ : InMux
    port map (
            O => \N__14209\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_8\
        );

    \I__1985\ : InMux
    port map (
            O => \N__14206\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_9\
        );

    \I__1984\ : InMux
    port map (
            O => \N__14203\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_10\
        );

    \I__1983\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14196\
        );

    \I__1982\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14193\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__14196\,
            I => \N__14190\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__14193\,
            I => \N__14187\
        );

    \I__1979\ : Span4Mux_h
    port map (
            O => \N__14190\,
            I => \N__14182\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__14187\,
            I => \N__14182\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__14182\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__14179\,
            I => \N__14176\
        );

    \I__1975\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14173\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__14173\,
            I => \N__14170\
        );

    \I__1973\ : Odrv12
    port map (
            O => \N__14170\,
            I => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\
        );

    \I__1972\ : InMux
    port map (
            O => \N__14167\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_11\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__14164\,
            I => \N__14161\
        );

    \I__1970\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14158\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__1968\ : Span4Mux_v
    port map (
            O => \N__14155\,
            I => \N__14152\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__14152\,
            I => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__14149\,
            I => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\
        );

    \I__1965\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14143\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__14143\,
            I => \ppm_encoder_1.un2_throttle_iv_1_5\
        );

    \I__1963\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14137\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__14137\,
            I => \N__14134\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__14134\,
            I => \ppm_encoder_1.throttle_RNIN3352Z0Z_0\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__14131\,
            I => \N__14128\
        );

    \I__1959\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14124\
        );

    \I__1958\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14121\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__14124\,
            I => \N__14118\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__14121\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__14118\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__14113\,
            I => \N__14110\
        );

    \I__1953\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14107\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__14107\,
            I => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\
        );

    \I__1951\ : InMux
    port map (
            O => \N__14104\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_0\
        );

    \I__1950\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14098\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14094\
        );

    \I__1948\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14091\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__14094\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__14091\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__14086\,
            I => \N__14083\
        );

    \I__1944\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14080\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__14080\,
            I => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\
        );

    \I__1942\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14074\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__14074\,
            I => \ppm_encoder_1.un1_init_pulses_10_2\
        );

    \I__1940\ : InMux
    port map (
            O => \N__14071\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_1\
        );

    \I__1939\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14065\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__14065\,
            I => \N__14061\
        );

    \I__1937\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14058\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__14061\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__14058\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__14053\,
            I => \N__14050\
        );

    \I__1933\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14047\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__14047\,
            I => \N__14044\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__14044\,
            I => \ppm_encoder_1.throttle_RNI82223Z0Z_3\
        );

    \I__1930\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14038\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__14038\,
            I => \N__14035\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__14035\,
            I => \ppm_encoder_1.un1_init_pulses_10_3\
        );

    \I__1927\ : InMux
    port map (
            O => \N__14032\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_2\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__14029\,
            I => \N__14026\
        );

    \I__1925\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14023\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__14023\,
            I => \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\
        );

    \I__1923\ : InMux
    port map (
            O => \N__14020\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_3\
        );

    \I__1922\ : InMux
    port map (
            O => \N__14017\,
            I => \N__14014\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__14014\,
            I => \ppm_encoder_1.un2_throttle_iv_1_8\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__14011\,
            I => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\
        );

    \I__1919\ : InMux
    port map (
            O => \N__14008\,
            I => \N__14005\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__14005\,
            I => \ppm_encoder_1.un2_throttle_iv_1_9\
        );

    \I__1917\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13999\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__13999\,
            I => \ppm_encoder_1.un2_throttle_iv_1_4\
        );

    \I__1915\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13991\
        );

    \I__1914\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13988\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__13994\,
            I => \N__13985\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__13991\,
            I => \N__13982\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__13988\,
            I => \N__13979\
        );

    \I__1910\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13976\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__13982\,
            I => \N__13973\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__13979\,
            I => \N__13970\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__13976\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__13973\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__13970\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__1904\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13957\
        );

    \I__1903\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13957\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__13957\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__1901\ : InMux
    port map (
            O => \N__13954\,
            I => \N__13951\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__13951\,
            I => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\
        );

    \I__1899\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13945\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__13945\,
            I => \N__13941\
        );

    \I__1897\ : InMux
    port map (
            O => \N__13944\,
            I => \N__13938\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__13941\,
            I => \N__13935\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__13938\,
            I => \N__13932\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__13935\,
            I => \N__13929\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__13932\,
            I => \N__13926\
        );

    \I__1892\ : Span4Mux_v
    port map (
            O => \N__13929\,
            I => \N__13923\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__13926\,
            I => \N__13920\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__13923\,
            I => throttle_command_12
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__13920\,
            I => throttle_command_12
        );

    \I__1888\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13912\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__13912\,
            I => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__13909\,
            I => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\
        );

    \I__1885\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13903\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__13903\,
            I => \ppm_encoder_1.un2_throttle_iv_1_12\
        );

    \I__1883\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13895\
        );

    \I__1882\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13890\
        );

    \I__1881\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13890\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__13895\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__13890\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__13885\,
            I => \ppm_encoder_1.N_303_cascade_\
        );

    \I__1877\ : InMux
    port map (
            O => \N__13882\,
            I => \N__13873\
        );

    \I__1876\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13873\
        );

    \I__1875\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13873\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__13873\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__13870\,
            I => \N__13867\
        );

    \I__1872\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13862\
        );

    \I__1871\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13859\
        );

    \I__1870\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13856\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__13862\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__13859\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__13856\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__13849\,
            I => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\
        );

    \I__1865\ : IoInMux
    port map (
            O => \N__13846\,
            I => \N__13843\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__13843\,
            I => \N__13840\
        );

    \I__1863\ : IoSpan4Mux
    port map (
            O => \N__13840\,
            I => \N__13837\
        );

    \I__1862\ : Span4Mux_s3_v
    port map (
            O => \N__13837\,
            I => \N__13833\
        );

    \I__1861\ : InMux
    port map (
            O => \N__13836\,
            I => \N__13830\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__13833\,
            I => \N__13823\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__13830\,
            I => \N__13823\
        );

    \I__1858\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13818\
        );

    \I__1857\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13818\
        );

    \I__1856\ : Sp12to4
    port map (
            O => \N__13823\,
            I => \N__13815\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__13818\,
            I => drone_frame_decoder_data_rdy_debug_c
        );

    \I__1854\ : Odrv12
    port map (
            O => \N__13815\,
            I => drone_frame_decoder_data_rdy_debug_c
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__13810\,
            I => \uart_pc.N_152_cascade_\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__13807\,
            I => \uart_pc.CO0_cascade_\
        );

    \I__1851\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13798\
        );

    \I__1850\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13798\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__13798\,
            I => \uart_pc.un1_state_7_0\
        );

    \I__1848\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13792\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__13792\,
            I => \N__13788\
        );

    \I__1846\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13785\
        );

    \I__1845\ : Span4Mux_h
    port map (
            O => \N__13788\,
            I => \N__13780\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__13785\,
            I => \N__13780\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__13780\,
            I => \N__13777\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__13777\,
            I => \N__13774\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__13774\,
            I => throttle_command_9
        );

    \I__1840\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13768\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__13768\,
            I => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\
        );

    \I__1838\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13762\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__13762\,
            I => \N__13759\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__13759\,
            I => \N__13756\
        );

    \I__1835\ : Sp12to4
    port map (
            O => \N__13756\,
            I => \N__13752\
        );

    \I__1834\ : InMux
    port map (
            O => \N__13755\,
            I => \N__13749\
        );

    \I__1833\ : Span12Mux_s2_h
    port map (
            O => \N__13752\,
            I => \N__13744\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__13749\,
            I => \N__13744\
        );

    \I__1831\ : Span12Mux_v
    port map (
            O => \N__13744\,
            I => \N__13741\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__13741\,
            I => throttle_command_11
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__13738\,
            I => \N__13735\
        );

    \I__1828\ : InMux
    port map (
            O => \N__13735\,
            I => \N__13732\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__13732\,
            I => \N__13729\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__13729\,
            I => alt_command_7
        );

    \I__1825\ : CEMux
    port map (
            O => \N__13726\,
            I => \N__13723\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__13723\,
            I => \N__13718\
        );

    \I__1823\ : CEMux
    port map (
            O => \N__13722\,
            I => \N__13715\
        );

    \I__1822\ : CEMux
    port map (
            O => \N__13721\,
            I => \N__13712\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__13718\,
            I => \N__13707\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__13715\,
            I => \N__13707\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__13712\,
            I => \N__13704\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__13707\,
            I => \N__13699\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__13704\,
            I => \N__13699\
        );

    \I__1816\ : Span4Mux_s2_h
    port map (
            O => \N__13699\,
            I => \N__13696\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__13696\,
            I => \dron_frame_decoder_1.N_238_0\
        );

    \I__1814\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13690\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__13690\,
            I => \N__13686\
        );

    \I__1812\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13677\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__13686\,
            I => \N__13674\
        );

    \I__1810\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13663\
        );

    \I__1809\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13663\
        );

    \I__1808\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13663\
        );

    \I__1807\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13663\
        );

    \I__1806\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13663\
        );

    \I__1805\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13660\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__13677\,
            I => \dron_frame_decoder_1.N_237\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__13674\,
            I => \dron_frame_decoder_1.N_237\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__13663\,
            I => \dron_frame_decoder_1.N_237\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__13660\,
            I => \dron_frame_decoder_1.N_237\
        );

    \I__1800\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13647\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__13650\,
            I => \N__13644\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__13647\,
            I => \N__13640\
        );

    \I__1797\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13635\
        );

    \I__1796\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13635\
        );

    \I__1795\ : Odrv12
    port map (
            O => \N__13640\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__13635\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__1793\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13627\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__13627\,
            I => \dron_frame_decoder_1.un1_sink_data_valid_5_0_0\
        );

    \I__1791\ : InMux
    port map (
            O => \N__13624\,
            I => \N__13621\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__13621\,
            I => \N__13616\
        );

    \I__1789\ : InMux
    port map (
            O => \N__13620\,
            I => \N__13611\
        );

    \I__1788\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13611\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__13616\,
            I => \N__13608\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__13611\,
            I => \dron_frame_decoder_1.stateZ0Z_7\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__13608\,
            I => \dron_frame_decoder_1.stateZ0Z_7\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__13603\,
            I => \N__13599\
        );

    \I__1783\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13590\
        );

    \I__1782\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13590\
        );

    \I__1781\ : InMux
    port map (
            O => \N__13598\,
            I => \N__13590\
        );

    \I__1780\ : InMux
    port map (
            O => \N__13597\,
            I => \N__13587\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13584\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__13587\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__13584\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__13579\,
            I => \dron_frame_decoder_1.un1_sink_data_valid_5_0_0_cascade_\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__13576\,
            I => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_\
        );

    \I__1774\ : CEMux
    port map (
            O => \N__13573\,
            I => \N__13569\
        );

    \I__1773\ : CEMux
    port map (
            O => \N__13572\,
            I => \N__13565\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__13569\,
            I => \N__13562\
        );

    \I__1771\ : CEMux
    port map (
            O => \N__13568\,
            I => \N__13559\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__13565\,
            I => \N__13556\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__13562\,
            I => \N__13553\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__13559\,
            I => \N__13550\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__13556\,
            I => \N__13547\
        );

    \I__1766\ : Span4Mux_s3_h
    port map (
            O => \N__13553\,
            I => \N__13544\
        );

    \I__1765\ : Sp12to4
    port map (
            O => \N__13550\,
            I => \N__13541\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__13547\,
            I => \dron_frame_decoder_1.N_230_0\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__13544\,
            I => \dron_frame_decoder_1.N_230_0\
        );

    \I__1762\ : Odrv12
    port map (
            O => \N__13541\,
            I => \dron_frame_decoder_1.N_230_0\
        );

    \I__1761\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13527\
        );

    \I__1760\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13527\
        );

    \I__1759\ : InMux
    port map (
            O => \N__13532\,
            I => \N__13522\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__13527\,
            I => \N__13518\
        );

    \I__1757\ : InMux
    port map (
            O => \N__13526\,
            I => \N__13515\
        );

    \I__1756\ : InMux
    port map (
            O => \N__13525\,
            I => \N__13512\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__13522\,
            I => \N__13509\
        );

    \I__1754\ : InMux
    port map (
            O => \N__13521\,
            I => \N__13506\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__13518\,
            I => \N__13501\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__13515\,
            I => \N__13501\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__13512\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__13509\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__13506\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__13501\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__1747\ : IoInMux
    port map (
            O => \N__13492\,
            I => \N__13489\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__13489\,
            I => \N__13486\
        );

    \I__1745\ : IoSpan4Mux
    port map (
            O => \N__13486\,
            I => \N__13479\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__13485\,
            I => \N__13475\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__13484\,
            I => \N__13472\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__13483\,
            I => \N__13469\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__13482\,
            I => \N__13465\
        );

    \I__1740\ : Sp12to4
    port map (
            O => \N__13479\,
            I => \N__13461\
        );

    \I__1739\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13451\
        );

    \I__1738\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13451\
        );

    \I__1737\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13451\
        );

    \I__1736\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13451\
        );

    \I__1735\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13448\
        );

    \I__1734\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13445\
        );

    \I__1733\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13442\
        );

    \I__1732\ : Span12Mux_s9_v
    port map (
            O => \N__13461\,
            I => \N__13438\
        );

    \I__1731\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13435\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__13451\,
            I => \N__13430\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__13448\,
            I => \N__13430\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__13445\,
            I => \N__13425\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__13442\,
            I => \N__13425\
        );

    \I__1726\ : InMux
    port map (
            O => \N__13441\,
            I => \N__13420\
        );

    \I__1725\ : Span12Mux_h
    port map (
            O => \N__13438\,
            I => \N__13415\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__13435\,
            I => \N__13415\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__13430\,
            I => \N__13410\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__13425\,
            I => \N__13410\
        );

    \I__1721\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13405\
        );

    \I__1720\ : InMux
    port map (
            O => \N__13423\,
            I => \N__13405\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__13420\,
            I => uart_drone_data_rdy_debug_c
        );

    \I__1718\ : Odrv12
    port map (
            O => \N__13415\,
            I => uart_drone_data_rdy_debug_c
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__13410\,
            I => uart_drone_data_rdy_debug_c
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__13405\,
            I => uart_drone_data_rdy_debug_c
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__13396\,
            I => \dron_frame_decoder_1.state_ns_i_a2_1_1_0_cascade_\
        );

    \I__1714\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13390\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__13390\,
            I => \dron_frame_decoder_1.N_239\
        );

    \I__1712\ : InMux
    port map (
            O => \N__13387\,
            I => \N__13382\
        );

    \I__1711\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13375\
        );

    \I__1710\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13375\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__13382\,
            I => \N__13372\
        );

    \I__1708\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13367\
        );

    \I__1707\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13367\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__13375\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__13372\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__13367\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__1703\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13357\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__13357\,
            I => \dron_frame_decoder_1.state_ns_i_a2_0_2_0\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__13354\,
            I => \dron_frame_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_\
        );

    \I__1700\ : InMux
    port map (
            O => \N__13351\,
            I => \N__13348\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__13348\,
            I => \N__13344\
        );

    \I__1698\ : InMux
    port map (
            O => \N__13347\,
            I => \N__13341\
        );

    \I__1697\ : Span4Mux_s3_h
    port map (
            O => \N__13344\,
            I => \N__13335\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__13341\,
            I => \N__13335\
        );

    \I__1695\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13332\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__13335\,
            I => \dron_frame_decoder_1.N_243\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__13332\,
            I => \dron_frame_decoder_1.N_243\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__13327\,
            I => \N__13324\
        );

    \I__1691\ : InMux
    port map (
            O => \N__13324\,
            I => \N__13321\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13318\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__13318\,
            I => alt_command_4
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__13315\,
            I => \N__13312\
        );

    \I__1687\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13309\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13306\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__13306\,
            I => alt_command_5
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__13303\,
            I => \N__13300\
        );

    \I__1683\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13297\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__13297\,
            I => \N__13294\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__13294\,
            I => alt_command_6
        );

    \I__1680\ : InMux
    port map (
            O => \N__13291\,
            I => \N__13288\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__13288\,
            I => \dron_frame_decoder_1.state_ns_0_a3_0_3_3\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__13285\,
            I => \N__13281\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__13284\,
            I => \N__13278\
        );

    \I__1676\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13273\
        );

    \I__1675\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13273\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__13273\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__1673\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13264\
        );

    \I__1672\ : InMux
    port map (
            O => \N__13269\,
            I => \N__13264\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__13264\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__13261\,
            I => \dron_frame_decoder_1.N_217_cascade_\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__13258\,
            I => \N__13254\
        );

    \I__1668\ : InMux
    port map (
            O => \N__13257\,
            I => \N__13250\
        );

    \I__1667\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13247\
        );

    \I__1666\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13244\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__13250\,
            I => \N__13241\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__13247\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__13244\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__13241\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__1661\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__13231\,
            I => \dron_frame_decoder_1.N_219\
        );

    \I__1659\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__13225\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_9\
        );

    \I__1657\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13213\
        );

    \I__1656\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13213\
        );

    \I__1655\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13213\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__13213\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__1653\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13207\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__13207\,
            I => \N__13204\
        );

    \I__1651\ : Span4Mux_s2_v
    port map (
            O => \N__13204\,
            I => \N__13201\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__13201\,
            I => \N__13198\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__13198\,
            I => \ppm_encoder_1.N_299\
        );

    \I__1648\ : InMux
    port map (
            O => \N__13195\,
            I => \N__13191\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__13194\,
            I => \N__13188\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__13191\,
            I => \N__13185\
        );

    \I__1645\ : InMux
    port map (
            O => \N__13188\,
            I => \N__13182\
        );

    \I__1644\ : Span4Mux_s3_h
    port map (
            O => \N__13185\,
            I => \N__13179\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__13182\,
            I => alt_kp_7
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__13179\,
            I => alt_kp_7
        );

    \I__1641\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13170\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__13173\,
            I => \N__13167\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__13170\,
            I => \N__13164\
        );

    \I__1638\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13161\
        );

    \I__1637\ : Span4Mux_s3_h
    port map (
            O => \N__13164\,
            I => \N__13158\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__13161\,
            I => alt_kp_5
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__13158\,
            I => alt_kp_5
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__13153\,
            I => \dron_frame_decoder_1.state_ns_0_a3_0_0_3_cascade_\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__13150\,
            I => \dron_frame_decoder_1.state_ns_0_a3_0_0_1_cascade_\
        );

    \I__1632\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13144\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__13144\,
            I => \dron_frame_decoder_1.state_ns_0_a3_0_3_1\
        );

    \I__1630\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13138\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__13138\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__13135\,
            I => \N__13130\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__13134\,
            I => \N__13125\
        );

    \I__1626\ : InMux
    port map (
            O => \N__13133\,
            I => \N__13118\
        );

    \I__1625\ : InMux
    port map (
            O => \N__13130\,
            I => \N__13118\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \N__13115\
        );

    \I__1623\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13104\
        );

    \I__1622\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13104\
        );

    \I__1621\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13104\
        );

    \I__1620\ : InMux
    port map (
            O => \N__13123\,
            I => \N__13104\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__13118\,
            I => \N__13101\
        );

    \I__1618\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13096\
        );

    \I__1617\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13096\
        );

    \I__1616\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13093\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__13104\,
            I => \N__13090\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__13101\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__13096\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__13093\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__13090\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__1610\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13078\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__13078\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\
        );

    \I__1608\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13072\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__13072\,
            I => \N__13069\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__13069\,
            I => \ppm_encoder_1.un1_init_pulses_11_17\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__13066\,
            I => \N__13063\
        );

    \I__1604\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13060\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13060\,
            I => \N__13057\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__13057\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_17\
        );

    \I__1601\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13051\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__13051\,
            I => \ppm_encoder_1.un1_init_pulses_11_8\
        );

    \I__1599\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13045\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__13045\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_8\
        );

    \I__1597\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13033\
        );

    \I__1596\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13033\
        );

    \I__1595\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13033\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__13033\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__1593\ : InMux
    port map (
            O => \N__13030\,
            I => \N__13027\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__13027\,
            I => \ppm_encoder_1.un1_init_pulses_11_9\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__13024\,
            I => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__13021\,
            I => \ppm_encoder_1.un1_init_pulses_0_cascade_\
        );

    \I__1589\ : InMux
    port map (
            O => \N__13018\,
            I => \N__13015\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__13015\,
            I => \ppm_encoder_1.un1_init_pulses_10_0\
        );

    \I__1587\ : InMux
    port map (
            O => \N__13012\,
            I => \N__13009\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__13009\,
            I => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\
        );

    \I__1585\ : InMux
    port map (
            O => \N__13006\,
            I => \N__13003\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__13003\,
            I => \N__13000\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__13000\,
            I => \N__12996\
        );

    \I__1582\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12993\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__12996\,
            I => \N__12988\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__12993\,
            I => \N__12988\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__12988\,
            I => \N__12985\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__12985\,
            I => \N__12982\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__12982\,
            I => throttle_command_0
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__12979\,
            I => \N__12976\
        );

    \I__1575\ : InMux
    port map (
            O => \N__12976\,
            I => \N__12964\
        );

    \I__1574\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12964\
        );

    \I__1573\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12964\
        );

    \I__1572\ : InMux
    port map (
            O => \N__12973\,
            I => \N__12964\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__12964\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__12961\,
            I => \N__12958\
        );

    \I__1569\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12955\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__12955\,
            I => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__12952\,
            I => \N__12949\
        );

    \I__1566\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12946\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__12946\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__12943\,
            I => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__12940\,
            I => \N__12937\
        );

    \I__1562\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12934\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__12934\,
            I => \N__12931\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__12931\,
            I => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\
        );

    \I__1559\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12925\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__12925\,
            I => \N__12922\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__12922\,
            I => \ppm_encoder_1.un1_init_pulses_11_2\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__12919\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\
        );

    \I__1555\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12913\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__12913\,
            I => \N__12910\
        );

    \I__1553\ : Odrv12
    port map (
            O => \N__12910\,
            I => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\
        );

    \I__1552\ : InMux
    port map (
            O => \N__12907\,
            I => \N__12904\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__12904\,
            I => \N__12901\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__12901\,
            I => \N__12897\
        );

    \I__1549\ : InMux
    port map (
            O => \N__12900\,
            I => \N__12894\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__12897\,
            I => \N__12889\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__12894\,
            I => \N__12889\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__12889\,
            I => \N__12886\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__12886\,
            I => \N__12883\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__12883\,
            I => throttle_command_2
        );

    \I__1543\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12877\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__12877\,
            I => \N__12874\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__12874\,
            I => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__12871\,
            I => \ppm_encoder_1.PPM_STATE_58_d_cascade_\
        );

    \I__1539\ : InMux
    port map (
            O => \N__12868\,
            I => \N__12860\
        );

    \I__1538\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12860\
        );

    \I__1537\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12855\
        );

    \I__1536\ : InMux
    port map (
            O => \N__12865\,
            I => \N__12855\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__12860\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__12855\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__1533\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12846\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__12849\,
            I => \N__12843\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__12846\,
            I => \N__12839\
        );

    \I__1530\ : InMux
    port map (
            O => \N__12843\,
            I => \N__12834\
        );

    \I__1529\ : InMux
    port map (
            O => \N__12842\,
            I => \N__12834\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__12839\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__12834\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__12829\,
            I => \N__12825\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__12828\,
            I => \N__12822\
        );

    \I__1524\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12818\
        );

    \I__1523\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12813\
        );

    \I__1522\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12813\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__12818\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__12813\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__1519\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12803\
        );

    \I__1518\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12800\
        );

    \I__1517\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12797\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__12803\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__12800\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__12797\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__1513\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12786\
        );

    \I__1512\ : InMux
    port map (
            O => \N__12789\,
            I => \N__12783\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__12786\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__12783\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__12778\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\
        );

    \I__1508\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12771\
        );

    \I__1507\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12768\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__12771\,
            I => \N__12765\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__12768\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__12765\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__12760\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__12757\,
            I => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\
        );

    \I__1501\ : InMux
    port map (
            O => \N__12754\,
            I => \N__12751\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__12751\,
            I => \ppm_encoder_1.un2_throttle_iv_1_7\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__12748\,
            I => \N__12745\
        );

    \I__1498\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12740\
        );

    \I__1497\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12737\
        );

    \I__1496\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12734\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__12740\,
            I => \N__12731\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__12737\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__12734\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__12731\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__1491\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12719\
        );

    \I__1490\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12714\
        );

    \I__1489\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12714\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__12719\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__12714\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__12709\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__12706\,
            I => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\
        );

    \I__1484\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12700\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__12700\,
            I => \N__12696\
        );

    \I__1482\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12693\
        );

    \I__1481\ : Span4Mux_v
    port map (
            O => \N__12696\,
            I => \N__12688\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__12693\,
            I => \N__12688\
        );

    \I__1479\ : Span4Mux_v
    port map (
            O => \N__12688\,
            I => \N__12685\
        );

    \I__1478\ : Span4Mux_v
    port map (
            O => \N__12685\,
            I => \N__12682\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__12682\,
            I => throttle_command_1
        );

    \I__1476\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12676\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__12676\,
            I => \N__12673\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__12673\,
            I => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\
        );

    \I__1473\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12667\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__12667\,
            I => \N__12663\
        );

    \I__1471\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12660\
        );

    \I__1470\ : Span4Mux_h
    port map (
            O => \N__12663\,
            I => \N__12657\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__12660\,
            I => \N__12654\
        );

    \I__1468\ : Sp12to4
    port map (
            O => \N__12657\,
            I => \N__12649\
        );

    \I__1467\ : Span12Mux_h
    port map (
            O => \N__12654\,
            I => \N__12649\
        );

    \I__1466\ : Odrv12
    port map (
            O => \N__12649\,
            I => throttle_command_10
        );

    \I__1465\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12643\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__12643\,
            I => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\
        );

    \I__1463\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12636\
        );

    \I__1462\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12633\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__12636\,
            I => \N__12628\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12628\
        );

    \I__1459\ : Span4Mux_v
    port map (
            O => \N__12628\,
            I => \N__12625\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__12625\,
            I => \N__12622\
        );

    \I__1457\ : Span4Mux_v
    port map (
            O => \N__12622\,
            I => \N__12619\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__12619\,
            I => throttle_command_13
        );

    \I__1455\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12613\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__12613\,
            I => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\
        );

    \I__1453\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12607\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__12607\,
            I => \N__12603\
        );

    \I__1451\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12600\
        );

    \I__1450\ : Span4Mux_v
    port map (
            O => \N__12603\,
            I => \N__12595\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__12600\,
            I => \N__12595\
        );

    \I__1448\ : Span4Mux_v
    port map (
            O => \N__12595\,
            I => \N__12592\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__12592\,
            I => throttle_command_4
        );

    \I__1446\ : InMux
    port map (
            O => \N__12589\,
            I => \N__12586\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__12586\,
            I => \N__12583\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__12583\,
            I => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\
        );

    \I__1443\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12577\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__12577\,
            I => \N__12574\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__12574\,
            I => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\
        );

    \I__1440\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12568\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__12568\,
            I => \N__12564\
        );

    \I__1438\ : InMux
    port map (
            O => \N__12567\,
            I => \N__12561\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__12564\,
            I => \N__12556\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__12561\,
            I => \N__12556\
        );

    \I__1435\ : Span4Mux_v
    port map (
            O => \N__12556\,
            I => \N__12553\
        );

    \I__1434\ : Span4Mux_v
    port map (
            O => \N__12553\,
            I => \N__12550\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__12550\,
            I => throttle_command_5
        );

    \I__1432\ : InMux
    port map (
            O => \N__12547\,
            I => \N__12544\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__12544\,
            I => \N__12540\
        );

    \I__1430\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12537\
        );

    \I__1429\ : Span4Mux_v
    port map (
            O => \N__12540\,
            I => \N__12534\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__12537\,
            I => \N__12531\
        );

    \I__1427\ : Span4Mux_v
    port map (
            O => \N__12534\,
            I => \N__12526\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__12531\,
            I => \N__12526\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__12526\,
            I => \N__12523\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__12523\,
            I => throttle_command_8
        );

    \I__1423\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12517\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__12517\,
            I => \N__12514\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__12514\,
            I => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\
        );

    \I__1420\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12508\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__12508\,
            I => \N__12505\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__12505\,
            I => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\
        );

    \I__1417\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12499\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__12499\,
            I => \N__12495\
        );

    \I__1415\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12492\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__12495\,
            I => \N__12487\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__12492\,
            I => \N__12487\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__12487\,
            I => \N__12484\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__12484\,
            I => \N__12481\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__12481\,
            I => throttle_command_7
        );

    \I__1409\ : InMux
    port map (
            O => \N__12478\,
            I => \N__12474\
        );

    \I__1408\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12471\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__12474\,
            I => \N__12466\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__12471\,
            I => \N__12466\
        );

    \I__1405\ : Span4Mux_v
    port map (
            O => \N__12466\,
            I => \N__12463\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__12463\,
            I => \N__12460\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__12460\,
            I => throttle_command_6
        );

    \I__1402\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12454\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__12454\,
            I => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\
        );

    \I__1400\ : InMux
    port map (
            O => \N__12451\,
            I => \ppm_encoder_1.un1_throttle_cry_5\
        );

    \I__1399\ : InMux
    port map (
            O => \N__12448\,
            I => \ppm_encoder_1.un1_throttle_cry_6\
        );

    \I__1398\ : InMux
    port map (
            O => \N__12445\,
            I => \bfn_2_20_0_\
        );

    \I__1397\ : InMux
    port map (
            O => \N__12442\,
            I => \ppm_encoder_1.un1_throttle_cry_8\
        );

    \I__1396\ : InMux
    port map (
            O => \N__12439\,
            I => \ppm_encoder_1.un1_throttle_cry_9\
        );

    \I__1395\ : InMux
    port map (
            O => \N__12436\,
            I => \ppm_encoder_1.un1_throttle_cry_10\
        );

    \I__1394\ : InMux
    port map (
            O => \N__12433\,
            I => \ppm_encoder_1.un1_throttle_cry_11\
        );

    \I__1393\ : InMux
    port map (
            O => \N__12430\,
            I => \ppm_encoder_1.un1_throttle_cry_12\
        );

    \I__1392\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12424\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__12424\,
            I => \N__12421\
        );

    \I__1390\ : Span4Mux_v
    port map (
            O => \N__12421\,
            I => \N__12418\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__12418\,
            I => \N__12415\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__12415\,
            I => throttle_command_14
        );

    \I__1387\ : InMux
    port map (
            O => \N__12412\,
            I => \ppm_encoder_1.un1_throttle_cry_13\
        );

    \I__1386\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12406\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__12406\,
            I => drone_altitude_i_9
        );

    \I__1384\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12400\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__12400\,
            I => drone_altitude_14
        );

    \I__1382\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12394\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__12394\,
            I => \dron_frame_decoder_1.drone_altitude_9\
        );

    \I__1380\ : InMux
    port map (
            O => \N__12391\,
            I => \ppm_encoder_1.un1_throttle_cry_0\
        );

    \I__1379\ : InMux
    port map (
            O => \N__12388\,
            I => \ppm_encoder_1.un1_throttle_cry_1\
        );

    \I__1378\ : InMux
    port map (
            O => \N__12385\,
            I => \N__12381\
        );

    \I__1377\ : InMux
    port map (
            O => \N__12384\,
            I => \N__12378\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__12381\,
            I => \N__12375\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__12378\,
            I => \N__12372\
        );

    \I__1374\ : Span12Mux_s11_v
    port map (
            O => \N__12375\,
            I => \N__12367\
        );

    \I__1373\ : Span12Mux_h
    port map (
            O => \N__12372\,
            I => \N__12367\
        );

    \I__1372\ : Odrv12
    port map (
            O => \N__12367\,
            I => throttle_command_3
        );

    \I__1371\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12361\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__12361\,
            I => \N__12358\
        );

    \I__1369\ : Span4Mux_v
    port map (
            O => \N__12358\,
            I => \N__12355\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__12355\,
            I => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\
        );

    \I__1367\ : InMux
    port map (
            O => \N__12352\,
            I => \ppm_encoder_1.un1_throttle_cry_2\
        );

    \I__1366\ : InMux
    port map (
            O => \N__12349\,
            I => \ppm_encoder_1.un1_throttle_cry_3\
        );

    \I__1365\ : InMux
    port map (
            O => \N__12346\,
            I => \ppm_encoder_1.un1_throttle_cry_4\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__12343\,
            I => \N__12339\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__12342\,
            I => \N__12336\
        );

    \I__1362\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12333\
        );

    \I__1361\ : InMux
    port map (
            O => \N__12336\,
            I => \N__12330\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__12333\,
            I => alt_command_3
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__12330\,
            I => alt_command_3
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__12325\,
            I => \N__12321\
        );

    \I__1357\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12318\
        );

    \I__1356\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12315\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__12318\,
            I => alt_command_1
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__12315\,
            I => alt_command_1
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__12310\,
            I => \Commands_frame_decoder.source_CH1data8lto7Z0Z_1_cascade_\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__12307\,
            I => \Commands_frame_decoder.source_CH1data8_cascade_\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__12304\,
            I => \N__12300\
        );

    \I__1350\ : InMux
    port map (
            O => \N__12303\,
            I => \N__12297\
        );

    \I__1349\ : InMux
    port map (
            O => \N__12300\,
            I => \N__12294\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__12297\,
            I => alt_command_0
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__12294\,
            I => alt_command_0
        );

    \I__1346\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12280\
        );

    \I__1345\ : InMux
    port map (
            O => \N__12288\,
            I => \N__12280\
        );

    \I__1344\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12280\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__12280\,
            I => \Commands_frame_decoder.source_CH1data8\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__12277\,
            I => \N__12274\
        );

    \I__1341\ : InMux
    port map (
            O => \N__12274\,
            I => \N__12270\
        );

    \I__1340\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12267\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__12270\,
            I => \N__12264\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__12267\,
            I => alt_command_2
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__12264\,
            I => alt_command_2
        );

    \I__1336\ : InMux
    port map (
            O => \N__12259\,
            I => \N__12256\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__12256\,
            I => \Commands_frame_decoder.source_CH1data8lt7_0\
        );

    \I__1334\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12250\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__12250\,
            I => \dron_frame_decoder_1.drone_altitude_8\
        );

    \I__1332\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12244\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__12244\,
            I => drone_altitude_i_8
        );

    \I__1330\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12238\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__12238\,
            I => \dron_frame_decoder_1.drone_altitude_6\
        );

    \I__1328\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12232\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__12232\,
            I => drone_altitude_i_6
        );

    \I__1326\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12226\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__12226\,
            I => drone_altitude_1
        );

    \I__1324\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12220\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__12220\,
            I => \pid_alt.error_axbZ0Z_1\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__12217\,
            I => \dron_frame_decoder_1.source_Altitude8lto3Z0Z_0_cascade_\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__12214\,
            I => \dron_frame_decoder_1.source_Altitude8lt7_0_cascade_\
        );

    \I__1320\ : InMux
    port map (
            O => \N__12211\,
            I => \N__12208\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__12208\,
            I => drone_altitude_2
        );

    \I__1318\ : InMux
    port map (
            O => \N__12205\,
            I => \N__12202\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__12202\,
            I => \pid_alt.error_axbZ0Z_2\
        );

    \I__1316\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12188\
        );

    \I__1315\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12188\
        );

    \I__1314\ : InMux
    port map (
            O => \N__12197\,
            I => \N__12188\
        );

    \I__1313\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12183\
        );

    \I__1312\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12183\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__12188\,
            I => \dron_frame_decoder_1.source_Altitude8lt7_0\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__12183\,
            I => \dron_frame_decoder_1.source_Altitude8lt7_0\
        );

    \I__1309\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12175\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__12175\,
            I => drone_altitude_3
        );

    \I__1307\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12169\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__12169\,
            I => \pid_alt.error_axbZ0Z_3\
        );

    \I__1305\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12163\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__12163\,
            I => \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__12160\,
            I => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10_cascade_\
        );

    \I__1302\ : InMux
    port map (
            O => \N__12157\,
            I => \N__12154\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__12154\,
            I => \dron_frame_decoder_1.WDT10lto13_1\
        );

    \I__1300\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12148\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__12148\,
            I => \dron_frame_decoder_1.WDT10lt14_0\
        );

    \I__1298\ : InMux
    port map (
            O => \N__12145\,
            I => \N__12140\
        );

    \I__1297\ : InMux
    port map (
            O => \N__12144\,
            I => \N__12137\
        );

    \I__1296\ : InMux
    port map (
            O => \N__12143\,
            I => \N__12134\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__12140\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__12137\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__12134\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__12127\,
            I => \dron_frame_decoder_1.WDT10lt14_0_cascade_\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__12124\,
            I => \N__12120\
        );

    \I__1290\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12116\
        );

    \I__1289\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12111\
        );

    \I__1288\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12111\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__12116\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__12111\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__12106\,
            I => \N__12102\
        );

    \I__1284\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12099\
        );

    \I__1283\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12096\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__12099\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__12096\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__1280\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12088\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__12088\,
            I => \N__12085\
        );

    \I__1278\ : Span4Mux_s2_h
    port map (
            O => \N__12085\,
            I => \N__12081\
        );

    \I__1277\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12078\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__12081\,
            I => drone_altitude_0
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__12078\,
            I => drone_altitude_0
        );

    \I__1274\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12069\
        );

    \I__1273\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12066\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__12069\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__12066\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__1270\ : InMux
    port map (
            O => \N__12061\,
            I => \N__12058\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__12058\,
            I => \dron_frame_decoder_1.drone_altitude_4\
        );

    \I__1268\ : InMux
    port map (
            O => \N__12055\,
            I => \N__12052\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__12052\,
            I => drone_altitude_i_4
        );

    \I__1266\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12046\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__12046\,
            I => \dron_frame_decoder_1.drone_altitude_5\
        );

    \I__1264\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12040\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__12040\,
            I => drone_altitude_i_5
        );

    \I__1262\ : InMux
    port map (
            O => \N__12037\,
            I => \N__12034\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__12034\,
            I => \N__12030\
        );

    \I__1260\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12027\
        );

    \I__1259\ : Span4Mux_s2_h
    port map (
            O => \N__12030\,
            I => \N__12024\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__12027\,
            I => alt_kp_3
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__12024\,
            I => alt_kp_3
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__12019\,
            I => \N__12015\
        );

    \I__1255\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12012\
        );

    \I__1254\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12009\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__12012\,
            I => \N__12006\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__12009\,
            I => alt_kp_6
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__12006\,
            I => alt_kp_6
        );

    \I__1250\ : SRMux
    port map (
            O => \N__12001\,
            I => \N__11997\
        );

    \I__1249\ : SRMux
    port map (
            O => \N__12000\,
            I => \N__11994\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__11997\,
            I => \N__11991\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__11994\,
            I => \N__11988\
        );

    \I__1246\ : Span4Mux_s2_h
    port map (
            O => \N__11991\,
            I => \N__11985\
        );

    \I__1245\ : Span4Mux_s2_h
    port map (
            O => \N__11988\,
            I => \N__11982\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__11985\,
            I => \N__11979\
        );

    \I__1243\ : Span4Mux_h
    port map (
            O => \N__11982\,
            I => \N__11976\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__11979\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__11976\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__1240\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11967\
        );

    \I__1239\ : InMux
    port map (
            O => \N__11970\,
            I => \N__11964\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__11967\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__11964\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__1236\ : InMux
    port map (
            O => \N__11959\,
            I => \N__11955\
        );

    \I__1235\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11952\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__11955\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__11952\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__1232\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11943\
        );

    \I__1231\ : InMux
    port map (
            O => \N__11946\,
            I => \N__11940\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__11943\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__11940\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__11935\,
            I => \N__11931\
        );

    \I__1227\ : InMux
    port map (
            O => \N__11934\,
            I => \N__11928\
        );

    \I__1226\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11925\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__11928\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__11925\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__1223\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11916\
        );

    \I__1222\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11913\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__11916\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__11913\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__1219\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11903\
        );

    \I__1218\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11898\
        );

    \I__1217\ : InMux
    port map (
            O => \N__11906\,
            I => \N__11898\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__11903\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__11898\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__1214\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11889\
        );

    \I__1213\ : InMux
    port map (
            O => \N__11892\,
            I => \N__11886\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__11889\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__11886\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__11881\,
            I => \N__11877\
        );

    \I__1209\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11874\
        );

    \I__1208\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11871\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__11874\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__11871\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__1205\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11861\
        );

    \I__1204\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11856\
        );

    \I__1203\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11856\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__11861\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__11856\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__1200\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11847\
        );

    \I__1199\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11844\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__11847\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__11844\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__1196\ : InMux
    port map (
            O => \N__11839\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13\
        );

    \I__1195\ : InMux
    port map (
            O => \N__11836\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_14\
        );

    \I__1194\ : InMux
    port map (
            O => \N__11833\,
            I => \bfn_1_30_0_\
        );

    \I__1193\ : InMux
    port map (
            O => \N__11830\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_16\
        );

    \I__1192\ : InMux
    port map (
            O => \N__11827\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_17\
        );

    \I__1191\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11821\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__11821\,
            I => \N__11817\
        );

    \I__1189\ : InMux
    port map (
            O => \N__11820\,
            I => \N__11814\
        );

    \I__1188\ : Span4Mux_s2_h
    port map (
            O => \N__11817\,
            I => \N__11811\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__11814\,
            I => alt_kp_0
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__11811\,
            I => alt_kp_0
        );

    \I__1185\ : InMux
    port map (
            O => \N__11806\,
            I => \N__11802\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__11805\,
            I => \N__11799\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__11802\,
            I => \N__11796\
        );

    \I__1182\ : InMux
    port map (
            O => \N__11799\,
            I => \N__11793\
        );

    \I__1181\ : Span4Mux_s2_h
    port map (
            O => \N__11796\,
            I => \N__11790\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__11793\,
            I => alt_kp_2
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__11790\,
            I => alt_kp_2
        );

    \I__1178\ : InMux
    port map (
            O => \N__11785\,
            I => \N__11782\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__11782\,
            I => \N__11778\
        );

    \I__1176\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11775\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__11778\,
            I => \N__11772\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__11775\,
            I => alt_kp_1
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__11772\,
            I => alt_kp_1
        );

    \I__1172\ : CEMux
    port map (
            O => \N__11767\,
            I => \N__11763\
        );

    \I__1171\ : CEMux
    port map (
            O => \N__11766\,
            I => \N__11760\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__11763\,
            I => \N__11755\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__11760\,
            I => \N__11752\
        );

    \I__1168\ : CEMux
    port map (
            O => \N__11759\,
            I => \N__11749\
        );

    \I__1167\ : CEMux
    port map (
            O => \N__11758\,
            I => \N__11746\
        );

    \I__1166\ : Span4Mux_s3_h
    port map (
            O => \N__11755\,
            I => \N__11743\
        );

    \I__1165\ : Span4Mux_s3_h
    port map (
            O => \N__11752\,
            I => \N__11740\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__11749\,
            I => \N__11737\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__11746\,
            I => \N__11734\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__11743\,
            I => \pid_alt.source_p_enZ0\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__11740\,
            I => \pid_alt.source_p_enZ0\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__11737\,
            I => \pid_alt.source_p_enZ0\
        );

    \I__1159\ : Odrv12
    port map (
            O => \N__11734\,
            I => \pid_alt.source_p_enZ0\
        );

    \I__1158\ : InMux
    port map (
            O => \N__11725\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_4\
        );

    \I__1157\ : InMux
    port map (
            O => \N__11722\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_5\
        );

    \I__1156\ : InMux
    port map (
            O => \N__11719\,
            I => \N__11716\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__11716\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_7\
        );

    \I__1154\ : InMux
    port map (
            O => \N__11713\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_6\
        );

    \I__1153\ : InMux
    port map (
            O => \N__11710\,
            I => \bfn_1_29_0_\
        );

    \I__1152\ : InMux
    port map (
            O => \N__11707\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_8\
        );

    \I__1151\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11701\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__11701\,
            I => \N__11698\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__11698\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_10\
        );

    \I__1148\ : InMux
    port map (
            O => \N__11695\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_9\
        );

    \I__1147\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11689\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__11689\,
            I => \N__11686\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__11686\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_11\
        );

    \I__1144\ : InMux
    port map (
            O => \N__11683\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_10\
        );

    \I__1143\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11677\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__11677\,
            I => \N__11674\
        );

    \I__1141\ : Span4Mux_v
    port map (
            O => \N__11674\,
            I => \N__11671\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__11671\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_12\
        );

    \I__1139\ : InMux
    port map (
            O => \N__11668\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_11\
        );

    \I__1138\ : InMux
    port map (
            O => \N__11665\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_12\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__1136\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11656\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__11656\,
            I => \N__11653\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__11653\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\
        );

    \I__1133\ : InMux
    port map (
            O => \N__11650\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_0\
        );

    \I__1132\ : InMux
    port map (
            O => \N__11647\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_1\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__11644\,
            I => \N__11641\
        );

    \I__1130\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11638\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__11638\,
            I => \N__11635\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__11635\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_3\
        );

    \I__1127\ : InMux
    port map (
            O => \N__11632\,
            I => \N__11629\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__11629\,
            I => \N__11626\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__11626\,
            I => \ppm_encoder_1.un1_init_pulses_11_3\
        );

    \I__1124\ : InMux
    port map (
            O => \N__11623\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_2\
        );

    \I__1123\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11617\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__11617\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_4\
        );

    \I__1121\ : InMux
    port map (
            O => \N__11614\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_3\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__11611\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__11608\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__11605\,
            I => \N__11601\
        );

    \I__1117\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11596\
        );

    \I__1116\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11596\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__11596\,
            I => \N__11593\
        );

    \I__1114\ : Odrv12
    port map (
            O => \N__11593\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__1113\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11587\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__11587\,
            I => \ppm_encoder_1.un2_throttle_iv_1_6\
        );

    \I__1111\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11579\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__11583\,
            I => \N__11576\
        );

    \I__1109\ : InMux
    port map (
            O => \N__11582\,
            I => \N__11573\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__11579\,
            I => \N__11570\
        );

    \I__1107\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11567\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__11573\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__11570\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__11567\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__1103\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11557\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__11557\,
            I => \N__11552\
        );

    \I__1101\ : InMux
    port map (
            O => \N__11556\,
            I => \N__11547\
        );

    \I__1100\ : InMux
    port map (
            O => \N__11555\,
            I => \N__11547\
        );

    \I__1099\ : Odrv12
    port map (
            O => \N__11552\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__11547\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__11542\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \ppm_encoder_1.un2_throttle_iv_1_13_cascade_\
        );

    \I__1095\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11533\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__11533\,
            I => \ppm_encoder_1.un2_throttle_iv_0_13\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__11530\,
            I => \N__11525\
        );

    \I__1092\ : InMux
    port map (
            O => \N__11529\,
            I => \N__11522\
        );

    \I__1091\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11519\
        );

    \I__1090\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11516\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__11522\,
            I => \N__11511\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__11519\,
            I => \N__11511\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__11516\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__1086\ : Odrv12
    port map (
            O => \N__11511\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__11506\,
            I => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\
        );

    \I__1084\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11500\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__11500\,
            I => \N__11497\
        );

    \I__1082\ : Odrv12
    port map (
            O => \N__11497\,
            I => drone_altitude_i_7
        );

    \I__1081\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11491\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__11491\,
            I => \dron_frame_decoder_1.drone_altitude_7\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__11488\,
            I => \ppm_encoder_1.N_297_cascade_\
        );

    \I__1078\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11482\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__11482\,
            I => \dron_frame_decoder_1.drone_altitude_11\
        );

    \I__1076\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11476\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__11476\,
            I => \pid_alt.error_axbZ0Z_12\
        );

    \I__1074\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11470\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__11470\,
            I => drone_altitude_12
        );

    \I__1072\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__11464\,
            I => \pid_alt.error_axbZ0Z_13\
        );

    \I__1070\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11458\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__11458\,
            I => drone_altitude_13
        );

    \I__1068\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11452\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__11452\,
            I => \N__11449\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__11449\,
            I => \pid_alt.error_axbZ0Z_14\
        );

    \I__1065\ : InMux
    port map (
            O => \N__11446\,
            I => \N__11443\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__11443\,
            I => \N__11440\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__11440\,
            I => drone_altitude_15
        );

    \I__1062\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__11434\,
            I => \N__11431\
        );

    \I__1060\ : Span4Mux_s1_h
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__11428\,
            I => \pid_alt.error_10\
        );

    \I__1058\ : InMux
    port map (
            O => \N__11425\,
            I => \pid_alt.error_cry_9\
        );

    \I__1057\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11419\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11416\
        );

    \I__1055\ : Span4Mux_s1_h
    port map (
            O => \N__11416\,
            I => \N__11413\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__11413\,
            I => \pid_alt.error_11\
        );

    \I__1053\ : InMux
    port map (
            O => \N__11410\,
            I => \pid_alt.error_cry_10\
        );

    \I__1052\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11404\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__11404\,
            I => \N__11401\
        );

    \I__1050\ : Span4Mux_s1_h
    port map (
            O => \N__11401\,
            I => \N__11398\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__11398\,
            I => \pid_alt.error_12\
        );

    \I__1048\ : InMux
    port map (
            O => \N__11395\,
            I => \pid_alt.error_cry_11\
        );

    \I__1047\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11389\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__11389\,
            I => \N__11386\
        );

    \I__1045\ : Span4Mux_s1_h
    port map (
            O => \N__11386\,
            I => \N__11383\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__11383\,
            I => \pid_alt.error_13\
        );

    \I__1043\ : InMux
    port map (
            O => \N__11380\,
            I => \pid_alt.error_cry_12\
        );

    \I__1042\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11374\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__11374\,
            I => \N__11371\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__11371\,
            I => \N__11368\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__11368\,
            I => \pid_alt.error_14\
        );

    \I__1038\ : InMux
    port map (
            O => \N__11365\,
            I => \pid_alt.error_cry_13\
        );

    \I__1037\ : InMux
    port map (
            O => \N__11362\,
            I => \pid_alt.error_cry_14\
        );

    \I__1036\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11356\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__11356\,
            I => \N__11353\
        );

    \I__1034\ : Span4Mux_v
    port map (
            O => \N__11353\,
            I => \N__11350\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__11350\,
            I => \pid_alt.error_15\
        );

    \I__1032\ : InMux
    port map (
            O => \N__11347\,
            I => \N__11344\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__11344\,
            I => drone_altitude_i_10
        );

    \I__1030\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11338\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__11338\,
            I => \dron_frame_decoder_1.drone_altitude_10\
        );

    \I__1028\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11332\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__11332\,
            I => drone_altitude_i_11
        );

    \I__1026\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11326\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11323\
        );

    \I__1024\ : Span4Mux_s1_h
    port map (
            O => \N__11323\,
            I => \N__11320\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__11320\,
            I => \pid_alt.error_2\
        );

    \I__1022\ : InMux
    port map (
            O => \N__11317\,
            I => \pid_alt.error_cry_1\
        );

    \I__1021\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11311\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__11311\,
            I => \N__11308\
        );

    \I__1019\ : Span4Mux_s1_h
    port map (
            O => \N__11308\,
            I => \N__11305\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__11305\,
            I => \pid_alt.error_3\
        );

    \I__1017\ : InMux
    port map (
            O => \N__11302\,
            I => \pid_alt.error_cry_2\
        );

    \I__1016\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11296\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__1014\ : Span4Mux_v
    port map (
            O => \N__11293\,
            I => \N__11290\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__11290\,
            I => \pid_alt.error_4\
        );

    \I__1012\ : InMux
    port map (
            O => \N__11287\,
            I => \pid_alt.error_cry_3\
        );

    \I__1011\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__11278\,
            I => \pid_alt.error_5\
        );

    \I__1008\ : InMux
    port map (
            O => \N__11275\,
            I => \pid_alt.error_cry_4\
        );

    \I__1007\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__1005\ : Span4Mux_s1_h
    port map (
            O => \N__11266\,
            I => \N__11263\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__11263\,
            I => \pid_alt.error_6\
        );

    \I__1003\ : InMux
    port map (
            O => \N__11260\,
            I => \pid_alt.error_cry_5\
        );

    \I__1002\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11254\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__11254\,
            I => \N__11251\
        );

    \I__1000\ : Span4Mux_s1_h
    port map (
            O => \N__11251\,
            I => \N__11248\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__11248\,
            I => \pid_alt.error_7\
        );

    \I__998\ : InMux
    port map (
            O => \N__11245\,
            I => \pid_alt.error_cry_6\
        );

    \I__997\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11239\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__11239\,
            I => \N__11236\
        );

    \I__995\ : Span4Mux_s2_h
    port map (
            O => \N__11236\,
            I => \N__11233\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__11233\,
            I => \pid_alt.error_8\
        );

    \I__993\ : InMux
    port map (
            O => \N__11230\,
            I => \bfn_1_16_0_\
        );

    \I__992\ : InMux
    port map (
            O => \N__11227\,
            I => \N__11224\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__11224\,
            I => \N__11221\
        );

    \I__990\ : Span4Mux_v
    port map (
            O => \N__11221\,
            I => \N__11218\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__11218\,
            I => \pid_alt.error_9\
        );

    \I__988\ : InMux
    port map (
            O => \N__11215\,
            I => \pid_alt.error_cry_8\
        );

    \I__987\ : InMux
    port map (
            O => \N__11212\,
            I => \bfn_1_14_0_\
        );

    \I__986\ : InMux
    port map (
            O => \N__11209\,
            I => \dron_frame_decoder_1.un1_WDT_cry_8\
        );

    \I__985\ : InMux
    port map (
            O => \N__11206\,
            I => \dron_frame_decoder_1.un1_WDT_cry_9\
        );

    \I__984\ : InMux
    port map (
            O => \N__11203\,
            I => \dron_frame_decoder_1.un1_WDT_cry_10\
        );

    \I__983\ : InMux
    port map (
            O => \N__11200\,
            I => \dron_frame_decoder_1.un1_WDT_cry_11\
        );

    \I__982\ : InMux
    port map (
            O => \N__11197\,
            I => \dron_frame_decoder_1.un1_WDT_cry_12\
        );

    \I__981\ : InMux
    port map (
            O => \N__11194\,
            I => \dron_frame_decoder_1.un1_WDT_cry_13\
        );

    \I__980\ : InMux
    port map (
            O => \N__11191\,
            I => \dron_frame_decoder_1.un1_WDT_cry_14\
        );

    \I__979\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11185\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__11185\,
            I => \N__11182\
        );

    \I__977\ : Span4Mux_s1_h
    port map (
            O => \N__11182\,
            I => \N__11179\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__11179\,
            I => \pid_alt.error_1\
        );

    \I__975\ : InMux
    port map (
            O => \N__11176\,
            I => \pid_alt.error_cry_0\
        );

    \I__974\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__11170\,
            I => \dron_frame_decoder_1.WDTZ0Z_0\
        );

    \I__972\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11164\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__11164\,
            I => \dron_frame_decoder_1.WDTZ0Z_1\
        );

    \I__970\ : InMux
    port map (
            O => \N__11161\,
            I => \dron_frame_decoder_1.un1_WDT_cry_0\
        );

    \I__969\ : InMux
    port map (
            O => \N__11158\,
            I => \N__11155\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__11155\,
            I => \dron_frame_decoder_1.WDTZ0Z_2\
        );

    \I__967\ : InMux
    port map (
            O => \N__11152\,
            I => \dron_frame_decoder_1.un1_WDT_cry_1\
        );

    \I__966\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11146\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__11146\,
            I => \dron_frame_decoder_1.WDTZ0Z_3\
        );

    \I__964\ : InMux
    port map (
            O => \N__11143\,
            I => \dron_frame_decoder_1.un1_WDT_cry_2\
        );

    \I__963\ : InMux
    port map (
            O => \N__11140\,
            I => \dron_frame_decoder_1.un1_WDT_cry_3\
        );

    \I__962\ : InMux
    port map (
            O => \N__11137\,
            I => \dron_frame_decoder_1.un1_WDT_cry_4\
        );

    \I__961\ : InMux
    port map (
            O => \N__11134\,
            I => \dron_frame_decoder_1.un1_WDT_cry_5\
        );

    \I__960\ : InMux
    port map (
            O => \N__11131\,
            I => \dron_frame_decoder_1.un1_WDT_cry_6\
        );

    \I__959\ : InMux
    port map (
            O => \N__11128\,
            I => \N__11125\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__11125\,
            I => \pid_alt.O_11\
        );

    \I__957\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11119\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__11119\,
            I => \pid_alt.O_13\
        );

    \I__955\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11113\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__11113\,
            I => \N__11110\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__11110\,
            I => \pid_alt.O_18\
        );

    \I__952\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11104\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__11104\,
            I => \pid_alt.O_14\
        );

    \I__950\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11098\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__11098\,
            I => \pid_alt.O_4\
        );

    \I__948\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11092\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__11092\,
            I => \pid_alt.O_5\
        );

    \I__946\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11086\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__11086\,
            I => \pid_alt.O_9\
        );

    \I__944\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11080\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__11080\,
            I => \pid_alt.O_15\
        );

    \I__942\ : InMux
    port map (
            O => \N__11077\,
            I => \N__11074\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__11074\,
            I => \pid_alt.O_8\
        );

    \I__940\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11068\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__11068\,
            I => \N__11065\
        );

    \I__938\ : Odrv4
    port map (
            O => \N__11065\,
            I => \pid_alt.O_17\
        );

    \I__937\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11059\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__11059\,
            I => \pid_alt.O_6\
        );

    \I__935\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11053\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__11053\,
            I => \pid_alt.O_7\
        );

    \I__933\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11047\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__11047\,
            I => \N__11044\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__11044\,
            I => \pid_alt.O_10\
        );

    \I__930\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11038\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__11038\,
            I => \N__11035\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__11035\,
            I => \pid_alt.O_16\
        );

    \I__927\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11029\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__11029\,
            I => \pid_alt.O_12\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un3_source_data_0_cry_7\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un2_source_data_0_cry_8\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un3_source_data_0_cry_7\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un2_source_data_0_cry_8\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un3_source_data_0_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un2_source_data_0_cry_8\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_2_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_throttle_cry_7\,
            carryinitout => \bfn_2_20_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_rudder_cry_13\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_elevator_cry_13\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_aileron_cry_13\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_3_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_25_0_\
        );

    \IN_MUX_bfv_3_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            carryinitout => \bfn_3_26_0_\
        );

    \IN_MUX_bfv_3_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            carryinitout => \bfn_3_27_0_\
        );

    \IN_MUX_bfv_1_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_28_0_\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_1_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            carryinitout => \bfn_1_30_0_\
        );

    \IN_MUX_bfv_4_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_29_0_\
        );

    \IN_MUX_bfv_4_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.counter24_0_data_tmp_7\,
            carryinitout => \bfn_4_30_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.error_cry_7\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_5_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_19_0_\
        );

    \IN_MUX_bfv_7_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_28_0_\
        );

    \IN_MUX_bfv_7_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_7\,
            carryinitout => \bfn_7_29_0_\
        );

    \IN_MUX_bfv_7_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_15\,
            carryinitout => \bfn_7_30_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \dron_frame_decoder_1.un1_WDT_cry_7\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_4_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Commands_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_4_19_0_\
        );

    \reset_module_System.reset_RNITC69\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26679\,
            GLOBALBUFFEROUTPUT => reset_system_g
        );

    \pc_frame_decoder_dv_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26833\,
            GLOBALBUFFEROUTPUT => pc_frame_decoder_dv_0_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18883\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_168_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pid_alt.source_p_ess_13_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11071\,
            lcout => throttle_command_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29387\,
            ce => \N__11766\,
            sr => \N__28714\
        );

    \pid_alt.source_p_ess_2_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11062\,
            lcout => throttle_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29387\,
            ce => \N__11766\,
            sr => \N__28714\
        );

    \pid_alt.source_p_ess_3_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11056\,
            lcout => throttle_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29387\,
            ce => \N__11766\,
            sr => \N__28714\
        );

    \pid_alt.source_p_ess_6_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11050\,
            lcout => throttle_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29387\,
            ce => \N__11766\,
            sr => \N__28714\
        );

    \pid_alt.source_p_9_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28954\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11041\,
            lcout => throttle_command_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29386\,
            ce => \N__11758\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_5_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28951\,
            in2 => \_gnd_net_\,
            in3 => \N__11032\,
            lcout => throttle_command_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29386\,
            ce => \N__11758\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_4_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11128\,
            lcout => throttle_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29386\,
            ce => \N__11758\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_1_6_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28950\,
            in2 => \_gnd_net_\,
            in3 => \N__11122\,
            lcout => throttle_command_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29386\,
            ce => \N__11758\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_10_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11116\,
            lcout => throttle_command_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29386\,
            ce => \N__11758\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_7_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28956\,
            in2 => \_gnd_net_\,
            in3 => \N__11107\,
            lcout => throttle_command_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29384\,
            ce => \N__11759\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11101\,
            lcout => throttle_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29384\,
            ce => \N__11759\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_1_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28955\,
            in2 => \_gnd_net_\,
            in3 => \N__11095\,
            lcout => throttle_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29384\,
            ce => \N__11759\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_1_3_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__28959\,
            in1 => \N__11089\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => throttle_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29384\,
            ce => \N__11759\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28957\,
            in2 => \_gnd_net_\,
            in3 => \N__11083\,
            lcout => throttle_command_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29384\,
            ce => \N__11759\,
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_1_2_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28963\,
            in2 => \_gnd_net_\,
            in3 => \N__11077\,
            lcout => throttle_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29381\,
            ce => \N__11767\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_0_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11173\,
            in2 => \N__12106\,
            in3 => \N__12105\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_0\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_1_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11167\,
            in2 => \_gnd_net_\,
            in3 => \N__11161\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_0\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_1\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_2_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11158\,
            in2 => \_gnd_net_\,
            in3 => \N__11152\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_1\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_2\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_3_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11149\,
            in2 => \_gnd_net_\,
            in3 => \N__11143\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_2\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_3\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_4_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11920\,
            in2 => \_gnd_net_\,
            in3 => \N__11140\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_3\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_4\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_5_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11947\,
            in2 => \_gnd_net_\,
            in3 => \N__11137\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_4\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_5\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_6_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11971\,
            in2 => \_gnd_net_\,
            in3 => \N__11134\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_5\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_6\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_7_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11851\,
            in2 => \_gnd_net_\,
            in3 => \N__11131\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_6\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_7\,
            clk => \N__29378\,
            ce => 'H',
            sr => \N__12000\
        );

    \dron_frame_decoder_1.WDT_8_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11959\,
            in2 => \_gnd_net_\,
            in3 => \N__11212\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_8\,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \dron_frame_decoder_1.WDT_9_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11934\,
            in2 => \_gnd_net_\,
            in3 => \N__11209\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_8\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_9\,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \dron_frame_decoder_1.WDT_10_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11893\,
            in2 => \_gnd_net_\,
            in3 => \N__11206\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_9\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_10\,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \dron_frame_decoder_1.WDT_11_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11866\,
            in2 => \_gnd_net_\,
            in3 => \N__11203\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_10\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_11\,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \dron_frame_decoder_1.WDT_12_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11908\,
            in2 => \_gnd_net_\,
            in3 => \N__11200\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_11\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_12\,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \dron_frame_decoder_1.WDT_13_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11880\,
            in2 => \_gnd_net_\,
            in3 => \N__11197\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_12\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_13\,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \dron_frame_decoder_1.WDT_14_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12123\,
            in2 => \_gnd_net_\,
            in3 => \N__11194\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_13\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_14\,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \dron_frame_decoder_1.WDT_15_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12145\,
            in2 => \_gnd_net_\,
            in3 => \N__11191\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29375\,
            ce => 'H',
            sr => \N__12001\
        );

    \pid_alt.error_cry_0_c_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12072\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \pid_alt.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_RNI1N2F_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12223\,
            in2 => \_gnd_net_\,
            in3 => \N__11176\,
            lcout => \pid_alt.error_1\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_0\,
            carryout => \pid_alt.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_1_c_RNI3Q3F_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12205\,
            in2 => \_gnd_net_\,
            in3 => \N__11317\,
            lcout => \pid_alt.error_2\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_1\,
            carryout => \pid_alt.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_2_c_RNI5T4F_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12172\,
            in2 => \_gnd_net_\,
            in3 => \N__11302\,
            lcout => \pid_alt.error_3\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_2\,
            carryout => \pid_alt.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_3_c_RNIKE1T_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12055\,
            in2 => \N__12304\,
            in3 => \N__11287\,
            lcout => \pid_alt.error_4\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_3\,
            carryout => \pid_alt.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_4_c_RNINI2T_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12043\,
            in2 => \N__12325\,
            in3 => \N__11275\,
            lcout => \pid_alt.error_5\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_4\,
            carryout => \pid_alt.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_5_c_RNIQM3T_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12235\,
            in2 => \N__12277\,
            in3 => \N__11260\,
            lcout => \pid_alt.error_6\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_5\,
            carryout => \pid_alt.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_6_c_RNITQ4T_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11503\,
            in2 => \N__12342\,
            in3 => \N__11245\,
            lcout => \pid_alt.error_7\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_6\,
            carryout => \pid_alt.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_7_c_RNI9LEM_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12247\,
            in2 => \N__13327\,
            in3 => \N__11230\,
            lcout => \pid_alt.error_8\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pid_alt.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_8_c_RNICPFM_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12409\,
            in2 => \N__13315\,
            in3 => \N__11215\,
            lcout => \pid_alt.error_9\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_8\,
            carryout => \pid_alt.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_9_c_RNIMMUJ_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11347\,
            in2 => \N__13303\,
            in3 => \N__11425\,
            lcout => \pid_alt.error_10\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_9\,
            carryout => \pid_alt.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_10_c_RNI0SDO_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11335\,
            in2 => \N__13738\,
            in3 => \N__11410\,
            lcout => \pid_alt.error_11\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_10\,
            carryout => \pid_alt.error_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_11_c_RNI5JAH_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11479\,
            in2 => \_gnd_net_\,
            in3 => \N__11395\,
            lcout => \pid_alt.error_12\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_11\,
            carryout => \pid_alt.error_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_12_c_RNI7MBH_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11467\,
            in2 => \_gnd_net_\,
            in3 => \N__11380\,
            lcout => \pid_alt.error_13\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_12\,
            carryout => \pid_alt.error_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_13_c_RNI9PCH_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11455\,
            in2 => \_gnd_net_\,
            in3 => \N__11365\,
            lcout => \pid_alt.error_14\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_13\,
            carryout => \pid_alt.error_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_14_c_RNIBSDH_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11446\,
            in2 => \_gnd_net_\,
            in3 => \N__11362\,
            lcout => \pid_alt.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11341\,
            lcout => drone_altitude_i_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_10_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15289\,
            lcout => \dron_frame_decoder_1.drone_altitude_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29363\,
            ce => \N__13568\,
            sr => \N__28750\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11485\,
            lcout => drone_altitude_i_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_11_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15256\,
            lcout => \dron_frame_decoder_1.drone_altitude_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29363\,
            ce => \N__13568\,
            sr => \N__28750\
        );

    \pid_alt.error_axb_12_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11473\,
            lcout => \pid_alt.error_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_12_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15192\,
            lcout => drone_altitude_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29363\,
            ce => \N__13568\,
            sr => \N__28750\
        );

    \pid_alt.error_axb_13_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11461\,
            lcout => \pid_alt.error_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_13_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15132\,
            lcout => drone_altitude_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29363\,
            ce => \N__13568\,
            sr => \N__28750\
        );

    \pid_alt.error_axb_14_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12403\,
            lcout => \pid_alt.error_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_15_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15015\,
            lcout => drone_altitude_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29357\,
            ce => \N__13572\,
            sr => \N__28756\
        );

    \dron_frame_decoder_1.source_Altitude_esr_8_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14847\,
            lcout => \dron_frame_decoder_1.drone_altitude_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29357\,
            ce => \N__13572\,
            sr => \N__28756\
        );

    \ppm_encoder_1.throttle_6_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__12457\,
            in1 => \N__12478\,
            in2 => \N__11530\,
            in3 => \N__24864\,
            lcout => \ppm_encoder_1.throttleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29350\,
            ce => 'H',
            sr => \N__28763\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11494\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_7_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15014\,
            lcout => \dron_frame_decoder_1.drone_altitude_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29345\,
            ce => \N__13722\,
            sr => \N__28769\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22772\,
            in1 => \N__11529\,
            in2 => \_gnd_net_\,
            in3 => \N__11560\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20959\,
            in2 => \N__11488\,
            in3 => \N__11584\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22761\,
            in1 => \N__13866\,
            in2 => \_gnd_net_\,
            in3 => \N__19801\,
            lcout => \ppm_encoder_1.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__22762\,
            in1 => \N__28964\,
            in2 => \N__20980\,
            in3 => \N__23732\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110110"
        )
    port map (
            in0 => \N__23731\,
            in1 => \N__17818\,
            in2 => \N__28979\,
            in3 => \N__20773\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__18562\,
            in1 => \N__28968\,
            in2 => \N__20979\,
            in3 => \N__23617\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18561\,
            in1 => \N__17801\,
            in2 => \N__20572\,
            in3 => \N__17857\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_158_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__16150\,
            in1 => \N__23613\,
            in2 => \_gnd_net_\,
            in3 => \N__20782\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010101010"
        )
    port map (
            in0 => \N__17858\,
            in1 => \N__22798\,
            in2 => \N__20972\,
            in3 => \N__20568\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20067\,
            in1 => \N__23612\,
            in2 => \_gnd_net_\,
            in3 => \N__20781\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_12_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20783\,
            in1 => \_gnd_net_\,
            in2 => \N__23724\,
            in3 => \N__20066\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI47DH2_13_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__15965\,
            in1 => \N__25006\,
            in2 => \N__16054\,
            in3 => \N__20095\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIKVRT5_13_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__16351\,
            in1 => \_gnd_net_\,
            in2 => \N__11539\,
            in3 => \N__11536\,
            lcout => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIK8JI2_13_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100110001"
        )
    port map (
            in0 => \N__15845\,
            in1 => \N__15726\,
            in2 => \N__20136\,
            in3 => \N__21016\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIO1KK2_6_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__11528\,
            in1 => \N__21072\,
            in2 => \N__15745\,
            in3 => \N__15844\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIEDI96_6_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18361\,
            in2 => \N__11506\,
            in3 => \N__11590\,
            lcout => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI8GVN2_6_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__11555\,
            in1 => \N__15964\,
            in2 => \N__11583\,
            in3 => \N__16031\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_6_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__11582\,
            in1 => \N__24954\,
            in2 => \_gnd_net_\,
            in3 => \N__24172\,
            lcout => \ppm_encoder_1.aileronZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29314\,
            ce => 'H',
            sr => \N__28782\
        );

    \ppm_encoder_1.elevator_6_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__11556\,
            in1 => \N__24955\,
            in2 => \_gnd_net_\,
            in3 => \N__25996\,
            lcout => \ppm_encoder_1.elevatorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29314\,
            ce => 'H',
            sr => \N__28782\
        );

    \ppm_encoder_1.init_pulses_3_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18250\,
            in1 => \N__11632\,
            in2 => \N__18062\,
            in3 => \N__14041\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29306\,
            ce => 'H',
            sr => \N__28786\
        );

    \ppm_encoder_1.throttle_RNIT9352_3_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101001100101"
        )
    port map (
            in0 => \N__18461\,
            in1 => \N__18629\,
            in2 => \N__15865\,
            in3 => \N__16443\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI82223_3_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11542\,
            in3 => \N__14064\,
            lcout => \ppm_encoder_1.throttle_RNI82223Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__18460\,
            in1 => \N__23601\,
            in2 => \_gnd_net_\,
            in3 => \N__20685\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20686\,
            in1 => \_gnd_net_\,
            in2 => \N__23702\,
            in3 => \N__18462\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_3_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__12385\,
            in1 => \N__12364\,
            in2 => \N__24967\,
            in3 => \N__18630\,
            lcout => \ppm_encoder_1.throttleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29306\,
            ce => 'H',
            sr => \N__28786\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__16149\,
            in1 => \N__23653\,
            in2 => \_gnd_net_\,
            in3 => \N__20702\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17842\,
            in2 => \_gnd_net_\,
            in3 => \N__12867\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16313\,
            in2 => \N__11611\,
            in3 => \N__12789\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__23652\,
            in1 => \_gnd_net_\,
            in2 => \N__11608\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__23849\,
            in1 => \N__13113\,
            in2 => \_gnd_net_\,
            in3 => \N__23654\,
            lcout => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23655\,
            in1 => \N__28962\,
            in2 => \N__11605\,
            in3 => \N__17843\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__28961\,
            in1 => \N__11604\,
            in2 => \N__12829\,
            in3 => \N__23657\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23656\,
            in1 => \N__26697\,
            in2 => \N__20593\,
            in3 => \N__12868\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__20554\,
            in1 => \N__18676\,
            in2 => \N__20381\,
            in3 => \N__12774\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_4_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24481\,
            lcout => \ppm_encoder_1.rudderZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29288\,
            ce => \N__25065\,
            sr => \N__28792\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__18675\,
            in1 => \N__23763\,
            in2 => \_gnd_net_\,
            in3 => \N__20689\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20690\,
            in1 => \_gnd_net_\,
            in2 => \N__23810\,
            in3 => \N__20439\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20438\,
            in1 => \N__23767\,
            in2 => \_gnd_net_\,
            in3 => \N__20691\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20692\,
            in1 => \_gnd_net_\,
            in2 => \N__23811\,
            in3 => \N__16194\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__16195\,
            in1 => \N__23771\,
            in2 => \_gnd_net_\,
            in3 => \N__20693\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13012\,
            in2 => \N__11662\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_28_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_1_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16225\,
            in2 => \_gnd_net_\,
            in3 => \N__11650\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_2_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13081\,
            in2 => \N__12940\,
            in3 => \N__11647\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_3_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11644\,
            in3 => \N__11623\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_4_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11620\,
            in2 => \_gnd_net_\,
            in3 => \N__11614\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_5_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17731\,
            in2 => \_gnd_net_\,
            in3 => \N__11725\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_6_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12880\,
            in2 => \N__12952\,
            in3 => \N__11722\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_7_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11719\,
            in2 => \_gnd_net_\,
            in3 => \N__11713\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_8_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13048\,
            in2 => \_gnd_net_\,
            in3 => \N__11710\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_8\,
            ltout => OPEN,
            carryin => \bfn_1_29_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_9_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13228\,
            in2 => \_gnd_net_\,
            in3 => \N__11707\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_10_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11704\,
            in2 => \_gnd_net_\,
            in3 => \N__11695\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_11_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11692\,
            in2 => \_gnd_net_\,
            in3 => \N__11683\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_12_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11680\,
            in2 => \_gnd_net_\,
            in3 => \N__11668\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_13_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13141\,
            in2 => \N__12961\,
            in3 => \N__11665\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_14_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18277\,
            in2 => \_gnd_net_\,
            in3 => \N__11839\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_15_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16471\,
            in2 => \_gnd_net_\,
            in3 => \N__11836\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_16_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18265\,
            in3 => \N__11833\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_16\,
            ltout => OPEN,
            carryin => \bfn_1_30_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_17_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13066\,
            in3 => \N__11830\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_18_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__23780\,
            in1 => \N__17565\,
            in2 => \N__20807\,
            in3 => \N__11827\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset1data_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__28941\,
            in1 => \N__11820\,
            in2 => \N__16676\,
            in3 => \N__29846\,
            lcout => alt_kp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset1data_2_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__28355\,
            in1 => \N__16672\,
            in2 => \N__11805\,
            in3 => \N__28944\,
            lcout => alt_kp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset1data_1_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__28942\,
            in1 => \N__11781\,
            in2 => \N__16677\,
            in3 => \N__27767\,
            lcout => alt_kp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_p_en_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13836\,
            in2 => \_gnd_net_\,
            in3 => \N__28940\,
            lcout => \pid_alt.source_p_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset1data_3_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__28943\,
            in1 => \N__12033\,
            in2 => \N__16678\,
            in3 => \N__28113\,
            lcout => alt_kp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset1data_5_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__28230\,
            in1 => \N__16665\,
            in2 => \N__12019\,
            in3 => \N__28978\,
            lcout => alt_kp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_1_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__13147\,
            in1 => \N__13680\,
            in2 => \N__13258\,
            in3 => \N__13351\,
            lcout => \dron_frame_decoder_1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29379\,
            ce => 'H',
            sr => \N__28720\
        );

    \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13464\,
            in2 => \_gnd_net_\,
            in3 => \N__28932\,
            lcout => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__12151\,
            in1 => \N__12144\,
            in2 => \N__12124\,
            in3 => \N__13468\,
            lcout => \dron_frame_decoder_1.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11906\,
            in1 => \N__11864\,
            in2 => \_gnd_net_\,
            in3 => \N__11970\,
            lcout => \dron_frame_decoder_1.WDT10lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11958\,
            in1 => \N__11946\,
            in2 => \N__11935\,
            in3 => \N__11919\,
            lcout => \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__11907\,
            in1 => \N__11892\,
            in2 => \N__11881\,
            in3 => \N__11865\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__11850\,
            in1 => \N__12166\,
            in2 => \N__12160\,
            in3 => \N__12157\,
            lcout => \dron_frame_decoder_1.WDT10lt14_0\,
            ltout => \dron_frame_decoder_1.WDT10lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12143\,
            in2 => \N__12127\,
            in3 => \N__12119\,
            lcout => \dron_frame_decoder_1.WDT10_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12197\,
            in1 => \N__15011\,
            in2 => \N__14848\,
            in3 => \N__15088\,
            lcout => drone_altitude_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__13721\,
            sr => \N__28730\
        );

    \pid_alt.error_cry_0_c_inv_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__12073\,
            in1 => \N__27273\,
            in2 => \_gnd_net_\,
            in3 => \N__12084\,
            lcout => \pid_alt.drone_altitude_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_4_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12198\,
            in1 => \N__15087\,
            in2 => \N__15199\,
            in3 => \N__15013\,
            lcout => \dron_frame_decoder_1.drone_altitude_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__13721\,
            sr => \N__28730\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12061\,
            lcout => drone_altitude_i_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_5_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12199\,
            in1 => \N__15012\,
            in2 => \N__15136\,
            in3 => \N__15089\,
            lcout => \dron_frame_decoder_1.drone_altitude_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__13721\,
            sr => \N__28730\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12049\,
            lcout => drone_altitude_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_6_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15090\,
            lcout => \dron_frame_decoder_1.drone_altitude_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__13721\,
            sr => \N__28730\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12241\,
            lcout => drone_altitude_i_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_1_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12195\,
            in1 => \N__15006\,
            in2 => \N__14815\,
            in3 => \N__15084\,
            lcout => drone_altitude_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29369\,
            ce => \N__13726\,
            sr => \N__28734\
        );

    \pid_alt.error_axb_1_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12229\,
            lcout => \pid_alt.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude8lto3_0_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15254\,
            in2 => \_gnd_net_\,
            in3 => \N__15287\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.source_Altitude8lto3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude8lto5_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__15125\,
            in1 => \N__14810\,
            in2 => \N__12217\,
            in3 => \N__15191\,
            lcout => \dron_frame_decoder_1.source_Altitude8lt7_0\,
            ltout => \dron_frame_decoder_1.source_Altitude8lt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_2_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__15086\,
            in1 => \N__15007\,
            in2 => \N__12214\,
            in3 => \N__15288\,
            lcout => drone_altitude_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29369\,
            ce => \N__13726\,
            sr => \N__28734\
        );

    \pid_alt.error_axb_2_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12211\,
            lcout => \pid_alt.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_3_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__12196\,
            in1 => \N__15255\,
            in2 => \N__15016\,
            in3 => \N__15085\,
            lcout => drone_altitude_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29369\,
            ce => \N__13726\,
            sr => \N__28734\
        );

    \pid_alt.error_axb_3_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12178\,
            lcout => \pid_alt.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_3_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__12289\,
            in1 => \N__16894\,
            in2 => \N__12343\,
            in3 => \N__28098\,
            lcout => alt_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29364\,
            ce => 'H',
            sr => \N__28739\
        );

    \Commands_frame_decoder.source_CH1data_1_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__12287\,
            in1 => \N__16892\,
            in2 => \N__27769\,
            in3 => \N__12324\,
            lcout => alt_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29364\,
            ce => 'H',
            sr => \N__28739\
        );

    \Commands_frame_decoder.source_CH1data8lto7_1_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27812\,
            in2 => \_gnd_net_\,
            in3 => \N__27622\,
            lcout => \Commands_frame_decoder.source_CH1data8lto7Z0Z_1\,
            ltout => \Commands_frame_decoder.source_CH1data8lto7Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data8lto7_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12259\,
            in1 => \N__28220\,
            in2 => \N__12310\,
            in3 => \N__27977\,
            lcout => \Commands_frame_decoder.source_CH1data8\,
            ltout => \Commands_frame_decoder.source_CH1data8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_0_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__16891\,
            in1 => \N__29845\,
            in2 => \N__12307\,
            in3 => \N__12303\,
            lcout => alt_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29364\,
            ce => 'H',
            sr => \N__28739\
        );

    \Commands_frame_decoder.source_CH1data_2_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__12288\,
            in1 => \N__16893\,
            in2 => \N__28362\,
            in3 => \N__12273\,
            lcout => alt_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29364\,
            ce => 'H',
            sr => \N__28739\
        );

    \Commands_frame_decoder.source_CH1data8lto3_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__28064\,
            in1 => \N__28308\,
            in2 => \_gnd_net_\,
            in3 => \N__27718\,
            lcout => \Commands_frame_decoder.source_CH1data8lt7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_4_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__17036\,
            in1 => \N__16999\,
            in2 => \N__17647\,
            in3 => \N__27825\,
            lcout => uart_pc_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12253\,
            lcout => drone_altitude_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12397\,
            lcout => drone_altitude_i_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_14_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15091\,
            lcout => drone_altitude_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29351\,
            ce => \N__13573\,
            sr => \N__28751\
        );

    \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14814\,
            lcout => \dron_frame_decoder_1.drone_altitude_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29351\,
            ce => \N__13573\,
            sr => \N__28751\
        );

    \ppm_encoder_1.un1_throttle_cry_0_c_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12999\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12699\,
            in2 => \N__27207\,
            in3 => \N__12391\,
            lcout => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_0\,
            carryout => \ppm_encoder_1.un1_throttle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12900\,
            in2 => \_gnd_net_\,
            in3 => \N__12388\,
            lcout => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_1\,
            carryout => \ppm_encoder_1.un1_throttle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12384\,
            in2 => \N__27208\,
            in3 => \N__12352\,
            lcout => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_2\,
            carryout => \ppm_encoder_1.un1_throttle_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12606\,
            in2 => \_gnd_net_\,
            in3 => \N__12349\,
            lcout => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_3\,
            carryout => \ppm_encoder_1.un1_throttle_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12567\,
            in2 => \_gnd_net_\,
            in3 => \N__12346\,
            lcout => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_4\,
            carryout => \ppm_encoder_1.un1_throttle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12477\,
            in2 => \N__27209\,
            in3 => \N__12451\,
            lcout => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_5\,
            carryout => \ppm_encoder_1.un1_throttle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12498\,
            in2 => \_gnd_net_\,
            in3 => \N__12448\,
            lcout => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_6\,
            carryout => \ppm_encoder_1.un1_throttle_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12543\,
            in2 => \_gnd_net_\,
            in3 => \N__12445\,
            lcout => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_20_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13791\,
            in2 => \_gnd_net_\,
            in3 => \N__12442\,
            lcout => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_8\,
            carryout => \ppm_encoder_1.un1_throttle_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12666\,
            in2 => \_gnd_net_\,
            in3 => \N__12439\,
            lcout => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_9\,
            carryout => \ppm_encoder_1.un1_throttle_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13755\,
            in2 => \_gnd_net_\,
            in3 => \N__12436\,
            lcout => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_10\,
            carryout => \ppm_encoder_1.un1_throttle_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13944\,
            in2 => \_gnd_net_\,
            in3 => \N__12433\,
            lcout => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_11\,
            carryout => \ppm_encoder_1.un1_throttle_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12639\,
            in2 => \N__27206\,
            in3 => \N__12430\,
            lcout => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_12\,
            carryout => \ppm_encoder_1.un1_throttle_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_14_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12427\,
            in2 => \_gnd_net_\,
            in3 => \N__12412\,
            lcout => \ppm_encoder_1.throttleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29340\,
            ce => \N__25066\,
            sr => \N__28764\
        );

    \ppm_encoder_1.throttle_1_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__24842\,
            in1 => \N__12703\,
            in2 => \N__14466\,
            in3 => \N__12679\,
            lcout => \ppm_encoder_1.throttleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29333\,
            ce => 'H',
            sr => \N__28770\
        );

    \ppm_encoder_1.throttle_10_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__12670\,
            in1 => \N__12646\,
            in2 => \N__22712\,
            in3 => \N__24840\,
            lcout => \ppm_encoder_1.throttleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29333\,
            ce => 'H',
            sr => \N__28770\
        );

    \ppm_encoder_1.throttle_13_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__24841\,
            in1 => \N__12640\,
            in2 => \N__20129\,
            in3 => \N__12616\,
            lcout => \ppm_encoder_1.throttleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29333\,
            ce => 'H',
            sr => \N__28770\
        );

    \ppm_encoder_1.throttle_4_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__24843\,
            in1 => \N__12610\,
            in2 => \N__13994\,
            in3 => \N__12589\,
            lcout => \ppm_encoder_1.throttleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29333\,
            ce => 'H',
            sr => \N__28770\
        );

    \ppm_encoder_1.throttle_5_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__12580\,
            in1 => \N__12571\,
            in2 => \N__24911\,
            in3 => \N__18605\,
            lcout => \ppm_encoder_1.throttleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29326\,
            ce => 'H',
            sr => \N__28774\
        );

    \ppm_encoder_1.throttle_8_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__12547\,
            in1 => \N__12520\,
            in2 => \N__13870\,
            in3 => \N__24853\,
            lcout => \ppm_encoder_1.throttleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29326\,
            ce => 'H',
            sr => \N__28774\
        );

    \ppm_encoder_1.throttle_7_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__12511\,
            in1 => \N__12502\,
            in2 => \N__24912\,
            in3 => \N__12744\,
            lcout => \ppm_encoder_1.throttleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29326\,
            ce => 'H',
            sr => \N__28774\
        );

    \ppm_encoder_1.elevator_7_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__24589\,
            in1 => \N__25966\,
            in2 => \N__24910\,
            in3 => \N__12724\,
            lcout => \ppm_encoder_1.elevatorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29326\,
            ce => 'H',
            sr => \N__28774\
        );

    \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__20408\,
            in1 => \N__15746\,
            in2 => \N__12748\,
            in3 => \N__15848\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14335\,
            in2 => \N__12757\,
            in3 => \N__12754\,
            lcout => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__12722\,
            in1 => \N__20150\,
            in2 => \N__16055\,
            in3 => \N__15970\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12743\,
            in1 => \N__22763\,
            in2 => \_gnd_net_\,
            in3 => \N__12723\,
            lcout => \ppm_encoder_1.N_298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_7_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__20151\,
            in1 => \N__22495\,
            in2 => \N__24908\,
            in3 => \N__24130\,
            lcout => \ppm_encoder_1.aileronZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29315\,
            ce => 'H',
            sr => \N__28776\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12850\,
            in1 => \N__12807\,
            in2 => \N__16319\,
            in3 => \N__23552\,
            lcout => \ppm_encoder_1.init_pulses_1_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__23556\,
            in1 => \N__12790\,
            in2 => \N__12709\,
            in3 => \N__15977\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIALN65_1_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001111"
        )
    port map (
            in0 => \N__14462\,
            in1 => \N__16264\,
            in2 => \N__12706\,
            in3 => \N__15847\,
            lcout => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18538\,
            in1 => \N__17809\,
            in2 => \N__23629\,
            in3 => \N__16311\,
            lcout => \ppm_encoder_1.init_pulses_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17941\,
            in2 => \_gnd_net_\,
            in3 => \N__18902\,
            lcout => \ppm_encoder_1.PPM_STATE_58_d\,
            ltout => \ppm_encoder_1.PPM_STATE_58_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18537\,
            in1 => \N__17808\,
            in2 => \N__12871\,
            in3 => \N__16312\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_1_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__18694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18904\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29307\,
            ce => 'H',
            sr => \N__28780\
        );

    \ppm_encoder_1.PPM_STATE_0_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__18903\,
            in1 => \N__18693\,
            in2 => \N__17951\,
            in3 => \N__18976\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29307\,
            ce => 'H',
            sr => \N__28780\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20666\,
            in2 => \_gnd_net_\,
            in3 => \N__23557\,
            lcout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12821\,
            in2 => \_gnd_net_\,
            in3 => \N__12865\,
            lcout => \ppm_encoder_1.N_226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011110110"
        )
    port map (
            in0 => \N__12808\,
            in1 => \N__23560\,
            in2 => \N__28980\,
            in3 => \N__20667\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__23559\,
            in1 => \N__20958\,
            in2 => \N__12849\,
            in3 => \N__28972\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__12866\,
            in1 => \N__12842\,
            in2 => \N__12828\,
            in3 => \N__12806\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__23558\,
            in1 => \_gnd_net_\,
            in2 => \N__12778\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.init_pulses_3_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__13995\,
            in1 => \N__12775\,
            in2 => \N__12760\,
            in3 => \N__15846\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__14002\,
            in1 => \N__18655\,
            in2 => \N__12943\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23651\,
            in1 => \N__15902\,
            in2 => \N__13135\,
            in3 => \N__16440\,
            lcout => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_2_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18227\,
            in1 => \N__12928\,
            in2 => \N__18026\,
            in3 => \N__14077\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29289\,
            ce => 'H',
            sr => \N__28787\
        );

    \ppm_encoder_1.throttle_RNIR7352_2_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__14378\,
            in1 => \N__15864\,
            in2 => \N__15909\,
            in3 => \N__16441\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI5V123_2_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12919\,
            in3 => \N__14097\,
            lcout => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIANUS_2_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__23650\,
            in1 => \N__20687\,
            in2 => \_gnd_net_\,
            in3 => \N__15901\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_2_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__12916\,
            in1 => \N__12907\,
            in2 => \N__24966\,
            in3 => \N__14379\,
            lcout => \ppm_encoder_1.throttleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29289\,
            ce => 'H',
            sr => \N__28787\
        );

    \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16442\,
            in1 => \N__13133\,
            in2 => \N__23798\,
            in3 => \N__21102\,
            lcout => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_0_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__13114\,
            in1 => \N__23761\,
            in2 => \N__12979\,
            in3 => \N__16448\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_0_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__13018\,
            in1 => \N__18010\,
            in2 => \N__13024\,
            in3 => \N__18243\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29283\,
            ce => 'H',
            sr => \N__28789\
        );

    \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12973\,
            in1 => \N__23760\,
            in2 => \_gnd_net_\,
            in3 => \N__20688\,
            lcout => \ppm_encoder_1.un1_init_pulses_0\,
            ltout => \ppm_encoder_1.un1_init_pulses_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_0_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18485\,
            in2 => \N__13021\,
            in3 => \N__15863\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12974\,
            in1 => \N__23762\,
            in2 => \N__13129\,
            in3 => \N__16447\,
            lcout => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIN3352_0_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \N__14127\,
            in1 => \N__18484\,
            in2 => \_gnd_net_\,
            in3 => \N__15862\,
            lcout => \ppm_encoder_1.throttle_RNIN3352Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_0_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__18486\,
            in1 => \N__24907\,
            in2 => \_gnd_net_\,
            in3 => \N__13006\,
            lcout => \ppm_encoder_1.throttleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29283\,
            ce => 'H',
            sr => \N__28789\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__20361\,
            in1 => \N__20555\,
            in2 => \_gnd_net_\,
            in3 => \N__12975\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__13128\,
            in1 => \N__21043\,
            in2 => \N__23809\,
            in3 => \N__16457\,
            lcout => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13124\,
            in2 => \_gnd_net_\,
            in3 => \N__23754\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__23755\,
            in1 => \_gnd_net_\,
            in2 => \N__13134\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23753\,
            in2 => \_gnd_net_\,
            in3 => \N__13123\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_17_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__18063\,
            in1 => \N__18244\,
            in2 => \N__14401\,
            in3 => \N__13075\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29277\,
            ce => 'H',
            sr => \N__28793\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22914\,
            in1 => \N__23756\,
            in2 => \_gnd_net_\,
            in3 => \N__20759\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_8_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18248\,
            in1 => \N__13054\,
            in2 => \N__18112\,
            in3 => \N__14266\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29270\,
            ce => 'H',
            sr => \N__28796\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__13040\,
            in1 => \_gnd_net_\,
            in2 => \N__23812\,
            in3 => \N__20792\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__20790\,
            in1 => \N__23772\,
            in2 => \_gnd_net_\,
            in3 => \N__13041\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__13042\,
            in1 => \N__20570\,
            in2 => \N__20382\,
            in3 => \N__19834\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_9_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18249\,
            in1 => \N__13030\,
            in2 => \N__18113\,
            in3 => \N__14221\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29270\,
            ce => 'H',
            sr => \N__28796\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__13220\,
            in1 => \_gnd_net_\,
            in2 => \N__23813\,
            in3 => \N__20793\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__20791\,
            in1 => \N__23773\,
            in2 => \_gnd_net_\,
            in3 => \N__13221\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__13222\,
            in1 => \N__20571\,
            in2 => \N__20383\,
            in3 => \N__19756\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20957\,
            in1 => \N__13210\,
            in2 => \_gnd_net_\,
            in3 => \N__15490\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset1data_6_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__16664\,
            in1 => \N__27632\,
            in2 => \N__13194\,
            in3 => \N__28977\,
            lcout => alt_kp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset1data_1_4_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__16663\,
            in1 => \N__27869\,
            in2 => \N__13173\,
            in3 => \N__28976\,
            lcout => alt_kp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_1_3_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15252\,
            in2 => \_gnd_net_\,
            in3 => \N__15189\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_a3_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_3_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15083\,
            in1 => \N__13253\,
            in2 => \N__13153\,
            in3 => \N__14809\,
            lcout => \dron_frame_decoder_1.state_ns_0_a3_0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_1_1_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14808\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15082\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_a3_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_1_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15190\,
            in1 => \N__15253\,
            in2 => \N__13150\,
            in3 => \N__13387\,
            lcout => \dron_frame_decoder_1.state_ns_0_a3_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_5_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__13683\,
            in1 => \N__13270\,
            in2 => \N__13483\,
            in3 => \N__13597\,
            lcout => \dron_frame_decoder_1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \N__28721\
        );

    \dron_frame_decoder_1.state_6_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__13684\,
            in1 => \N__13619\,
            in2 => \N__13484\,
            in3 => \N__13525\,
            lcout => \dron_frame_decoder_1.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \N__28721\
        );

    \dron_frame_decoder_1.state_3_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__13291\,
            in1 => \N__13682\,
            in2 => \N__13285\,
            in3 => \N__13347\,
            lcout => \dron_frame_decoder_1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \N__28721\
        );

    \dron_frame_decoder_1.state_7_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__13685\,
            in1 => \N__13620\,
            in2 => \N__13485\,
            in3 => \N__13651\,
            lcout => \dron_frame_decoder_1.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \N__28721\
        );

    \dron_frame_decoder_1.state_2_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__13269\,
            in1 => \N__13681\,
            in2 => \N__13284\,
            in3 => \N__13478\,
            lcout => \dron_frame_decoder_1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \N__28721\
        );

    \dron_frame_decoder_1.state_RNO_0_0_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__13360\,
            in1 => \N__13393\,
            in2 => \N__14872\,
            in3 => \N__13340\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.N_217_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_0_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__13386\,
            in1 => \N__13234\,
            in2 => \N__13261\,
            in3 => \N__13689\,
            lcout => \dron_frame_decoder_1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29370\,
            ce => 'H',
            sr => \N__28725\
        );

    \dron_frame_decoder_1.state_RNO_1_0_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13521\,
            in1 => \N__13385\,
            in2 => \N__13482\,
            in3 => \N__13257\,
            lcout => \dron_frame_decoder_1.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_5_0_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15049\,
            in2 => \_gnd_net_\,
            in3 => \N__15165\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_i_a2_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_2_0_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14793\,
            in1 => \N__13380\,
            in2 => \N__13396\,
            in3 => \N__15234\,
            lcout => \dron_frame_decoder_1.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_1_2_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27621\,
            in2 => \_gnd_net_\,
            in3 => \N__29831\,
            lcout => \Commands_frame_decoder.state_1_ns_0_a4_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_3_0_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__13526\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13381\,
            lcout => \dron_frame_decoder_1.state_ns_i_a2_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14971\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_i_a2_2_0_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15107\,
            in1 => \N__14831\,
            in2 => \N__13354\,
            in3 => \N__15283\,
            lcout => \dron_frame_decoder_1.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_ns_i_a2_3_1_0_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27957\,
            in2 => \_gnd_net_\,
            in3 => \N__27714\,
            lcout => \Commands_frame_decoder.state_1_ns_i_a2_3_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_esr_4_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27956\,
            lcout => alt_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29359\,
            ce => \N__16918\,
            sr => \N__28735\
        );

    \Commands_frame_decoder.source_CH1data_esr_5_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27826\,
            lcout => alt_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29359\,
            ce => \N__16918\,
            sr => \N__28735\
        );

    \Commands_frame_decoder.source_CH1data_esr_6_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28168\,
            lcout => alt_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29359\,
            ce => \N__16918\,
            sr => \N__28735\
        );

    \Commands_frame_decoder.source_CH1data_esr_7_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27623\,
            lcout => alt_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29359\,
            ce => \N__16918\,
            sr => \N__28735\
        );

    \dron_frame_decoder_1.state_RNI0TLI1_5_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__13534\,
            in1 => \N__13630\,
            in2 => \N__13603\,
            in3 => \N__28933\,
            lcout => \dron_frame_decoder_1.N_238_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_4_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__13424\,
            in1 => \N__13602\,
            in2 => \N__13650\,
            in3 => \N__13693\,
            lcout => \dron_frame_decoder_1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29352\,
            ce => 'H',
            sr => \N__28740\
        );

    \dron_frame_decoder_1.state_RNI6P6K_4_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13643\,
            in2 => \_gnd_net_\,
            in3 => \N__13423\,
            lcout => \dron_frame_decoder_1.un1_sink_data_valid_5_0_0\,
            ltout => \dron_frame_decoder_1.un1_sink_data_valid_5_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI3T3K1_7_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13624\,
            in1 => \N__13598\,
            in2 => \N__13579\,
            in3 => \N__13533\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI0AAT1_7_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13576\,
            in3 => \N__26687\,
            lcout => \dron_frame_decoder_1.N_230_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_data_valid_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__13828\,
            in1 => \N__13532\,
            in2 => \_gnd_net_\,
            in3 => \N__13441\,
            lcout => drone_frame_decoder_data_rdy_debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29346\,
            ce => 'H',
            sr => \N__28745\
        );

    \uart_pc.bit_Count_0_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__19370\,
            in1 => \N__19486\,
            in2 => \N__17283\,
            in3 => \N__19558\,
            lcout => \uart_pc.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29346\,
            ce => 'H',
            sr => \N__28745\
        );

    \uart_drone.data_rdy_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21760\,
            lcout => uart_drone_data_rdy_debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29346\,
            ce => 'H',
            sr => \N__28745\
        );

    \pid_alt.source_data_valid_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13829\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => pid_altitude_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29346\,
            ce => 'H',
            sr => \N__28745\
        );

    \Commands_frame_decoder.WDT_RNII19A1_4_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15435\,
            in1 => \N__15309\,
            in2 => \N__15421\,
            in3 => \N__15324\,
            lcout => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNI4U6E1_2_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17320\,
            in1 => \N__17370\,
            in2 => \_gnd_net_\,
            in3 => \N__17248\,
            lcout => \uart_pc.N_152\,
            ltout => \uart_pc.N_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIUPE73_3_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19482\,
            in2 => \N__13810\,
            in3 => \N__19555\,
            lcout => \uart_pc.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_2_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17321\,
            in1 => \N__17371\,
            in2 => \_gnd_net_\,
            in3 => \N__17249\,
            lcout => \uart_pc.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNO_0_2_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__17281\,
            in1 => \N__19556\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \uart_pc.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_2_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__13804\,
            in1 => \N__17386\,
            in2 => \N__13807\,
            in3 => \N__17339\,
            lcout => \uart_pc.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29334\,
            ce => 'H',
            sr => \N__28757\
        );

    \uart_pc.bit_Count_1_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__17282\,
            in1 => \N__19557\,
            in2 => \N__17348\,
            in3 => \N__13803\,
            lcout => \uart_pc.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29334\,
            ce => 'H',
            sr => \N__28757\
        );

    \ppm_encoder_1.throttle_9_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__13795\,
            in1 => \N__13771\,
            in2 => \N__24870\,
            in3 => \N__15456\,
            lcout => \ppm_encoder_1.throttleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29327\,
            ce => 'H',
            sr => \N__28765\
        );

    \ppm_encoder_1.throttle_11_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__13765\,
            in1 => \N__13954\,
            in2 => \N__24868\,
            in3 => \N__17918\,
            lcout => \ppm_encoder_1.throttleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29327\,
            ce => 'H',
            sr => \N__28765\
        );

    \ppm_encoder_1.throttle_12_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__13948\,
            in1 => \N__13915\,
            in2 => \N__24869\,
            in3 => \N__13900\,
            lcout => \ppm_encoder_1.throttleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29327\,
            ce => 'H',
            sr => \N__28765\
        );

    \ppm_encoder_1.throttle_RNII6JI2_12_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__20040\,
            in1 => \N__13898\,
            in2 => \N__15881\,
            in3 => \N__15769\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIFQRT5_12_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__14200\,
            in1 => \_gnd_net_\,
            in2 => \N__13909\,
            in3 => \N__13906\,
            lcout => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI25DH2_12_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__22875\,
            in1 => \N__13880\,
            in2 => \N__16065\,
            in3 => \N__15991\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13899\,
            in1 => \N__22876\,
            in2 => \_gnd_net_\,
            in3 => \N__22799\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20938\,
            in1 => \_gnd_net_\,
            in2 => \N__13885\,
            in3 => \N__13881\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_12_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__13882\,
            in1 => \N__23926\,
            in2 => \N__24909\,
            in3 => \N__22420\,
            lcout => \ppm_encoder_1.aileronZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29316\,
            ce => 'H',
            sr => \N__28771\
        );

    \ppm_encoder_1.throttle_RNIS5KK2_8_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__13865\,
            in1 => \N__15765\,
            in2 => \N__19830\,
            in3 => \N__15851\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIONI96_8_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14296\,
            in2 => \N__13849\,
            in3 => \N__14017\,
            lcout => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNICKVN2_8_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__19797\,
            in1 => \N__15479\,
            in2 => \N__15989\,
            in3 => \N__16042\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIU7KK2_9_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__15852\,
            in1 => \N__15457\,
            in2 => \N__15772\,
            in3 => \N__19749\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNITSI96_9_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14251\,
            in2 => \N__14011\,
            in3 => \N__14008\,
            lcout => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__15850\,
            in1 => \N__20184\,
            in2 => \N__15771\,
            in3 => \N__19900\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIEMVN2_9_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__19614\,
            in1 => \N__19875\,
            in2 => \N__15990\,
            in3 => \N__16043\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__13962\,
            in1 => \N__14427\,
            in2 => \N__15988\,
            in3 => \N__16041\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_4_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24208\,
            lcout => \ppm_encoder_1.aileronZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29299\,
            ce => \N__25050\,
            sr => \N__28777\
        );

    \ppm_encoder_1.elevator_esr_4_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24508\,
            lcout => \ppm_encoder_1.elevatorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29299\,
            ce => \N__25050\,
            sr => \N__28777\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13996\,
            in1 => \N__13963\,
            in2 => \_gnd_net_\,
            in3 => \N__18563\,
            lcout => \ppm_encoder_1.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__17715\,
            in1 => \N__18612\,
            in2 => \N__15757\,
            in3 => \N__15849\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__17752\,
            in1 => \_gnd_net_\,
            in2 => \N__14149\,
            in3 => \N__14146\,
            lcout => \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__18582\,
            in1 => \N__18507\,
            in2 => \N__16056\,
            in3 => \N__15969\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIVO123_0_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14140\,
            in2 => \N__14131\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_25_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_1_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16260\,
            in2 => \N__14113\,
            in3 => \N__14104\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_2_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14101\,
            in2 => \N__14086\,
            in3 => \N__14071\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_3_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14068\,
            in2 => \N__14053\,
            in3 => \N__14032\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_4_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18654\,
            in2 => \N__14029\,
            in3 => \N__14020\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_5_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17745\,
            in2 => \N__14365\,
            in3 => \N__14356\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_6_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18357\,
            in2 => \N__14353\,
            in3 => \N__14338\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_7_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14334\,
            in2 => \N__14311\,
            in3 => \N__14299\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_8_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14292\,
            in2 => \N__14278\,
            in3 => \N__14254\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_8\,
            ltout => OPEN,
            carryin => \bfn_3_26_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_9_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14247\,
            in2 => \N__14233\,
            in3 => \N__14209\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_10_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15687\,
            in2 => \N__15661\,
            in3 => \N__14206\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_11_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16104\,
            in2 => \N__16078\,
            in3 => \N__14203\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_12_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14199\,
            in2 => \N__14179\,
            in3 => \N__14167\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_13_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16344\,
            in2 => \N__14164\,
            in3 => \N__14413\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_14_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18294\,
            in2 => \N__15616\,
            in3 => \N__14410\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_15_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16504\,
            in2 => \N__16381\,
            in3 => \N__14407\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_16_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14524\,
            in2 => \_gnd_net_\,
            in3 => \N__14404\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_16\,
            ltout => OPEN,
            carryin => \bfn_3_27_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_17_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14386\,
            in2 => \_gnd_net_\,
            in3 => \N__14392\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_18_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16405\,
            in2 => \_gnd_net_\,
            in3 => \N__14389\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22913\,
            in1 => \N__23795\,
            in2 => \_gnd_net_\,
            in3 => \N__20798\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22856\,
            in2 => \N__16333\,
            in3 => \N__20885\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010111110"
        )
    port map (
            in0 => \N__28960\,
            in1 => \N__23796\,
            in2 => \N__20931\,
            in3 => \N__20799\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__20921\,
            in1 => \N__22855\,
            in2 => \_gnd_net_\,
            in3 => \N__14380\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22955\,
            in1 => \N__23794\,
            in2 => \_gnd_net_\,
            in3 => \N__20797\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_16_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18231\,
            in1 => \N__14518\,
            in2 => \N__18094\,
            in3 => \N__14506\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29271\,
            ce => 'H',
            sr => \N__28790\
        );

    \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__21147\,
            in1 => \N__14488\,
            in2 => \N__14476\,
            in3 => \N__22591\,
            lcout => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_8_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23106\,
            in1 => \N__14500\,
            in2 => \_gnd_net_\,
            in3 => \N__14494\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29267\,
            ce => \N__23061\,
            sr => \N__28794\
        );

    \ppm_encoder_1.pulses2count_esr_9_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23107\,
            in1 => \N__15643\,
            in2 => \_gnd_net_\,
            in3 => \N__14482\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29267\,
            ce => \N__23061\,
            sr => \N__28794\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__20932\,
            in1 => \N__22857\,
            in2 => \_gnd_net_\,
            in3 => \N__14467\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20933\,
            in1 => \N__14440\,
            in2 => \_gnd_net_\,
            in3 => \N__14431\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14559\,
            in2 => \_gnd_net_\,
            in3 => \N__14580\,
            lcout => OPEN,
            ltout => \reset_module_System.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__16782\,
            in1 => \N__16702\,
            in2 => \N__14416\,
            in3 => \N__16597\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__16701\,
            in1 => \N__14536\,
            in2 => \N__16783\,
            in3 => \N__16596\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIR9N6_1_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14576\,
            lcout => \reset_module_System.reset6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14637\,
            in1 => \N__14652\,
            in2 => \N__14623\,
            in3 => \N__14670\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIA72I1_16_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__14710\,
            in1 => \N__14731\,
            in2 => \N__14596\,
            in3 => \N__14593\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIMJ304_12_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14758\,
            in1 => \N__14557\,
            in2 => \N__14587\,
            in3 => \N__14881\,
            lcout => \reset_module_System.reset6_19\,
            ltout => \reset_module_System.reset6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__14558\,
            in1 => \N__16777\,
            in2 => \N__14584\,
            in3 => \N__16700\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14581\,
            in2 => \N__14560\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16794\,
            in2 => \_gnd_net_\,
            in3 => \N__14530\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16824\,
            in2 => \_gnd_net_\,
            in3 => \N__14527\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__29374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14686\,
            in2 => \_gnd_net_\,
            in3 => \N__14674\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__29374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14671\,
            in2 => \_gnd_net_\,
            in3 => \N__14659\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__29374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16836\,
            in2 => \_gnd_net_\,
            in3 => \N__14656\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__29374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14653\,
            in2 => \_gnd_net_\,
            in3 => \N__14641\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__29374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14638\,
            in2 => \_gnd_net_\,
            in3 => \N__14626\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__29374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14619\,
            in2 => \_gnd_net_\,
            in3 => \N__14605\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16740\,
            in2 => \_gnd_net_\,
            in3 => \N__14602\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16713\,
            in2 => \_gnd_net_\,
            in3 => \N__14599\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14754\,
            in2 => \_gnd_net_\,
            in3 => \N__14743\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14893\,
            in2 => \_gnd_net_\,
            in3 => \N__14740\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16752\,
            in2 => \_gnd_net_\,
            in3 => \N__14737\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14917\,
            in2 => \_gnd_net_\,
            in3 => \N__14734\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14730\,
            in2 => \_gnd_net_\,
            in3 => \N__14716\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16725\,
            in2 => \_gnd_net_\,
            in3 => \N__14713\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__29365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14709\,
            in2 => \_gnd_net_\,
            in3 => \N__14695\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__29365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14926\,
            in2 => \_gnd_net_\,
            in3 => \N__14692\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__29365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16809\,
            in2 => \_gnd_net_\,
            in3 => \N__14689\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__29365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14904\,
            in2 => \_gnd_net_\,
            in3 => \N__14929\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14925\,
            in1 => \N__14916\,
            in2 => \N__14905\,
            in3 => \N__14892\,
            lcout => \reset_module_System.reset6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_4_0_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15233\,
            in1 => \N__15050\,
            in2 => \N__14799\,
            in3 => \N__15169\,
            lcout => \dron_frame_decoder_1.state_ns_i_a2_0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIES9Q1_2_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__21756\,
            in1 => \N__17135\,
            in2 => \_gnd_net_\,
            in3 => \N__26647\,
            lcout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\,
            ltout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIRC5U2_2_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__17136\,
            in1 => \_gnd_net_\,
            in2 => \N__14860\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.state_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_5_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__28203\,
            in1 => \N__17037\,
            in2 => \N__17593\,
            in3 => \N__16987\,
            lcout => uart_pc_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_0_2_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__28312\,
            in1 => \N__27857\,
            in2 => \N__14857\,
            in3 => \N__24361\,
            lcout => \Commands_frame_decoder.state_1_ns_0_a4_0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_esr_0_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21505\,
            lcout => uart_drone_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_drone.data_esr_1_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21487\,
            lcout => uart_drone_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_drone.data_esr_2_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21841\,
            lcout => uart_drone_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_drone.data_esr_3_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_drone_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_drone.data_esr_4_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21655\,
            lcout => uart_drone_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_drone.data_esr_5_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17088\,
            lcout => uart_drone_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_drone.data_esr_6_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17073\,
            lcout => uart_drone_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_drone.data_esr_7_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17058\,
            lcout => uart_drone_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29353\,
            ce => \N__14950\,
            sr => \N__14944\
        );

    \uart_pc.data_3_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__16993\,
            in1 => \N__28063\,
            in2 => \N__17698\,
            in3 => \N__17024\,
            lcout => uart_pc_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26646\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19327\,
            lcout => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\,
            ltout => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__17188\,
            in1 => \N__16992\,
            in2 => \N__14932\,
            in3 => \N__27713\,
            lcout => uart_pc_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_4_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19328\,
            in1 => \N__16991\,
            in2 => \N__27976\,
            in3 => \N__17671\,
            lcout => uart_pc_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_0_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15358\,
            in2 => \N__17415\,
            in3 => \N__17416\,
            lcout => \Commands_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_0\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_1_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15352\,
            in2 => \_gnd_net_\,
            in3 => \N__15346\,
            lcout => \Commands_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_0\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_1\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_2_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15343\,
            in2 => \_gnd_net_\,
            in3 => \N__15337\,
            lcout => \Commands_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_1\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_2\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_3_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15334\,
            in2 => \_gnd_net_\,
            in3 => \N__15328\,
            lcout => \Commands_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_2\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_3\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_4_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15325\,
            in2 => \_gnd_net_\,
            in3 => \N__15313\,
            lcout => \Commands_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_3\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_4\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_5_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15310\,
            in2 => \_gnd_net_\,
            in3 => \N__15298\,
            lcout => \Commands_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_4\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_5\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_6_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15582\,
            in2 => \_gnd_net_\,
            in3 => \N__15295\,
            lcout => \Commands_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_5\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_6\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_7_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15552\,
            in2 => \_gnd_net_\,
            in3 => \N__15292\,
            lcout => \Commands_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_6\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_7\,
            clk => \N__29341\,
            ce => 'H',
            sr => \N__17112\
        );

    \Commands_frame_decoder.WDT_8_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15436\,
            in2 => \_gnd_net_\,
            in3 => \N__15424\,
            lcout => \Commands_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_19_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_8\,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_9_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15420\,
            in2 => \_gnd_net_\,
            in3 => \N__15406\,
            lcout => \Commands_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_8\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_9\,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_10_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15370\,
            in2 => \_gnd_net_\,
            in3 => \N__15403\,
            lcout => \Commands_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_9\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_10\,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_11_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15598\,
            in2 => \_gnd_net_\,
            in3 => \N__15400\,
            lcout => \Commands_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_10\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_11\,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_12_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15568\,
            in2 => \_gnd_net_\,
            in3 => \N__15397\,
            lcout => \Commands_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_11\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_12\,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_13_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15384\,
            in2 => \_gnd_net_\,
            in3 => \N__15394\,
            lcout => \Commands_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_12\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_13\,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_14_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22337\,
            in2 => \_gnd_net_\,
            in3 => \N__15391\,
            lcout => \Commands_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_13\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_14\,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_15_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17438\,
            in2 => \_gnd_net_\,
            in3 => \N__15388\,
            lcout => \Commands_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29335\,
            ce => 'H',
            sr => \N__17116\
        );

    \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__15566\,
            in1 => \N__15596\,
            in2 => \N__15385\,
            in3 => \N__15369\,
            lcout => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_1_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__17387\,
            in1 => \N__17322\,
            in2 => \_gnd_net_\,
            in3 => \N__17277\,
            lcout => \uart_pc.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_3_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__17278\,
            in1 => \_gnd_net_\,
            in2 => \N__17340\,
            in3 => \N__17388\,
            lcout => \uart_pc.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNID7P31_6_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15597\,
            in1 => \N__15583\,
            in2 => \_gnd_net_\,
            in3 => \N__15567\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.WDT8lto13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__15553\,
            in1 => \N__15538\,
            in2 => \N__15532\,
            in3 => \N__15529\,
            lcout => \Commands_frame_decoder.WDT8lt14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_4_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17389\,
            in1 => \N__17326\,
            in2 => \_gnd_net_\,
            in3 => \N__17279\,
            lcout => \uart_pc.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_5_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__17280\,
            in1 => \_gnd_net_\,
            in2 => \N__17341\,
            in3 => \N__17390\,
            lcout => \uart_pc.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110010011110100"
        )
    port map (
            in0 => \N__22510\,
            in1 => \N__15631\,
            in2 => \N__15507\,
            in3 => \N__17956\,
            lcout => ppm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29317\,
            ce => 'H',
            sr => \N__28758\
        );

    \ppm_encoder_1.aileron_8_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__22477\,
            in1 => \N__24091\,
            in2 => \N__24798\,
            in3 => \N__15483\,
            lcout => \ppm_encoder_1.aileronZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29317\,
            ce => 'H',
            sr => \N__28758\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22828\,
            in1 => \N__15455\,
            in2 => \_gnd_net_\,
            in3 => \N__19615\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20934\,
            in2 => \N__15646\,
            in3 => \N__19876\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_0_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18969\,
            in2 => \_gnd_net_\,
            in3 => \N__18935\,
            lcout => \ppm_encoder_1.N_139_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_5_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24265\,
            lcout => \ppm_encoder_1.aileronZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29300\,
            ce => \N__25042\,
            sr => \N__28772\
        );

    \ppm_encoder_1.elevator_esr_5_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24250\,
            lcout => \ppm_encoder_1.elevatorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29300\,
            ce => \N__25042\,
            sr => \N__28772\
        );

    \ppm_encoder_1.rudder_esr_5_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24232\,
            lcout => \ppm_encoder_1.rudderZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29300\,
            ce => \N__25042\,
            sr => \N__28772\
        );

    \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__18295\,
            in1 => \_gnd_net_\,
            in2 => \N__15625\,
            in3 => \N__15604\,
            lcout => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIU0DH2_10_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__22683\,
            in1 => \N__16061\,
            in2 => \N__19963\,
            in3 => \N__15993\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__15994\,
            in1 => \N__25099\,
            in2 => \N__16066\,
            in3 => \N__22387\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIG4JI2_11_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__17919\,
            in1 => \N__19710\,
            in2 => \N__15883\,
            in3 => \N__15770\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIALRT5_11_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__16105\,
            in1 => \_gnd_net_\,
            in2 => \N__16081\,
            in3 => \N__15922\,
            lcout => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI03DH2_11_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__24675\,
            in1 => \N__16060\,
            in2 => \N__17898\,
            in3 => \N__15992\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16148\,
            in1 => \N__20559\,
            in2 => \_gnd_net_\,
            in3 => \N__19711\,
            lcout => \ppm_encoder_1.N_318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000101"
        )
    port map (
            in0 => \N__20004\,
            in1 => \N__20551\,
            in2 => \N__20351\,
            in3 => \N__16243\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__20553\,
            in1 => \N__20322\,
            in2 => \N__15916\,
            in3 => \N__20005\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__20323\,
            in1 => \N__20552\,
            in2 => \N__16193\,
            in3 => \N__19639\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIE2JI2_10_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__22713\,
            in1 => \N__19638\,
            in2 => \N__15882\,
            in3 => \N__15761\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI5GRT5_10_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__15688\,
            in1 => \_gnd_net_\,
            in2 => \N__15670\,
            in3 => \N__15667\,
            lcout => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__20327\,
            in1 => \_gnd_net_\,
            in2 => \N__20010\,
            in3 => \N__15652\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_ctle_14_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24797\,
            in2 => \_gnd_net_\,
            in3 => \N__28925\,
            lcout => \ppm_encoder_1.pid_altitude_dv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17823\,
            in1 => \N__16326\,
            in2 => \N__18570\,
            in3 => \N__18937\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16288\,
            in3 => \N__18968\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1\,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_1_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__16285\,
            in1 => \N__18049\,
            in2 => \N__16279\,
            in3 => \N__16276\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29279\,
            ce => 'H',
            sr => \N__28781\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__16239\,
            in1 => \_gnd_net_\,
            in2 => \N__23799\,
            in3 => \N__20714\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__20713\,
            in1 => \N__23733\,
            in2 => \_gnd_net_\,
            in3 => \N__16238\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_10_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18198\,
            in1 => \N__16213\,
            in2 => \N__18079\,
            in3 => \N__16201\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29279\,
            ce => 'H',
            sr => \N__28781\
        );

    \ppm_encoder_1.init_pulses_11_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__18200\,
            in1 => \N__18045\,
            in2 => \N__16171\,
            in3 => \N__16156\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29279\,
            ce => 'H',
            sr => \N__28781\
        );

    \ppm_encoder_1.init_pulses_12_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18199\,
            in1 => \N__16123\,
            in2 => \N__18080\,
            in3 => \N__16111\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29279\,
            ce => 'H',
            sr => \N__28781\
        );

    \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23788\,
            in1 => \N__23885\,
            in2 => \N__20809\,
            in3 => \N__16458\,
            lcout => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_15_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__18205\,
            in1 => \N__18090\,
            in2 => \N__16492\,
            in3 => \N__16477\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29272\,
            ce => 'H',
            sr => \N__28783\
        );

    \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__23784\,
            in1 => \N__23886\,
            in2 => \_gnd_net_\,
            in3 => \N__20784\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_2_18_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__16459\,
            in1 => \N__17552\,
            in2 => \N__20806\,
            in3 => \N__23787\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_18_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18202\,
            in1 => \N__16399\,
            in2 => \N__18111\,
            in3 => \N__16387\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29272\,
            ce => 'H',
            sr => \N__28783\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23786\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_13_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18201\,
            in1 => \N__16369\,
            in2 => \N__18110\,
            in3 => \N__16357\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29272\,
            ce => 'H',
            sr => \N__28783\
        );

    \ppm_encoder_1.init_pulses_RNISFRP_13_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20785\,
            in1 => \N__21032\,
            in2 => \_gnd_net_\,
            in3 => \N__23785\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__16555\,
            in1 => \N__22633\,
            in2 => \N__16549\,
            in3 => \N__22612\,
            lcout => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_4_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__23096\,
            in1 => \_gnd_net_\,
            in2 => \N__16579\,
            in3 => \N__16567\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29268\,
            ce => \N__23052\,
            sr => \N__28788\
        );

    \ppm_encoder_1.pulses2count_esr_5_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18394\,
            in1 => \N__18496\,
            in2 => \_gnd_net_\,
            in3 => \N__23097\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29268\,
            ce => \N__23052\,
            sr => \N__28788\
        );

    \ppm_encoder_1.pulses2count_esr_10_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23093\,
            in1 => \N__19933\,
            in2 => \_gnd_net_\,
            in3 => \N__16540\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29268\,
            ce => \N__23052\,
            sr => \N__28788\
        );

    \ppm_encoder_1.pulses2count_esr_11_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23094\,
            in1 => \N__17872\,
            in2 => \_gnd_net_\,
            in3 => \N__16531\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29268\,
            ce => \N__23052\,
            sr => \N__28788\
        );

    \ppm_encoder_1.pulses2count_esr_12_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16522\,
            in1 => \N__23095\,
            in2 => \_gnd_net_\,
            in3 => \N__19975\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29268\,
            ce => \N__23052\,
            sr => \N__28788\
        );

    \ppm_encoder_1.counter24_0_I_1_c_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18778\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_29_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18445\,
            in2 => \N__27272\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_0\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16510\,
            in2 => \N__27266\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_1\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23236\,
            in2 => \N__27269\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_2\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16609\,
            in2 => \N__27267\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_3\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18724\,
            in2 => \N__27270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_4\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18712\,
            in2 => \N__27268\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_5\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22978\,
            in2 => \N__27271\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_6\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18847\,
            in2 => \N__27274\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_30_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18853\,
            in2 => \N__27275\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_8\,
            carryout => \ppm_encoder_1.counter24_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16600\,
            lcout => \ppm_encoder_1.counter24_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__16781\,
            in1 => \N__16699\,
            in2 => \_gnd_net_\,
            in3 => \N__16595\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNI08RE_4_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16852\,
            in2 => \_gnd_net_\,
            in3 => \N__29618\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__16837\,
            in1 => \N__16825\,
            in2 => \N__16813\,
            in3 => \N__16795\,
            lcout => \reset_module_System.reset6_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNILR1B2_2_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__19092\,
            in1 => \N__19339\,
            in2 => \_gnd_net_\,
            in3 => \N__26608\,
            lcout => \uart_pc.timer_Count_RNILR1B2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNISRMR1_10_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16756\,
            in1 => \N__16741\,
            in2 => \N__16729\,
            in3 => \N__16714\,
            lcout => \reset_module_System.reset6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_0_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__16971\,
            in1 => \N__17041\,
            in2 => \N__29826\,
            in3 => \N__17212\,
            lcout => uart_pc_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNIVM1O_6_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__25616\,
            in1 => \N__29600\,
            in2 => \_gnd_net_\,
            in3 => \N__28926\,
            lcout => \Commands_frame_decoder.state_1_RNIVM1OZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNI19RE_5_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16944\,
            in2 => \_gnd_net_\,
            in3 => \N__29587\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_6_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25612\,
            in2 => \N__16633\,
            in3 => \N__29459\,
            lcout => \Commands_frame_decoder.state_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29361\,
            ce => 'H',
            sr => \N__28717\
        );

    \Commands_frame_decoder.source_offset1data_4_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__16623\,
            in1 => \N__29588\,
            in2 => \N__25617\,
            in3 => \N__27972\,
            lcout => alt_kp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29361\,
            ce => 'H',
            sr => \N__28717\
        );

    \Commands_frame_decoder.state_1_5_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__16945\,
            in1 => \N__24652\,
            in2 => \_gnd_net_\,
            in3 => \N__29458\,
            lcout => \Commands_frame_decoder.state_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29361\,
            ce => 'H',
            sr => \N__28717\
        );

    \uart_pc.data_rdy_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19338\,
            lcout => uart_pc_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29361\,
            ce => 'H',
            sr => \N__28717\
        );

    \Commands_frame_decoder.state_1_ns_i_a2_3_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29591\,
            in1 => \N__28076\,
            in2 => \N__28175\,
            in3 => \N__16936\,
            lcout => \Commands_frame_decoder.N_323\,
            ltout => \Commands_frame_decoder.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_2_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__16906\,
            in1 => \N__16927\,
            in2 => \N__16921\,
            in3 => \N__29455\,
            lcout => \Commands_frame_decoder.state_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29354\,
            ce => 'H',
            sr => \N__28722\
        );

    \Commands_frame_decoder.state_1_RNIRI1O_2_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16878\,
            in2 => \_gnd_net_\,
            in3 => \N__28938\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNIU5RE_2_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16905\,
            in2 => \_gnd_net_\,
            in3 => \N__29589\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0\,
            ltout => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_3_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__29456\,
            in1 => \_gnd_net_\,
            in2 => \N__16867\,
            in3 => \N__16864\,
            lcout => \Commands_frame_decoder.state_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29354\,
            ce => 'H',
            sr => \N__28722\
        );

    \Commands_frame_decoder.state_1_RNIV6RE_3_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16863\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_4_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16851\,
            in2 => \N__16855\,
            in3 => \N__29457\,
            lcout => \Commands_frame_decoder.state_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29354\,
            ce => 'H',
            sr => \N__28722\
        );

    \uart_drone.data_Aux_5_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19165\,
            in1 => \N__21746\,
            in2 => \N__17089\,
            in3 => \N__21775\,
            lcout => \uart_drone.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29348\,
            ce => 'H',
            sr => \N__21586\
        );

    \uart_drone.data_Aux_6_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19228\,
            in1 => \N__21747\,
            in2 => \N__17074\,
            in3 => \N__21776\,
            lcout => \uart_drone.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29348\,
            ce => 'H',
            sr => \N__21586\
        );

    \uart_drone.data_Aux_7_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__21777\,
            in1 => \N__21748\,
            in2 => \N__17059\,
            in3 => \N__25525\,
            lcout => \uart_drone.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29348\,
            ce => 'H',
            sr => \N__21586\
        );

    \uart_pc.data_2_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__17025\,
            in1 => \N__16994\,
            in2 => \N__17158\,
            in3 => \N__28307\,
            lcout => uart_pc_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_0_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__21552\,
            in1 => \N__17516\,
            in2 => \N__19278\,
            in3 => \N__26625\,
            lcout => \uart_drone.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__29614\,
            in1 => \N__22338\,
            in2 => \N__17443\,
            in3 => \N__22305\,
            lcout => \Commands_frame_decoder.N_316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_1_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17515\,
            in2 => \_gnd_net_\,
            in3 => \N__17535\,
            lcout => OPEN,
            ltout => \uart_drone.timer_Count_RNO_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_1_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__26624\,
            in1 => \N__19274\,
            in2 => \N__17044\,
            in3 => \N__21553\,
            lcout => \uart_drone.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI9ADK1_4_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__19191\,
            in1 => \N__25582\,
            in2 => \N__17497\,
            in3 => \N__21887\,
            lcout => \uart_drone.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_6_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__17026\,
            in1 => \N__16995\,
            in2 => \N__17626\,
            in3 => \N__27577\,
            lcout => uart_pc_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_4_0_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17439\,
            in2 => \_gnd_net_\,
            in3 => \N__29613\,
            lcout => \Commands_frame_decoder.state_1_RNO_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_2_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__26622\,
            in1 => \N__17470\,
            in2 => \N__19291\,
            in3 => \N__21557\,
            lcout => \uart_drone.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_6_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__17273\,
            in1 => \N__17398\,
            in2 => \_gnd_net_\,
            in3 => \N__17350\,
            lcout => \uart_pc.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIDGR31_2_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__21917\,
            in1 => \N__17483\,
            in2 => \N__21999\,
            in3 => \N__21888\,
            lcout => \uart_drone.state_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.un1_state49_i_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29640\,
            in2 => \_gnd_net_\,
            in3 => \N__28929\,
            lcout => \Commands_frame_decoder.un1_state49_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI9E9J_2_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17484\,
            lcout => \uart_drone.N_126_li\,
            ltout => \uart_drone.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIAT1D1_4_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__21889\,
            in1 => \N__21985\,
            in2 => \N__17095\,
            in3 => \N__26621\,
            lcout => \uart_drone.N_143\,
            ltout => \uart_drone.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_3_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__19289\,
            in1 => \N__26626\,
            in2 => \N__17092\,
            in3 => \N__17461\,
            lcout => \uart_drone.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_4_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__17449\,
            in1 => \N__19290\,
            in2 => \N__21564\,
            in3 => \N__26623\,
            lcout => \uart_drone.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI5A9J_1_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__17520\,
            in1 => \N__17536\,
            in2 => \N__17521\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_5_19_0_\,
            carryout => \uart_drone.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_2_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17485\,
            in2 => \_gnd_net_\,
            in3 => \N__17464\,
            lcout => \uart_drone.timer_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_1\,
            carryout => \uart_drone.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_3_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21922\,
            in2 => \_gnd_net_\,
            in3 => \N__17455\,
            lcout => \uart_drone.timer_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_2\,
            carryout => \uart_drone.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_4_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21991\,
            in2 => \_gnd_net_\,
            in3 => \N__17452\,
            lcout => \uart_drone.timer_Count_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_RNIF92K5_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__22330\,
            in1 => \N__17432\,
            in2 => \N__27388\,
            in3 => \N__22298\,
            lcout => \Commands_frame_decoder.state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_0_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17397\,
            in1 => \N__17349\,
            in2 => \_gnd_net_\,
            in3 => \N__17284\,
            lcout => \uart_pc.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_0_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__17221\,
            in1 => \N__19133\,
            in2 => \N__17211\,
            in3 => \N__19428\,
            lcout => \uart_pc.data_AuxZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29318\,
            ce => 'H',
            sr => \N__19581\
        );

    \uart_pc.data_Aux_1_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__19429\,
            in1 => \N__17181\,
            in2 => \N__19152\,
            in3 => \N__17194\,
            lcout => \uart_pc.data_AuxZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29318\,
            ce => 'H',
            sr => \N__19581\
        );

    \uart_pc.data_Aux_2_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__17170\,
            in1 => \N__19137\,
            in2 => \N__17154\,
            in3 => \N__19430\,
            lcout => \uart_pc.data_AuxZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29318\,
            ce => 'H',
            sr => \N__19581\
        );

    \uart_pc.data_Aux_3_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__19431\,
            in1 => \N__17688\,
            in2 => \N__19153\,
            in3 => \N__17704\,
            lcout => \uart_pc.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29318\,
            ce => 'H',
            sr => \N__19581\
        );

    \uart_pc.data_Aux_4_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__17677\,
            in1 => \N__19141\,
            in2 => \N__17670\,
            in3 => \N__19432\,
            lcout => \uart_pc.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29318\,
            ce => 'H',
            sr => \N__19581\
        );

    \uart_pc.data_Aux_5_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__19433\,
            in1 => \N__17637\,
            in2 => \N__19154\,
            in3 => \N__17653\,
            lcout => \uart_pc.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29318\,
            ce => 'H',
            sr => \N__19581\
        );

    \uart_pc.data_Aux_7_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__19434\,
            in1 => \N__17616\,
            in2 => \N__19155\,
            in3 => \N__19378\,
            lcout => \uart_pc.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29318\,
            ce => 'H',
            sr => \N__19581\
        );

    \uart_pc.data_Aux_6_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__19156\,
            in1 => \N__17605\,
            in2 => \N__17586\,
            in3 => \N__19435\,
            lcout => \uart_pc.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29308\,
            ce => 'H',
            sr => \N__19585\
        );

    \ppm_encoder_1.pulses2count_18_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__23808\,
            in1 => \N__23850\,
            in2 => \N__17569\,
            in3 => \N__18867\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29290\,
            ce => 'H',
            sr => \N__28766\
        );

    \ppm_encoder_1.rudder_7_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__19393\,
            in1 => \N__24867\,
            in2 => \N__20412\,
            in3 => \N__25468\,
            lcout => \ppm_encoder_1.rudderZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29290\,
            ce => 'H',
            sr => \N__28766\
        );

    \ppm_encoder_1.rudder_6_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__24865\,
            in1 => \N__25132\,
            in2 => \_gnd_net_\,
            in3 => \N__21065\,
            lcout => \ppm_encoder_1.rudderZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29290\,
            ce => 'H',
            sr => \N__28766\
        );

    \ppm_encoder_1.aileron_11_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__23965\,
            in1 => \N__24866\,
            in2 => \N__17899\,
            in3 => \N__22435\,
            lcout => \ppm_encoder_1.aileronZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29290\,
            ce => 'H',
            sr => \N__28766\
        );

    \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21235\,
            in1 => \N__20224\,
            in2 => \N__21202\,
            in3 => \N__17952\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__17923\,
            in1 => \_gnd_net_\,
            in2 => \N__22846\,
            in3 => \N__24676\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__17894\,
            in1 => \_gnd_net_\,
            in2 => \N__17875\,
            in3 => \N__20948\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22815\,
            in1 => \N__17819\,
            in2 => \_gnd_net_\,
            in3 => \N__17859\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010101"
        )
    port map (
            in0 => \N__17860\,
            in1 => \_gnd_net_\,
            in2 => \N__17824\,
            in3 => \N__22816\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_5_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18209\,
            in1 => \N__17773\,
            in2 => \N__18114\,
            in3 => \N__17761\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29280\,
            ce => 'H',
            sr => \N__28775\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__18405\,
            in1 => \_gnd_net_\,
            in2 => \N__23823\,
            in3 => \N__20775\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20774\,
            in1 => \N__18404\,
            in2 => \_gnd_net_\,
            in3 => \N__23800\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__17719\,
            in1 => \N__20321\,
            in2 => \N__18409\,
            in3 => \N__20569\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_6_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18210\,
            in1 => \N__18385\,
            in2 => \N__18115\,
            in3 => \N__18370\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29280\,
            ce => 'H',
            sr => \N__28775\
        );

    \ppm_encoder_1.init_pulses_RNIERUS_6_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__21089\,
            in1 => \_gnd_net_\,
            in2 => \N__23824\,
            in3 => \N__20776\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_7_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__18340\,
            in1 => \N__18107\,
            in2 => \N__18328\,
            in3 => \N__18211\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29280\,
            ce => 'H',
            sr => \N__28775\
        );

    \ppm_encoder_1.init_pulses_14_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18203\,
            in1 => \N__18316\,
            in2 => \N__18108\,
            in3 => \N__18304\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29273\,
            ce => 'H',
            sr => \N__28778\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_14_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19913\,
            in1 => \N__23749\,
            in2 => \_gnd_net_\,
            in3 => \N__20780\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20778\,
            in1 => \_gnd_net_\,
            in2 => \N__23807\,
            in3 => \N__19914\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22968\,
            in1 => \N__23748\,
            in2 => \_gnd_net_\,
            in3 => \N__20779\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_4_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18204\,
            in1 => \N__18130\,
            in2 => \N__18109\,
            in3 => \N__17968\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29273\,
            ce => 'H',
            sr => \N__28778\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_4_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__18666\,
            in1 => \N__23744\,
            in2 => \_gnd_net_\,
            in3 => \N__20777\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__22849\,
            in1 => \N__20922\,
            in2 => \_gnd_net_\,
            in3 => \N__18637\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18616\,
            in1 => \N__18589\,
            in2 => \_gnd_net_\,
            in3 => \N__18571\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20923\,
            in1 => \_gnd_net_\,
            in2 => \N__18517\,
            in3 => \N__18514\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__20924\,
            in1 => \N__22848\,
            in2 => \_gnd_net_\,
            in3 => \N__18490\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__20360\,
            in1 => \N__20537\,
            in2 => \N__20017\,
            in3 => \N__18469\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21231\,
            in1 => \N__18928\,
            in2 => \N__21198\,
            in3 => \N__20220\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__18415\,
            in1 => \N__21191\,
            in2 => \N__18814\,
            in3 => \N__21230\,
            lcout => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_2_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23125\,
            in1 => \N__18439\,
            in2 => \_gnd_net_\,
            in3 => \N__18427\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29265\,
            ce => \N__23060\,
            sr => \N__28784\
        );

    \ppm_encoder_1.pulses2count_esr_3_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18829\,
            in1 => \N__23126\,
            in2 => \_gnd_net_\,
            in3 => \N__18820\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29265\,
            ce => \N__23060\,
            sr => \N__28784\
        );

    \ppm_encoder_1.pulses2count_esr_0_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__23123\,
            in1 => \_gnd_net_\,
            in2 => \N__18805\,
            in3 => \N__18796\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29265\,
            ce => \N__23060\,
            sr => \N__28784\
        );

    \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__20219\,
            in1 => \N__18784\,
            in2 => \N__18748\,
            in3 => \N__20244\,
            lcout => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_1_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23124\,
            in1 => \N__18772\,
            in2 => \_gnd_net_\,
            in3 => \N__18760\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29265\,
            ce => \N__23060\,
            sr => \N__28784\
        );

    \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__18739\,
            in1 => \N__21297\,
            in2 => \N__18733\,
            in3 => \N__21123\,
            lcout => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23314\,
            in1 => \N__18718\,
            in2 => \N__23170\,
            in3 => \N__22570\,
            lcout => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIK1KG_0_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21124\,
            in1 => \N__21148\,
            in2 => \N__21301\,
            in3 => \N__20248\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\,
            ltout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23386\,
            in1 => \N__18706\,
            in2 => \N__18697\,
            in3 => \N__22546\,
            lcout => \ppm_encoder_1.N_237\,
            ltout => \ppm_encoder_1.N_237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__26642\,
            in1 => \N__18958\,
            in2 => \N__18940\,
            in3 => \N__18936\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18868\,
            in2 => \_gnd_net_\,
            in3 => \N__23427\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22939\,
            in1 => \N__23470\,
            in2 => \N__22897\,
            in3 => \N__23449\,
            lcout => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_2__0__0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23353\,
            lcout => \uart_pc_sync.aux_2__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.Q_0__0_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18835\,
            lcout => uart_commands_input_debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_3__0__0_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18841\,
            lcout => \uart_pc_sync.aux_3__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH2data_esr_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29838\,
            lcout => \frame_decoder_CH2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29367\,
            ce => \N__21339\,
            sr => \N__28711\
        );

    \Commands_frame_decoder.source_CH2data_esr_5_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27871\,
            lcout => \frame_decoder_CH2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29355\,
            ce => \N__21338\,
            sr => \N__28715\
        );

    \Commands_frame_decoder.source_CH2data_esr_6_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28221\,
            lcout => \frame_decoder_CH2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29355\,
            ce => \N__21338\,
            sr => \N__28715\
        );

    \Commands_frame_decoder.source_CH2data_esr_4_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27989\,
            lcout => \frame_decoder_CH2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29355\,
            ce => \N__21338\,
            sr => \N__28715\
        );

    \Commands_frame_decoder.source_CH2data_esr_1_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27736\,
            lcout => \frame_decoder_CH2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29355\,
            ce => \N__21338\,
            sr => \N__28715\
        );

    \Commands_frame_decoder.source_CH2data_esr_3_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28105\,
            lcout => \frame_decoder_CH2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29355\,
            ce => \N__21338\,
            sr => \N__28715\
        );

    \Commands_frame_decoder.source_CH2data_esr_2_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28354\,
            lcout => \frame_decoder_CH2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29355\,
            ce => \N__21338\,
            sr => \N__28715\
        );

    \uart_drone.bit_Count_RNIJOJC1_2_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__26348\,
            in1 => \N__26271\,
            in2 => \_gnd_net_\,
            in3 => \N__26109\,
            lcout => \uart_drone.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNIUL1O_5_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__19018\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28935\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNISJ1O_3_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19009\,
            in2 => \_gnd_net_\,
            in3 => \N__28936\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_2_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__21619\,
            in1 => \N__21754\,
            in2 => \N__18994\,
            in3 => \N__28948\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_2_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__18993\,
            in1 => \N__22020\,
            in2 => \N__18997\,
            in3 => \N__21944\,
            lcout => \uart_drone.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_1_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__18992\,
            in1 => \N__19177\,
            in2 => \N__28981\,
            in3 => \N__21755\,
            lcout => \uart_drone.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__28949\,
            in1 => \N__19038\,
            in2 => \N__19213\,
            in3 => \N__19104\,
            lcout => \uart_pc.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_6_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__26353\,
            in1 => \N__26273\,
            in2 => \_gnd_net_\,
            in3 => \N__26111\,
            lcout => \uart_drone.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__19209\,
            in1 => \N__19094\,
            in2 => \_gnd_net_\,
            in3 => \N__28946\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_0_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__22242\,
            in1 => \N__19528\,
            in2 => \N__19216\,
            in3 => \N__19513\,
            lcout => \uart_pc.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_0_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__21750\,
            in1 => \N__19176\,
            in2 => \_gnd_net_\,
            in3 => \N__28945\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_0_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__19198\,
            in1 => \N__22019\,
            in2 => \N__19180\,
            in3 => \N__21881\,
            lcout => \uart_drone.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_5_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__26341\,
            in1 => \N__26272\,
            in2 => \_gnd_net_\,
            in3 => \N__26110\,
            lcout => \uart_drone.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_2_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__19250\,
            in1 => \N__19093\,
            in2 => \N__19039\,
            in3 => \N__28947\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_2_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__22243\,
            in1 => \N__19037\,
            in2 => \N__19021\,
            in3 => \N__22060\,
            lcout => \uart_pc.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_3_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__19249\,
            in1 => \N__19348\,
            in2 => \N__19300\,
            in3 => \N__26694\,
            lcout => \uart_pc.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNI5UFA2_3_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22053\,
            in1 => \_gnd_net_\,
            in2 => \N__22240\,
            in3 => \N__19377\,
            lcout => \uart_pc.N_144_1\,
            ltout => \uart_pc.N_144_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_4_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__22118\,
            in1 => \N__19475\,
            in2 => \N__19342\,
            in3 => \N__26695\,
            lcout => \uart_pc.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIPD2K1_2_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__22052\,
            in1 => \N__22271\,
            in2 => \N__22239\,
            in3 => \N__19508\,
            lcout => \uart_pc.state_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_3_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__22230\,
            in1 => \N__22054\,
            in2 => \N__19251\,
            in3 => \N__19474\,
            lcout => \uart_pc.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI40411_2_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__25567\,
            in1 => \N__22014\,
            in2 => \N__21630\,
            in3 => \N__21946\,
            lcout => \uart_drone.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIGRIF1_2_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110000"
        )
    port map (
            in0 => \N__22231\,
            in1 => \N__22055\,
            in2 => \N__19252\,
            in3 => \N__19473\,
            lcout => \uart_pc.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_3_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__25566\,
            in1 => \N__22015\,
            in2 => \N__21629\,
            in3 => \N__21945\,
            lcout => \uart_drone.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIMQ8T1_4_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__19524\,
            in1 => \N__19510\,
            in2 => \N__22238\,
            in3 => \N__26683\,
            lcout => \uart_pc.N_143\,
            ltout => \uart_pc.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_2_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__26685\,
            in1 => \N__22083\,
            in2 => \N__19588\,
            in3 => \N__22255\,
            lcout => \uart_pc.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIEAGS_4_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__19472\,
            in1 => \N__19512\,
            in2 => \_gnd_net_\,
            in3 => \N__28928\,
            lcout => \uart_pc.state_RNIEAGSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_4_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__26686\,
            in1 => \N__22180\,
            in2 => \N__22092\,
            in3 => \N__22117\,
            lcout => \uart_pc.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIITIF1_4_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110011"
        )
    port map (
            in0 => \N__22050\,
            in1 => \N__19465\,
            in2 => \N__22237\,
            in3 => \N__19509\,
            lcout => \uart_pc.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_0_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__26684\,
            in1 => \N__22084\,
            in2 => \N__22174\,
            in3 => \N__22116\,
            lcout => \uart_pc.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__22051\,
            in1 => \N__22272\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.N_126_li\,
            ltout => \uart_pc.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIBLRB2_4_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011101110"
        )
    port map (
            in0 => \N__19511\,
            in1 => \N__19471\,
            in2 => \N__19438\,
            in3 => \N__22282\,
            lcout => \uart_pc.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25131\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \ppm_encoder_1.un1_rudder_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25461\,
            in2 => \_gnd_net_\,
            in3 => \N__19381\,
            lcout => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_6\,
            carryout => \ppm_encoder_1.un1_rudder_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25437\,
            in2 => \_gnd_net_\,
            in3 => \N__19669\,
            lcout => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_7\,
            carryout => \ppm_encoder_1.un1_rudder_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25413\,
            in2 => \_gnd_net_\,
            in3 => \N__19666\,
            lcout => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_8\,
            carryout => \ppm_encoder_1.un1_rudder_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25389\,
            in2 => \_gnd_net_\,
            in3 => \N__19663\,
            lcout => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_9\,
            carryout => \ppm_encoder_1.un1_rudder_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25365\,
            in2 => \_gnd_net_\,
            in3 => \N__19660\,
            lcout => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_10\,
            carryout => \ppm_encoder_1.un1_rudder_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25341\,
            in2 => \_gnd_net_\,
            in3 => \N__19657\,
            lcout => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_11\,
            carryout => \ppm_encoder_1.un1_rudder_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25314\,
            in2 => \N__27276\,
            in3 => \N__19654\,
            lcout => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_12\,
            carryout => \ppm_encoder_1.un1_rudder_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_14_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25291\,
            in2 => \_gnd_net_\,
            in3 => \N__19651\,
            lcout => \ppm_encoder_1.rudderZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29301\,
            ce => \N__25076\,
            sr => \N__28746\
        );

    \ppm_encoder_1.rudder_10_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__19648\,
            in1 => \N__25393\,
            in2 => \N__19637\,
            in3 => \N__24950\,
            lcout => \ppm_encoder_1.rudderZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29291\,
            ce => 'H',
            sr => \N__28752\
        );

    \ppm_encoder_1.elevator_9_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__24553\,
            in1 => \N__25915\,
            in2 => \N__19613\,
            in3 => \N__24949\,
            lcout => \ppm_encoder_1.elevatorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29291\,
            ce => 'H',
            sr => \N__28752\
        );

    \ppm_encoder_1.aileron_10_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__24010\,
            in1 => \N__22450\,
            in2 => \N__24964\,
            in3 => \N__19952\,
            lcout => \ppm_encoder_1.aileronZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29291\,
            ce => 'H',
            sr => \N__28752\
        );

    \ppm_encoder_1.aileron_9_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__22462\,
            in1 => \N__24052\,
            in2 => \N__19874\,
            in3 => \N__24947\,
            lcout => \ppm_encoder_1.aileronZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29291\,
            ce => 'H',
            sr => \N__28752\
        );

    \ppm_encoder_1.rudder_8_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__19843\,
            in1 => \N__25441\,
            in2 => \N__24965\,
            in3 => \N__19817\,
            lcout => \ppm_encoder_1.rudderZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29291\,
            ce => 'H',
            sr => \N__28752\
        );

    \ppm_encoder_1.elevator_8_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__24568\,
            in1 => \N__25939\,
            in2 => \N__19796\,
            in3 => \N__24948\,
            lcout => \ppm_encoder_1.elevatorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29291\,
            ce => 'H',
            sr => \N__28752\
        );

    \ppm_encoder_1.rudder_9_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__19765\,
            in1 => \N__25417\,
            in2 => \N__19748\,
            in3 => \N__24940\,
            lcout => \ppm_encoder_1.rudderZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29284\,
            ce => 'H',
            sr => \N__28759\
        );

    \ppm_encoder_1.rudder_11_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__25369\,
            in1 => \N__19720\,
            in2 => \N__19709\,
            in3 => \N__24938\,
            lcout => \ppm_encoder_1.rudderZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29284\,
            ce => 'H',
            sr => \N__28759\
        );

    \ppm_encoder_1.rudder_12_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__25345\,
            in1 => \N__19687\,
            in2 => \N__24963\,
            in3 => \N__20039\,
            lcout => \ppm_encoder_1.rudderZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29284\,
            ce => 'H',
            sr => \N__28759\
        );

    \ppm_encoder_1.rudder_13_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__25321\,
            in1 => \N__19678\,
            in2 => \N__21015\,
            in3 => \N__24939\,
            lcout => \ppm_encoder_1.rudderZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29284\,
            ce => 'H',
            sr => \N__28759\
        );

    \ppm_encoder_1.aileron_13_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__22402\,
            in1 => \N__24307\,
            in2 => \N__24962\,
            in3 => \N__20087\,
            lcout => \ppm_encoder_1.aileronZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29284\,
            ce => 'H',
            sr => \N__28759\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25098\,
            in1 => \N__22850\,
            in2 => \_gnd_net_\,
            in3 => \N__20191\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20960\,
            in2 => \N__20170\,
            in3 => \N__22386\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20961\,
            in1 => \N__20167\,
            in2 => \_gnd_net_\,
            in3 => \N__20155\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22851\,
            in1 => \N__20137\,
            in2 => \_gnd_net_\,
            in3 => \N__25005\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20962\,
            in1 => \_gnd_net_\,
            in2 => \N__20098\,
            in3 => \N__20091\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20544\,
            in1 => \N__20068\,
            in2 => \_gnd_net_\,
            in3 => \N__20041\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20009\,
            in2 => \N__19978\,
            in3 => \N__20345\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20947\,
            in1 => \N__22657\,
            in2 => \_gnd_net_\,
            in3 => \N__19962\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__20514\,
            in1 => \N__19918\,
            in2 => \N__20379\,
            in3 => \N__19896\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__20517\,
            in1 => \N__21103\,
            in2 => \N__21076\,
            in3 => \N__20365\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101001111"
        )
    port map (
            in0 => \N__20515\,
            in1 => \N__21042\,
            in2 => \N__20380\,
            in3 => \N__21014\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23821\,
            lcout => \ppm_encoder_1.N_590_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__22858\,
            in1 => \N__20920\,
            in2 => \N__20545\,
            in3 => \N__20808\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__20516\,
            in1 => \N__26707\,
            in2 => \N__20575\,
            in3 => \N__23822\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__20513\,
            in1 => \N__20440\,
            in2 => \N__20416\,
            in3 => \N__20369\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_0_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20243\,
            in2 => \N__20265\,
            in3 => \N__20266\,
            lcout => \ppm_encoder_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_28_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_0\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_1_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20218\,
            in2 => \_gnd_net_\,
            in3 => \N__20194\,
            lcout => \ppm_encoder_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_0\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_1\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_2_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21229\,
            in2 => \_gnd_net_\,
            in3 => \N__21205\,
            lcout => \ppm_encoder_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_1\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_2\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_3_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21190\,
            in2 => \_gnd_net_\,
            in3 => \N__21166\,
            lcout => \ppm_encoder_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_2\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_3\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_4_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22611\,
            in2 => \_gnd_net_\,
            in3 => \N__21163\,
            lcout => \ppm_encoder_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_3\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_4\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_5_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22632\,
            in2 => \_gnd_net_\,
            in3 => \N__21160\,
            lcout => \ppm_encoder_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_4\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_5\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_6_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23254\,
            in2 => \_gnd_net_\,
            in3 => \N__21157\,
            lcout => \ppm_encoder_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_5\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_6\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_7_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23286\,
            in2 => \_gnd_net_\,
            in3 => \N__21154\,
            lcout => \ppm_encoder_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_6\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_7\,
            clk => \N__29262\,
            ce => 'H',
            sr => \N__21256\
        );

    \ppm_encoder_1.counter_8_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22590\,
            in2 => \_gnd_net_\,
            in3 => \N__21151\,
            lcout => \ppm_encoder_1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_29_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_8\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_9_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21146\,
            in2 => \_gnd_net_\,
            in3 => \N__21127\,
            lcout => \ppm_encoder_1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_8\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_9\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_10_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21122\,
            in2 => \_gnd_net_\,
            in3 => \N__21106\,
            lcout => \ppm_encoder_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_9\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_10\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_11_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21296\,
            in2 => \_gnd_net_\,
            in3 => \N__21280\,
            lcout => \ppm_encoder_1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_10\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_11\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_12_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22569\,
            in2 => \_gnd_net_\,
            in3 => \N__21277\,
            lcout => \ppm_encoder_1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_11\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_12\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_13_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23313\,
            in2 => \_gnd_net_\,
            in3 => \N__21274\,
            lcout => \ppm_encoder_1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_12\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_13\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_14_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22996\,
            in2 => \_gnd_net_\,
            in3 => \N__21271\,
            lcout => \ppm_encoder_1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_13\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_14\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_15_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23404\,
            in2 => \_gnd_net_\,
            in3 => \N__21268\,
            lcout => \ppm_encoder_1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_14\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_15\,
            clk => \N__29261\,
            ce => 'H',
            sr => \N__21255\
        );

    \ppm_encoder_1.counter_16_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23448\,
            in2 => \_gnd_net_\,
            in3 => \N__21265\,
            lcout => \ppm_encoder_1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_30_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_16\,
            clk => \N__29259\,
            ce => 'H',
            sr => \N__21254\
        );

    \ppm_encoder_1.counter_17_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23469\,
            in2 => \_gnd_net_\,
            in3 => \N__21262\,
            lcout => \ppm_encoder_1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_16\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_17\,
            clk => \N__29259\,
            ce => 'H',
            sr => \N__21254\
        );

    \ppm_encoder_1.counter_18_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23426\,
            in2 => \_gnd_net_\,
            in3 => \N__21259\,
            lcout => \ppm_encoder_1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29259\,
            ce => 'H',
            sr => \N__21254\
        );

    \uart_drone_sync.aux_0__0__0_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21241\,
            lcout => \uart_drone_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_2__0__0_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21358\,
            lcout => \uart_drone_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_1__0__0_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21364\,
            lcout => \uart_drone_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_3__0__0_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21352\,
            lcout => \uart_drone_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.Q_0__0_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21346\,
            lcout => uart_drone_input_debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH2data_ess_7_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27647\,
            lcout => \frame_decoder_CH2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29368\,
            ce => \N__21340\,
            sr => \N__28712\
        );

    \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23340\,
            in2 => \_gnd_net_\,
            in3 => \N__21309\,
            lcout => \scaler_2.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.N_521_i_l_ofx_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__21310\,
            in1 => \_gnd_net_\,
            in2 => \N__23344\,
            in3 => \_gnd_net_\,
            lcout => \scaler_2.N_521_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset2data_esr_6_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28213\,
            lcout => \frame_decoder_OFF2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29356\,
            ce => \N__24625\,
            sr => \N__28716\
        );

    \Commands_frame_decoder.source_offset2data_esr_3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28114\,
            lcout => \frame_decoder_OFF2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29356\,
            ce => \N__24625\,
            sr => \N__28716\
        );

    \Commands_frame_decoder.source_offset2data_esr_5_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27883\,
            lcout => \frame_decoder_OFF2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29356\,
            ce => \N__24625\,
            sr => \N__28716\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25198\,
            in2 => \N__25241\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21466\,
            in2 => \N__23332\,
            in3 => \N__21457\,
            lcout => \scaler_2.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_0\,
            carryout => \scaler_2.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21454\,
            in2 => \N__24181\,
            in3 => \N__21448\,
            lcout => \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_1\,
            carryout => \scaler_2.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21445\,
            in2 => \N__21439\,
            in3 => \N__21430\,
            lcout => \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_2\,
            carryout => \scaler_2.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21427\,
            in2 => \N__23323\,
            in3 => \N__21418\,
            lcout => \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_3\,
            carryout => \scaler_2.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21415\,
            in2 => \N__21409\,
            in3 => \N__21400\,
            lcout => \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_4\,
            carryout => \scaler_2.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21397\,
            in2 => \N__21391\,
            in3 => \N__21379\,
            lcout => \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_5\,
            carryout => \scaler_2.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21376\,
            in2 => \_gnd_net_\,
            in3 => \N__21367\,
            lcout => \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_6\,
            carryout => \scaler_2.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21520\,
            in2 => \N__27265\,
            in3 => \N__21511\,
            lcout => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21508\,
            lcout => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_3_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__26349\,
            in1 => \N__26278\,
            in2 => \_gnd_net_\,
            in3 => \N__26113\,
            lcout => \uart_drone.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_ns_0_a4_0_0_1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27617\,
            in2 => \_gnd_net_\,
            in3 => \N__29827\,
            lcout => \Commands_frame_decoder.state_1_ns_0_a4_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIU8TV1_3_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25522\,
            in1 => \N__22021\,
            in2 => \_gnd_net_\,
            in3 => \N__21943\,
            lcout => \uart_drone.N_144_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_2_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__26112\,
            in1 => \N__26340\,
            in2 => \_gnd_net_\,
            in3 => \N__26274\,
            lcout => \uart_drone.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__25819\,
            in1 => \N__25861\,
            in2 => \_gnd_net_\,
            in3 => \N__26810\,
            lcout => \scaler_4.un2_source_data_0_cry_1_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_0_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__24214\,
            in1 => \N__21738\,
            in2 => \N__21504\,
            in3 => \N__21792\,
            lcout => \uart_drone.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29329\,
            ce => 'H',
            sr => \N__21576\
        );

    \uart_drone.data_Aux_1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__21793\,
            in1 => \N__26206\,
            in2 => \N__21483\,
            in3 => \N__21740\,
            lcout => \uart_drone.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29329\,
            ce => 'H',
            sr => \N__21576\
        );

    \uart_drone.data_Aux_2_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__21847\,
            in1 => \N__21739\,
            in2 => \N__21840\,
            in3 => \N__21794\,
            lcout => \uart_drone.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29329\,
            ce => 'H',
            sr => \N__21576\
        );

    \uart_drone.data_Aux_3_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__21795\,
            in1 => \N__21823\,
            in2 => \N__21813\,
            in3 => \N__21741\,
            lcout => \uart_drone.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29329\,
            ce => 'H',
            sr => \N__21576\
        );

    \uart_drone.data_Aux_4_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__21796\,
            in1 => \N__21637\,
            in2 => \N__21654\,
            in3 => \N__21742\,
            lcout => \uart_drone.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29329\,
            ce => 'H',
            sr => \N__21576\
        );

    \uart_drone.data_Aux_RNO_0_4_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__26243\,
            in1 => \N__26313\,
            in2 => \_gnd_net_\,
            in3 => \N__26095\,
            lcout => \uart_drone.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_0_1_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28310\,
            in1 => \N__27853\,
            in2 => \N__24394\,
            in3 => \N__24448\,
            lcout => \Commands_frame_decoder.state_1_ns_0_a4_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_3_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__21531\,
            in1 => \N__21631\,
            in2 => \N__21598\,
            in3 => \N__26692\,
            lcout => \uart_drone.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIOU0N_4_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__25571\,
            in1 => \N__21880\,
            in2 => \_gnd_net_\,
            in3 => \N__28931\,
            lcout => \uart_drone.state_RNIOU0NZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_1_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__22120\,
            in1 => \N__22091\,
            in2 => \N__22138\,
            in3 => \N__26693\,
            lcout => \uart_pc.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_4_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__26691\,
            in1 => \N__21565\,
            in2 => \N__25583\,
            in3 => \N__21532\,
            lcout => \uart_drone.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_1_0_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__22360\,
            in1 => \N__24393\,
            in2 => \N__22348\,
            in3 => \N__22309\,
            lcout => \Commands_frame_decoder.state_1_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIRP8S_1_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__22165\,
            in1 => \N__22149\,
            in2 => \N__22173\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \uart_pc.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_2_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22273\,
            in2 => \_gnd_net_\,
            in3 => \N__22249\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_1\,
            carryout => \uart_pc.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_3_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22056\,
            in2 => \_gnd_net_\,
            in3 => \N__22246\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_2\,
            carryout => \uart_pc.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_4_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22241\,
            in2 => \_gnd_net_\,
            in3 => \N__22183\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_1_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22169\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22150\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_3_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__22126\,
            in1 => \N__22119\,
            in2 => \N__22093\,
            in3 => \N__26696\,
            lcout => \uart_pc.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI62411_4_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__21998\,
            in1 => \N__21931\,
            in2 => \N__25578\,
            in3 => \N__21876\,
            lcout => \uart_drone.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_c_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24162\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24129\,
            in2 => \_gnd_net_\,
            in3 => \N__22480\,
            lcout => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_6\,
            carryout => \ppm_encoder_1.un1_aileron_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24084\,
            in2 => \_gnd_net_\,
            in3 => \N__22465\,
            lcout => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_7\,
            carryout => \ppm_encoder_1.un1_aileron_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24048\,
            in2 => \_gnd_net_\,
            in3 => \N__22453\,
            lcout => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_8\,
            carryout => \ppm_encoder_1.un1_aileron_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24003\,
            in2 => \_gnd_net_\,
            in3 => \N__22438\,
            lcout => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_9\,
            carryout => \ppm_encoder_1.un1_aileron_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23958\,
            in2 => \_gnd_net_\,
            in3 => \N__22423\,
            lcout => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_10\,
            carryout => \ppm_encoder_1.un1_aileron_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23919\,
            in2 => \_gnd_net_\,
            in3 => \N__22405\,
            lcout => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_11\,
            carryout => \ppm_encoder_1.un1_aileron_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24306\,
            in2 => \N__27296\,
            in3 => \N__22393\,
            lcout => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_12\,
            carryout => \ppm_encoder_1.un1_aileron_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_14_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24277\,
            in2 => \_gnd_net_\,
            in3 => \N__22390\,
            lcout => \ppm_encoder_1.aileronZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29292\,
            ce => \N__25078\,
            sr => \N__28753\
        );

    \ppm_encoder_1.elevator_10_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__25888\,
            in1 => \N__24535\,
            in2 => \N__24960\,
            in3 => \N__22676\,
            lcout => \ppm_encoder_1.elevatorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29285\,
            ce => 'H',
            sr => \N__28760\
        );

    \ppm_encoder_1.elevator_12_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__24520\,
            in1 => \N__26452\,
            in2 => \N__24959\,
            in3 => \N__22874\,
            lcout => \ppm_encoder_1.elevatorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29281\,
            ce => 'H',
            sr => \N__28767\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22847\,
            in1 => \N__22717\,
            in2 => \_gnd_net_\,
            in3 => \N__22684\,
            lcout => \ppm_encoder_1.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_7_LC_8_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23127\,
            in1 => \N__22651\,
            in2 => \_gnd_net_\,
            in3 => \N__22639\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29263\,
            ce => \N__23062\,
            sr => \N__28785\
        );

    \ppm_encoder_1.counter_RNIUS1G_4_LC_8_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23253\,
            in1 => \N__22631\,
            in2 => \N__23287\,
            in3 => \N__22610\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIAEV01_8_LC_8_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22589\,
            in1 => \N__22568\,
            in2 => \N__22549\,
            in3 => \N__23293\,
            lcout => \ppm_encoder_1.N_144_17\,
            ltout => \ppm_encoder_1.N_144_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_1_LC_8_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22534\,
            in1 => \N__22525\,
            in2 => \N__22513\,
            in3 => \N__23385\,
            lcout => \ppm_encoder_1.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_8_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28930\,
            in2 => \_gnd_net_\,
            in3 => \N__23797\,
            lcout => \ppm_encoder_1.N_590_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIDBJ8_13_LC_8_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22995\,
            in2 => \_gnd_net_\,
            in3 => \N__23312\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_8_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23200\,
            in1 => \N__23282\,
            in2 => \N__23266\,
            in3 => \N__23252\,
            lcout => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_6_LC_8_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23227\,
            in1 => \N__23137\,
            in2 => \_gnd_net_\,
            in3 => \N__23209\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29260\,
            ce => \N__23056\,
            sr => \N__28791\
        );

    \ppm_encoder_1.pulses2count_esr_13_LC_8_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23194\,
            in1 => \N__23135\,
            in2 => \_gnd_net_\,
            in3 => \N__23179\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29260\,
            ce => \N__23056\,
            sr => \N__28791\
        );

    \ppm_encoder_1.pulses2count_esr_14_LC_8_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23158\,
            in1 => \N__23146\,
            in2 => \_gnd_net_\,
            in3 => \N__23136\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29260\,
            ce => \N__23056\,
            sr => \N__28791\
        );

    \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23002\,
            in1 => \N__23402\,
            in2 => \N__23485\,
            in3 => \N__22994\,
            lcout => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_16_LC_8_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__22969\,
            in1 => \N__22938\,
            in2 => \N__23872\,
            in3 => \N__23827\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29258\,
            ce => 'H',
            sr => \N__28795\
        );

    \ppm_encoder_1.pulses2count_17_LC_8_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__23825\,
            in1 => \N__22924\,
            in2 => \N__22896\,
            in3 => \N__23870\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29258\,
            ce => 'H',
            sr => \N__28795\
        );

    \ppm_encoder_1.pulses2count_15_LC_8_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__23893\,
            in1 => \N__23484\,
            in2 => \N__23871\,
            in3 => \N__23826\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29258\,
            ce => 'H',
            sr => \N__28795\
        );

    \ppm_encoder_1.counter_RNI637H_18_LC_8_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23468\,
            in1 => \N__23447\,
            in2 => \N__23428\,
            in3 => \N__23403\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_0__0__0_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23365\,
            lcout => \uart_pc_sync.aux_0__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_1__0__0_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23359\,
            lcout => \uart_pc_sync.aux_1__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset2data_ess_7_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29362\,
            ce => \N__24617\,
            sr => \N__28713\
        );

    \Commands_frame_decoder.source_offset2data_esr_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29860\,
            lcout => \frame_decoder_OFF2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29349\,
            ce => \N__24624\,
            sr => \N__28718\
        );

    \Commands_frame_decoder.source_offset2data_esr_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27774\,
            lcout => \frame_decoder_OFF2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29349\,
            ce => \N__24624\,
            sr => \N__28718\
        );

    \Commands_frame_decoder.source_offset2data_esr_4_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27993\,
            lcout => \frame_decoder_OFF2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29349\,
            ce => \N__24624\,
            sr => \N__28718\
        );

    \Commands_frame_decoder.source_offset2data_esr_2_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28361\,
            lcout => \frame_decoder_OFF2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29349\,
            ce => \N__24624\,
            sr => \N__28718\
        );

    \scaler_2.un2_source_data_0_cry_1_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25261\,
            in2 => \N__25165\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_6_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24138\,
            in2 => \N__25271\,
            in3 => \N__24145\,
            lcout => scaler_2_data_6,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_1\,
            carryout => \scaler_2.un2_source_data_0_cry_2\,
            clk => \N__29344\,
            ce => \N__26374\,
            sr => \N__28723\
        );

    \scaler_2.source_data_1_esr_7_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24099\,
            in2 => \N__24142\,
            in3 => \N__24106\,
            lcout => scaler_2_data_7,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_2\,
            carryout => \scaler_2.un2_source_data_0_cry_3\,
            clk => \N__29344\,
            ce => \N__26374\,
            sr => \N__28723\
        );

    \scaler_2.source_data_1_esr_8_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24060\,
            in2 => \N__24103\,
            in3 => \N__24067\,
            lcout => scaler_2_data_8,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_3\,
            carryout => \scaler_2.un2_source_data_0_cry_4\,
            clk => \N__29344\,
            ce => \N__26374\,
            sr => \N__28723\
        );

    \scaler_2.source_data_1_esr_9_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24018\,
            in2 => \N__24064\,
            in3 => \N__24025\,
            lcout => scaler_2_data_9,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_4\,
            carryout => \scaler_2.un2_source_data_0_cry_5\,
            clk => \N__29344\,
            ce => \N__26374\,
            sr => \N__28723\
        );

    \scaler_2.source_data_1_esr_10_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23973\,
            in2 => \N__24022\,
            in3 => \N__23980\,
            lcout => scaler_2_data_10,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_5\,
            carryout => \scaler_2.un2_source_data_0_cry_6\,
            clk => \N__29344\,
            ce => \N__26374\,
            sr => \N__28723\
        );

    \scaler_2.source_data_1_esr_11_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23934\,
            in2 => \N__23977\,
            in3 => \N__23941\,
            lcout => scaler_2_data_11,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_6\,
            carryout => \scaler_2.un2_source_data_0_cry_7\,
            clk => \N__29344\,
            ce => \N__26374\,
            sr => \N__28723\
        );

    \scaler_2.source_data_1_esr_12_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24327\,
            in2 => \N__23938\,
            in3 => \N__23896\,
            lcout => scaler_2_data_12,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_7\,
            carryout => \scaler_2.un2_source_data_0_cry_8\,
            clk => \N__29344\,
            ce => \N__26374\,
            sr => \N__28723\
        );

    \scaler_2.source_data_1_esr_13_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24328\,
            in2 => \N__24316\,
            in3 => \N__24283\,
            lcout => scaler_2_data_13,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_9\,
            clk => \N__29338\,
            ce => \N__26377\,
            sr => \N__28726\
        );

    \scaler_2.source_data_1_esr_14_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24280\,
            lcout => scaler_2_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29338\,
            ce => \N__26377\,
            sr => \N__28726\
        );

    \scaler_2.source_data_1_esr_5_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25242\,
            in1 => \N__25276\,
            in2 => \_gnd_net_\,
            in3 => \N__25210\,
            lcout => scaler_2_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29330\,
            ce => \N__26380\,
            sr => \N__28731\
        );

    \scaler_3.source_data_1_esr_5_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27517\,
            in1 => \N__29734\,
            in2 => \_gnd_net_\,
            in3 => \N__27490\,
            lcout => scaler_3_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29330\,
            ce => \N__26380\,
            sr => \N__28731\
        );

    \scaler_4.source_data_1_esr_5_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25818\,
            in1 => \N__25852\,
            in2 => \_gnd_net_\,
            in3 => \N__26812\,
            lcout => scaler_4_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29330\,
            ce => \N__26380\,
            sr => \N__28731\
        );

    \uart_drone.data_Aux_RNO_0_0_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__26264\,
            in1 => \N__26335\,
            in2 => \_gnd_net_\,
            in3 => \N__26094\,
            lcout => \uart_drone.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27374\,
            lcout => \Commands_frame_decoder.preinitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29321\,
            ce => 'H',
            sr => \N__28736\
        );

    \scaler_2.source_data_1_4_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__27347\,
            in1 => \N__25243\,
            in2 => \N__24198\,
            in3 => \N__25209\,
            lcout => scaler_2_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29321\,
            ce => 'H',
            sr => \N__28736\
        );

    \scaler_3.source_data_1_4_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__27349\,
            in1 => \N__29730\,
            in2 => \N__24498\,
            in3 => \N__27489\,
            lcout => scaler_3_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29321\,
            ce => 'H',
            sr => \N__28736\
        );

    \scaler_4.source_data_1_4_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__27348\,
            in1 => \N__25860\,
            in2 => \N__24468\,
            in3 => \N__26811\,
            lcout => scaler_4_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29321\,
            ce => 'H',
            sr => \N__28736\
        );

    \Commands_frame_decoder.state_1_RNI2D06_1_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26183\,
            in2 => \_gnd_net_\,
            in3 => \N__24343\,
            lcout => \Commands_frame_decoder.N_282_0\,
            ltout => \Commands_frame_decoder.N_282_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_2_0_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28309\,
            in1 => \N__27852\,
            in2 => \N__24451\,
            in3 => \N__24447\,
            lcout => \Commands_frame_decoder.N_318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_3_0_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29847\,
            in1 => \N__28311\,
            in2 => \N__24353\,
            in3 => \N__24433\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNO_0_0_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010101"
        )
    port map (
            in0 => \N__26163\,
            in1 => \N__24381\,
            in2 => \N__24418\,
            in3 => \N__24415\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_1_ns_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_0_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__24409\,
            in1 => \N__24403\,
            in2 => \N__24397\,
            in3 => \N__29461\,
            lcout => \Commands_frame_decoder.state_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29310\,
            ce => 'H',
            sr => \N__28741\
        );

    \Commands_frame_decoder.state_1_10_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__29462\,
            in1 => \N__29698\,
            in2 => \N__26167\,
            in3 => \N__26184\,
            lcout => \Commands_frame_decoder.state_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29310\,
            ce => 'H',
            sr => \N__28741\
        );

    \Commands_frame_decoder.state_1_1_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24382\,
            in1 => \N__24367\,
            in2 => \N__24354\,
            in3 => \N__29460\,
            lcout => \Commands_frame_decoder.state_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29310\,
            ce => 'H',
            sr => \N__28741\
        );

    \uart_drone.bit_Count_2_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__25489\,
            in1 => \N__26737\,
            in2 => \N__26336\,
            in3 => \N__26253\,
            lcout => \uart_drone.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29302\,
            ce => 'H',
            sr => \N__28747\
        );

    \uart_drone.bit_Count_1_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__26252\,
            in1 => \N__25488\,
            in2 => \N__26149\,
            in3 => \N__26090\,
            lcout => \uart_drone.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29302\,
            ce => 'H',
            sr => \N__28747\
        );

    \ppm_encoder_1.un1_elevator_cry_6_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25986\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25959\,
            in2 => \_gnd_net_\,
            in3 => \N__24571\,
            lcout => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_6\,
            carryout => \ppm_encoder_1.un1_elevator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25935\,
            in2 => \_gnd_net_\,
            in3 => \N__24556\,
            lcout => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_7\,
            carryout => \ppm_encoder_1.un1_elevator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25911\,
            in2 => \_gnd_net_\,
            in3 => \N__24538\,
            lcout => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_8\,
            carryout => \ppm_encoder_1.un1_elevator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25887\,
            in2 => \_gnd_net_\,
            in3 => \N__24526\,
            lcout => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_9\,
            carryout => \ppm_encoder_1.un1_elevator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26478\,
            in2 => \_gnd_net_\,
            in3 => \N__24523\,
            lcout => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_10\,
            carryout => \ppm_encoder_1.un1_elevator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26451\,
            in2 => \_gnd_net_\,
            in3 => \N__24511\,
            lcout => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_11\,
            carryout => \ppm_encoder_1.un1_elevator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26421\,
            in2 => \N__27297\,
            in3 => \N__25105\,
            lcout => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_12\,
            carryout => \ppm_encoder_1.un1_elevator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_esr_14_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26392\,
            in2 => \_gnd_net_\,
            in3 => \N__25102\,
            lcout => \ppm_encoder_1.elevatorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29286\,
            ce => \N__25077\,
            sr => \N__28761\
        );

    \ppm_encoder_1.elevator_13_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__26425\,
            in1 => \N__25015\,
            in2 => \N__25001\,
            in3 => \N__24913\,
            lcout => \ppm_encoder_1.elevatorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29274\,
            ce => 'H',
            sr => \N__28773\
        );

    \ppm_encoder_1.elevator_11_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__26479\,
            in1 => \N__24976\,
            in2 => \N__24961\,
            in3 => \N__24674\,
            lcout => \ppm_encoder_1.elevatorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29266\,
            ce => 'H',
            sr => \N__28779\
        );

    \Commands_frame_decoder.state_1_RNITK1O_4_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24651\,
            in2 => \_gnd_net_\,
            in3 => \N__28934\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH4data_ess_7_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27648\,
            lcout => \frame_decoder_CH4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29339\,
            ce => \N__26773\,
            sr => \N__28719\
        );

    \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25155\,
            in2 => \_gnd_net_\,
            in3 => \N__24633\,
            lcout => \scaler_4.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.N_545_i_l_ofx_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25156\,
            in2 => \_gnd_net_\,
            in3 => \N__24634\,
            lcout => \scaler_4.N_545_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNI0O1O_7_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29505\,
            in2 => \_gnd_net_\,
            in3 => \N__28927\,
            lcout => \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__25275\,
            in1 => \N__25234\,
            in2 => \_gnd_net_\,
            in3 => \N__25208\,
            lcout => \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset4data_esr_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28356\,
            lcout => \frame_decoder_OFF4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29323\,
            ce => \N__29683\,
            sr => \N__28727\
        );

    \Commands_frame_decoder.source_offset4data_esr_4_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28001\,
            lcout => \frame_decoder_OFF4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29323\,
            ce => \N__29683\,
            sr => \N__28727\
        );

    \Commands_frame_decoder.source_offset4data_esr_0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29856\,
            lcout => \frame_decoder_OFF4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29323\,
            ce => \N__29683\,
            sr => \N__28727\
        );

    \Commands_frame_decoder.source_offset4data_esr_5_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27870\,
            lcout => \frame_decoder_OFF4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29323\,
            ce => \N__29683\,
            sr => \N__28727\
        );

    \Commands_frame_decoder.source_offset4data_esr_1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27768\,
            lcout => \frame_decoder_OFF4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29323\,
            ce => \N__29683\,
            sr => \N__28727\
        );

    \Commands_frame_decoder.source_offset4data_ess_7_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27639\,
            lcout => \frame_decoder_OFF4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29323\,
            ce => \N__29683\,
            sr => \N__28727\
        );

    \scaler_4.un2_source_data_0_cry_1_c_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25802\,
            in2 => \N__25147\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_6_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25767\,
            in2 => \N__25811\,
            in3 => \N__25108\,
            lcout => scaler_4_data_6,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_1\,
            carryout => \scaler_4.un2_source_data_0_cry_2\,
            clk => \N__29312\,
            ce => \N__26375\,
            sr => \N__28732\
        );

    \scaler_4.source_data_1_esr_7_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25746\,
            in2 => \N__25771\,
            in3 => \N__25444\,
            lcout => scaler_4_data_7,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_2\,
            carryout => \scaler_4.un2_source_data_0_cry_3\,
            clk => \N__29312\,
            ce => \N__26375\,
            sr => \N__28732\
        );

    \scaler_4.source_data_1_esr_8_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25713\,
            in2 => \N__25750\,
            in3 => \N__25420\,
            lcout => scaler_4_data_8,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_3\,
            carryout => \scaler_4.un2_source_data_0_cry_4\,
            clk => \N__29312\,
            ce => \N__26375\,
            sr => \N__28732\
        );

    \scaler_4.source_data_1_esr_9_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25683\,
            in2 => \N__25717\,
            in3 => \N__25396\,
            lcout => scaler_4_data_9,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_4\,
            carryout => \scaler_4.un2_source_data_0_cry_5\,
            clk => \N__29312\,
            ce => \N__26375\,
            sr => \N__28732\
        );

    \scaler_4.source_data_1_esr_10_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25659\,
            in2 => \N__25687\,
            in3 => \N__25372\,
            lcout => scaler_4_data_10,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_5\,
            carryout => \scaler_4.un2_source_data_0_cry_6\,
            clk => \N__29312\,
            ce => \N__26375\,
            sr => \N__28732\
        );

    \scaler_4.source_data_1_esr_11_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25638\,
            in2 => \N__25663\,
            in3 => \N__25348\,
            lcout => scaler_4_data_11,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_6\,
            carryout => \scaler_4.un2_source_data_0_cry_7\,
            clk => \N__29312\,
            ce => \N__26375\,
            sr => \N__28732\
        );

    \scaler_4.source_data_1_esr_12_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26022\,
            in2 => \N__25642\,
            in3 => \N__25324\,
            lcout => scaler_4_data_12,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_7\,
            carryout => \scaler_4.un2_source_data_0_cry_8\,
            clk => \N__29312\,
            ce => \N__26375\,
            sr => \N__28732\
        );

    \scaler_4.source_data_1_esr_13_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26023\,
            in2 => \N__26005\,
            in3 => \N__25297\,
            lcout => scaler_4_data_13,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_9\,
            clk => \N__29304\,
            ce => \N__26378\,
            sr => \N__28737\
        );

    \scaler_4.source_data_1_esr_14_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25294\,
            lcout => scaler_4_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29304\,
            ce => \N__26378\,
            sr => \N__28737\
        );

    \uart_drone.bit_Count_0_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001100100"
        )
    port map (
            in0 => \N__26148\,
            in1 => \N__26108\,
            in2 => \N__25588\,
            in3 => \N__25524\,
            lcout => \uart_drone.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29293\,
            ce => 'H',
            sr => \N__28742\
        );

    \Commands_frame_decoder.state_1_7_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__25480\,
            in1 => \N__29649\,
            in2 => \N__25627\,
            in3 => \N__29463\,
            lcout => \Commands_frame_decoder.state_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29293\,
            ce => 'H',
            sr => \N__28742\
        );

    \uart_drone.state_RNI63LK2_3_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__25587\,
            in1 => \N__26137\,
            in2 => \_gnd_net_\,
            in3 => \N__25523\,
            lcout => \uart_drone.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNI3BRE_7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25479\,
            in2 => \_gnd_net_\,
            in3 => \N__29648\,
            lcout => \Commands_frame_decoder.source_offset2data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH3data_esr_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29849\,
            lcout => \frame_decoder_CH3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29331\,
            ce => \N__27404\,
            sr => \N__28724\
        );

    \Commands_frame_decoder.source_CH4data_esr_2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28353\,
            lcout => \frame_decoder_CH4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29324\,
            ce => \N__26774\,
            sr => \N__28728\
        );

    \Commands_frame_decoder.source_CH4data_esr_3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28115\,
            lcout => \frame_decoder_CH4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29324\,
            ce => \N__26774\,
            sr => \N__28728\
        );

    \Commands_frame_decoder.source_CH4data_esr_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28000\,
            lcout => \frame_decoder_CH4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29324\,
            ce => \N__26774\,
            sr => \N__28728\
        );

    \Commands_frame_decoder.source_CH4data_esr_5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27890\,
            lcout => \frame_decoder_CH4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29324\,
            ce => \N__26774\,
            sr => \N__28728\
        );

    \Commands_frame_decoder.source_CH4data_esr_6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28231\,
            lcout => \frame_decoder_CH4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29324\,
            ce => \N__26774\,
            sr => \N__28728\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26793\,
            in2 => \N__25856\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25825\,
            in2 => \N__26824\,
            in3 => \N__25789\,
            lcout => \scaler_4.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_0\,
            carryout => \scaler_4.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25786\,
            in2 => \N__25780\,
            in3 => \N__25759\,
            lcout => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_1\,
            carryout => \scaler_4.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25756\,
            in2 => \N__28387\,
            in3 => \N__25738\,
            lcout => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_2\,
            carryout => \scaler_4.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25735\,
            in2 => \N__25729\,
            in3 => \N__25705\,
            lcout => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_3\,
            carryout => \scaler_4.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25702\,
            in2 => \N__25696\,
            in3 => \N__25675\,
            lcout => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_4\,
            carryout => \scaler_4.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25672\,
            in2 => \N__28375\,
            in3 => \N__25651\,
            lcout => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_5\,
            carryout => \scaler_4.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25648\,
            in2 => \_gnd_net_\,
            in3 => \N__25630\,
            lcout => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_6\,
            carryout => \scaler_4.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26032\,
            in2 => \N__27307\,
            in3 => \N__26011\,
            lcout => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26008\,
            lcout => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27508\,
            in2 => \N__27454\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.source_data_1_esr_6_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26973\,
            in2 => \N__27516\,
            in3 => \N__25969\,
            lcout => scaler_3_data_6,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_1\,
            carryout => \scaler_3.un2_source_data_0_cry_2\,
            clk => \N__29294\,
            ce => \N__26376\,
            sr => \N__28743\
        );

    \scaler_3.source_data_1_esr_7_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26952\,
            in2 => \N__26977\,
            in3 => \N__25942\,
            lcout => scaler_3_data_7,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_2\,
            carryout => \scaler_3.un2_source_data_0_cry_3\,
            clk => \N__29294\,
            ce => \N__26376\,
            sr => \N__28743\
        );

    \scaler_3.source_data_1_esr_8_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26931\,
            in2 => \N__26956\,
            in3 => \N__25918\,
            lcout => scaler_3_data_8,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_3\,
            carryout => \scaler_3.un2_source_data_0_cry_4\,
            clk => \N__29294\,
            ce => \N__26376\,
            sr => \N__28743\
        );

    \scaler_3.source_data_1_esr_9_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26907\,
            in2 => \N__26935\,
            in3 => \N__25891\,
            lcout => scaler_3_data_9,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_4\,
            carryout => \scaler_3.un2_source_data_0_cry_5\,
            clk => \N__29294\,
            ce => \N__26376\,
            sr => \N__28743\
        );

    \scaler_3.source_data_1_esr_10_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26886\,
            in2 => \N__26911\,
            in3 => \N__25864\,
            lcout => scaler_3_data_10,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_5\,
            carryout => \scaler_3.un2_source_data_0_cry_6\,
            clk => \N__29294\,
            ce => \N__26376\,
            sr => \N__28743\
        );

    \scaler_3.source_data_1_esr_11_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26871\,
            in2 => \N__26890\,
            in3 => \N__26455\,
            lcout => scaler_3_data_11,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_6\,
            carryout => \scaler_3.un2_source_data_0_cry_7\,
            clk => \N__29294\,
            ce => \N__26376\,
            sr => \N__28743\
        );

    \scaler_3.source_data_1_esr_12_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26859\,
            in2 => \N__26875\,
            in3 => \N__26428\,
            lcout => scaler_3_data_12,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_7\,
            carryout => \scaler_3.un2_source_data_0_cry_8\,
            clk => \N__29294\,
            ce => \N__26376\,
            sr => \N__28743\
        );

    \scaler_3.source_data_1_esr_13_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26860\,
            in2 => \N__26842\,
            in3 => \N__26398\,
            lcout => scaler_3_data_13,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_9\,
            clk => \N__29287\,
            ce => \N__26379\,
            sr => \N__28748\
        );

    \scaler_3.source_data_1_esr_14_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26395\,
            lcout => scaler_3_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29287\,
            ce => \N__26379\,
            sr => \N__28748\
        );

    \uart_drone.data_Aux_RNO_0_1_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__26073\,
            in1 => \N__26334\,
            in2 => \_gnd_net_\,
            in3 => \N__26263\,
            lcout => \uart_drone.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_data_valid_RNO_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__26194\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26713\,
            lcout => \Commands_frame_decoder.count_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNIDIPF_10_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29647\,
            in2 => \_gnd_net_\,
            in3 => \N__26193\,
            lcout => \Commands_frame_decoder.state_1_ns_i_a4_2_0_0\,
            ltout => \Commands_frame_decoder.state_1_ns_i_a4_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNI0PVH1_2_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__26521\,
            in1 => \N__26497\,
            in2 => \N__26170\,
            in3 => \N__27003\,
            lcout => \Commands_frame_decoder.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNO_0_2_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26147\,
            in2 => \_gnd_net_\,
            in3 => \N__26072\,
            lcout => \uart_drone.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count8_cry_0_c_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27042\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \Commands_frame_decoder.count8_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count8_cry_1_c_inv_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26728\,
            in2 => \_gnd_net_\,
            in3 => \N__26494\,
            lcout => \Commands_frame_decoder.count8_axb_1\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.count8_cry_0\,
            carryout => \Commands_frame_decoder.count8_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count8_cry_2_c_inv_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26722\,
            in2 => \N__27299\,
            in3 => \N__26519\,
            lcout => \Commands_frame_decoder.count_i_2\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.count8_cry_1\,
            carryout => \Commands_frame_decoder.count8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count8_THRU_LUT4_0_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26716\,
            lcout => \Commands_frame_decoder.count8_THRU_CO\,
            ltout => \Commands_frame_decoder.count8_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count8_cry_2_c_RNIARGV_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__26657\,
            in1 => \_gnd_net_\,
            in2 => \N__26527\,
            in3 => \N__27018\,
            lcout => \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0\,
            ltout => \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_2_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010100000"
        )
    port map (
            in0 => \N__26520\,
            in1 => \N__26506\,
            in2 => \N__26524\,
            in3 => \N__26496\,
            lcout => \Commands_frame_decoder.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNIT86R_0_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27017\,
            in2 => \_gnd_net_\,
            in3 => \N__27004\,
            lcout => \Commands_frame_decoder.CO0\,
            ltout => \Commands_frame_decoder.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_1_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27030\,
            in2 => \N__26500\,
            in3 => \N__26495\,
            lcout => \Commands_frame_decoder.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_ctle_14_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27346\,
            in2 => \_gnd_net_\,
            in3 => \N__28924\,
            lcout => pc_frame_decoder_dv_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH4data_esr_1_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27775\,
            lcout => \frame_decoder_CH4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29322\,
            ce => \N__26782\,
            sr => \N__28729\
        );

    \Commands_frame_decoder.source_CH4data_esr_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29848\,
            lcout => \frame_decoder_CH4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29311\,
            ce => \N__26781\,
            sr => \N__28733\
        );

    \Commands_frame_decoder.source_CH3data_esr_4_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28002\,
            lcout => \frame_decoder_CH3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29303\,
            ce => \N__27417\,
            sr => \N__28738\
        );

    \Commands_frame_decoder.source_CH3data_esr_2_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28360\,
            lcout => \frame_decoder_CH3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29303\,
            ce => \N__27417\,
            sr => \N__28738\
        );

    \Commands_frame_decoder.source_CH3data_esr_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28106\,
            lcout => \frame_decoder_CH3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29303\,
            ce => \N__27417\,
            sr => \N__28738\
        );

    \Commands_frame_decoder.source_CH3data_esr_5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27891\,
            lcout => \frame_decoder_CH3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29303\,
            ce => \N__27417\,
            sr => \N__28738\
        );

    \Commands_frame_decoder.source_CH3data_esr_6_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28228\,
            lcout => \frame_decoder_CH3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29303\,
            ce => \N__27417\,
            sr => \N__28738\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27487\,
            in2 => \N__29729\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27439\,
            in2 => \N__27658\,
            in3 => \N__26740\,
            lcout => \scaler_3.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_0\,
            carryout => \scaler_3.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26983\,
            in2 => \N__28240\,
            in3 => \N__26965\,
            lcout => \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_1\,
            carryout => \scaler_3.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26962\,
            in2 => \N__28012\,
            in3 => \N__26944\,
            lcout => \scaler_3.un3_source_data_0_cry_2_c_RNI780L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_2\,
            carryout => \scaler_3.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26941\,
            in2 => \N__27901\,
            in3 => \N__26923\,
            lcout => \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_3\,
            carryout => \scaler_3.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27781\,
            in2 => \N__26920\,
            in3 => \N__26899\,
            lcout => \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_4\,
            carryout => \scaler_3.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26896\,
            in2 => \N__28126\,
            in3 => \N__26878\,
            lcout => \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_5\,
            carryout => \scaler_3.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27445\,
            in2 => \_gnd_net_\,
            in3 => \N__26863\,
            lcout => \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_6\,
            carryout => \scaler_3.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27523\,
            in2 => \N__27306\,
            in3 => \N__26848\,
            lcout => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26845\,
            lcout => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.N_533_i_l_ofx_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__27430\,
            in1 => \_gnd_net_\,
            in2 => \N__27535\,
            in3 => \_gnd_net_\,
            lcout => \scaler_3.N_533_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__27515\,
            in1 => \N__29722\,
            in2 => \_gnd_net_\,
            in3 => \N__27488\,
            lcout => \scaler_3.un2_source_data_0_cry_1_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27531\,
            in2 => \_gnd_net_\,
            in3 => \N__27429\,
            lcout => \scaler_3.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH3data_esr_1_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27763\,
            lcout => \frame_decoder_CH3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29282\,
            ce => \N__27421\,
            sr => \N__28754\
        );

    \Commands_frame_decoder.source_CH3data_ess_7_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27605\,
            lcout => \frame_decoder_CH3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29282\,
            ce => \N__27421\,
            sr => \N__28754\
        );

    \Commands_frame_decoder.source_data_valid_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__27387\,
            in1 => \N__29658\,
            in2 => \N__27337\,
            in3 => \N__27355\,
            lcout => pc_frame_decoder_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29275\,
            ce => 'H',
            sr => \N__28762\
        );

    \Commands_frame_decoder.count8_cry_0_c_inv_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__27043\,
            in1 => \N__27298\,
            in2 => \_gnd_net_\,
            in3 => \N__27001\,
            lcout => \Commands_frame_decoder.count8_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_0_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27031\,
            in1 => \N__27019\,
            in2 => \_gnd_net_\,
            in3 => \N__27002\,
            lcout => \Commands_frame_decoder.count8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset4data_esr_3_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28117\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29313\,
            ce => \N__29682\,
            sr => \N__28744\
        );

    \Commands_frame_decoder.source_offset4data_esr_6_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28229\,
            lcout => \frame_decoder_OFF4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29313\,
            ce => \N__29682\,
            sr => \N__28744\
        );

    \Commands_frame_decoder.source_offset3data_esr_2_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28363\,
            lcout => \frame_decoder_OFF3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29305\,
            ce => \N__29527\,
            sr => \N__28749\
        );

    \Commands_frame_decoder.source_offset3data_esr_6_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28194\,
            lcout => \frame_decoder_OFF3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29305\,
            ce => \N__29527\,
            sr => \N__28749\
        );

    \Commands_frame_decoder.source_offset3data_esr_3_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28116\,
            lcout => \frame_decoder_OFF3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29305\,
            ce => \N__29527\,
            sr => \N__28749\
        );

    \Commands_frame_decoder.source_offset3data_esr_4_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28003\,
            lcout => \frame_decoder_OFF3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29305\,
            ce => \N__29527\,
            sr => \N__28749\
        );

    \Commands_frame_decoder.source_offset3data_esr_5_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27892\,
            lcout => \frame_decoder_OFF3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29305\,
            ce => \N__29527\,
            sr => \N__28749\
        );

    \Commands_frame_decoder.source_offset3data_esr_1_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27770\,
            lcout => \frame_decoder_OFF3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29305\,
            ce => \N__29527\,
            sr => \N__28749\
        );

    \Commands_frame_decoder.source_offset3data_ess_7_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27646\,
            lcout => \frame_decoder_OFF3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29295\,
            ce => \N__29523\,
            sr => \N__28755\
        );

    \Commands_frame_decoder.source_offset3data_esr_0_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29839\,
            lcout => \frame_decoder_OFF3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29295\,
            ce => \N__29523\,
            sr => \N__28755\
        );

    \Commands_frame_decoder.state_1_RNI5DRE_9_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29656\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNI2Q1O_9_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29686\,
            in3 => \N__28937\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNI4CRE_8_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29481\,
            in2 => \_gnd_net_\,
            in3 => \N__29659\,
            lcout => \Commands_frame_decoder.source_offset3data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_offset3data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_RNI1P1O_8_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29530\,
            in3 => \N__28939\,
            lcout => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_8_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__29482\,
            in1 => \N__29506\,
            in2 => \_gnd_net_\,
            in3 => \N__29469\,
            lcout => \Commands_frame_decoder.state_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29296\,
            ce => 'H',
            sr => \N__28768\
        );

    \Commands_frame_decoder.state_1_9_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__29470\,
            in1 => \N__29410\,
            in2 => \_gnd_net_\,
            in3 => \N__29404\,
            lcout => \Commands_frame_decoder.state_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29296\,
            ce => 'H',
            sr => \N__28768\
        );
end \INTERFACE\;
